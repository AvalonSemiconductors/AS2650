magic
tech gf180mcuD
magscale 1 10
timestamp 1700712075
<< metal1 >>
rect 77298 57038 77310 57090
rect 77362 57087 77374 57090
rect 78082 57087 78094 57090
rect 77362 57041 78094 57087
rect 77362 57038 77374 57041
rect 78082 57038 78094 57041
rect 78146 57038 78158 57090
rect 157378 57038 157390 57090
rect 157442 57087 157454 57090
rect 157938 57087 157950 57090
rect 157442 57041 157950 57087
rect 157442 57038 157454 57041
rect 157938 57038 157950 57041
rect 158002 57087 158014 57090
rect 158498 57087 158510 57090
rect 158002 57041 158510 57087
rect 158002 57038 158014 57041
rect 158498 57038 158510 57041
rect 158562 57038 158574 57090
rect 270834 57038 270846 57090
rect 270898 57087 270910 57090
rect 271506 57087 271518 57090
rect 270898 57041 271518 57087
rect 270898 57038 270910 57041
rect 271506 57038 271518 57041
rect 271570 57038 271582 57090
rect 11890 56590 11902 56642
rect 11954 56639 11966 56642
rect 13122 56639 13134 56642
rect 11954 56593 13134 56639
rect 11954 56590 11966 56593
rect 13122 56590 13134 56593
rect 13186 56590 13198 56642
rect 23538 56590 23550 56642
rect 23602 56639 23614 56642
rect 24098 56639 24110 56642
rect 23602 56593 24110 56639
rect 23602 56590 23614 56593
rect 24098 56590 24110 56593
rect 24162 56639 24174 56642
rect 24546 56639 24558 56642
rect 24162 56593 24558 56639
rect 24162 56590 24174 56593
rect 24546 56590 24558 56593
rect 24610 56590 24622 56642
rect 114930 56590 114942 56642
rect 114994 56639 115006 56642
rect 115490 56639 115502 56642
rect 114994 56593 115502 56639
rect 114994 56590 115006 56593
rect 115490 56590 115502 56593
rect 115554 56639 115566 56642
rect 115938 56639 115950 56642
rect 115554 56593 115950 56639
rect 115554 56590 115566 56593
rect 115938 56590 115950 56593
rect 116002 56590 116014 56642
rect 168690 56590 168702 56642
rect 168754 56639 168766 56642
rect 169586 56639 169598 56642
rect 168754 56593 169598 56639
rect 168754 56590 168766 56593
rect 169586 56590 169598 56593
rect 169650 56590 169662 56642
rect 190194 56590 190206 56642
rect 190258 56639 190270 56642
rect 191426 56639 191438 56642
rect 190258 56593 191438 56639
rect 190258 56590 190270 56593
rect 191426 56590 191438 56593
rect 191490 56639 191502 56642
rect 192210 56639 192222 56642
rect 191490 56593 192222 56639
rect 191490 56590 191502 56593
rect 192210 56590 192222 56593
rect 192274 56590 192286 56642
rect 222114 56590 222126 56642
rect 222178 56639 222190 56642
rect 223010 56639 223022 56642
rect 222178 56593 223022 56639
rect 222178 56590 222190 56593
rect 223010 56590 223022 56593
rect 223074 56590 223086 56642
rect 1344 56474 298592 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 81278 56474
rect 81330 56422 81382 56474
rect 81434 56422 81486 56474
rect 81538 56422 111998 56474
rect 112050 56422 112102 56474
rect 112154 56422 112206 56474
rect 112258 56422 142718 56474
rect 142770 56422 142822 56474
rect 142874 56422 142926 56474
rect 142978 56422 173438 56474
rect 173490 56422 173542 56474
rect 173594 56422 173646 56474
rect 173698 56422 204158 56474
rect 204210 56422 204262 56474
rect 204314 56422 204366 56474
rect 204418 56422 234878 56474
rect 234930 56422 234982 56474
rect 235034 56422 235086 56474
rect 235138 56422 265598 56474
rect 265650 56422 265702 56474
rect 265754 56422 265806 56474
rect 265858 56422 296318 56474
rect 296370 56422 296422 56474
rect 296474 56422 296526 56474
rect 296578 56422 298592 56474
rect 1344 56388 298592 56422
rect 12686 56306 12738 56318
rect 12686 56242 12738 56254
rect 18174 56306 18226 56318
rect 18174 56242 18226 56254
rect 18398 56306 18450 56318
rect 18398 56242 18450 56254
rect 19182 56306 19234 56318
rect 19182 56242 19234 56254
rect 24110 56306 24162 56318
rect 24110 56242 24162 56254
rect 24558 56306 24610 56318
rect 24558 56242 24610 56254
rect 28926 56306 28978 56318
rect 28926 56242 28978 56254
rect 29150 56306 29202 56318
rect 29150 56242 29202 56254
rect 34302 56306 34354 56318
rect 34302 56242 34354 56254
rect 34526 56306 34578 56318
rect 34526 56242 34578 56254
rect 39342 56306 39394 56318
rect 39342 56242 39394 56254
rect 39902 56306 39954 56318
rect 39902 56242 39954 56254
rect 45054 56306 45106 56318
rect 45054 56242 45106 56254
rect 45278 56306 45330 56318
rect 45278 56242 45330 56254
rect 50766 56306 50818 56318
rect 50766 56242 50818 56254
rect 51214 56306 51266 56318
rect 51214 56242 51266 56254
rect 55806 56306 55858 56318
rect 55806 56242 55858 56254
rect 56030 56306 56082 56318
rect 56030 56242 56082 56254
rect 61182 56306 61234 56318
rect 61182 56242 61234 56254
rect 61406 56306 61458 56318
rect 61406 56242 61458 56254
rect 109566 56306 109618 56318
rect 109566 56242 109618 56254
rect 109790 56306 109842 56318
rect 109790 56242 109842 56254
rect 115502 56306 115554 56318
rect 115502 56242 115554 56254
rect 115950 56306 116002 56318
rect 115950 56242 116002 56254
rect 120318 56306 120370 56318
rect 120318 56242 120370 56254
rect 120542 56306 120594 56318
rect 120542 56242 120594 56254
rect 125694 56306 125746 56318
rect 125694 56242 125746 56254
rect 125918 56306 125970 56318
rect 125918 56242 125970 56254
rect 130734 56306 130786 56318
rect 130734 56242 130786 56254
rect 136446 56306 136498 56318
rect 136446 56242 136498 56254
rect 142158 56306 142210 56318
rect 142158 56242 142210 56254
rect 147198 56306 147250 56318
rect 147198 56242 147250 56254
rect 152574 56306 152626 56318
rect 152574 56242 152626 56254
rect 157390 56306 157442 56318
rect 157390 56242 157442 56254
rect 163326 56306 163378 56318
rect 163326 56242 163378 56254
rect 168814 56306 168866 56318
rect 168814 56242 168866 56254
rect 174078 56306 174130 56318
rect 174078 56242 174130 56254
rect 179454 56306 179506 56318
rect 179454 56242 179506 56254
rect 184830 56306 184882 56318
rect 184830 56242 184882 56254
rect 192222 56306 192274 56318
rect 192222 56242 192274 56254
rect 195470 56306 195522 56318
rect 195470 56242 195522 56254
rect 208350 56306 208402 56318
rect 208350 56242 208402 56254
rect 211710 56306 211762 56318
rect 211710 56242 211762 56254
rect 211934 56306 211986 56318
rect 211934 56242 211986 56254
rect 217086 56306 217138 56318
rect 217086 56242 217138 56254
rect 222126 56306 222178 56318
rect 222126 56242 222178 56254
rect 223022 56306 223074 56318
rect 223022 56242 223074 56254
rect 227838 56306 227890 56318
rect 227838 56242 227890 56254
rect 233550 56306 233602 56318
rect 233550 56242 233602 56254
rect 238590 56306 238642 56318
rect 238590 56242 238642 56254
rect 238814 56306 238866 56318
rect 238814 56242 238866 56254
rect 243966 56306 244018 56318
rect 243966 56242 244018 56254
rect 244190 56306 244242 56318
rect 244190 56242 244242 56254
rect 248782 56306 248834 56318
rect 248782 56242 248834 56254
rect 249566 56306 249618 56318
rect 249566 56242 249618 56254
rect 254718 56306 254770 56318
rect 254718 56242 254770 56254
rect 260094 56306 260146 56318
rect 260094 56242 260146 56254
rect 265470 56306 265522 56318
rect 265470 56242 265522 56254
rect 271518 56306 271570 56318
rect 271518 56242 271570 56254
rect 276222 56306 276274 56318
rect 276222 56242 276274 56254
rect 286862 56306 286914 56318
rect 286862 56242 286914 56254
rect 287310 56306 287362 56318
rect 287310 56242 287362 56254
rect 292350 56306 292402 56318
rect 292350 56242 292402 56254
rect 292574 56306 292626 56318
rect 292574 56242 292626 56254
rect 131294 56194 131346 56206
rect 13122 56142 13134 56194
rect 13186 56142 13198 56194
rect 126242 56142 126254 56194
rect 126306 56142 126318 56194
rect 131294 56130 131346 56142
rect 131630 56194 131682 56206
rect 131630 56130 131682 56142
rect 136670 56194 136722 56206
rect 136670 56130 136722 56142
rect 142606 56194 142658 56206
rect 142606 56130 142658 56142
rect 147422 56194 147474 56206
rect 147422 56130 147474 56142
rect 152798 56194 152850 56206
rect 152798 56130 152850 56142
rect 153134 56194 153186 56206
rect 153134 56130 153186 56142
rect 158174 56194 158226 56206
rect 158174 56130 158226 56142
rect 158510 56194 158562 56206
rect 158510 56130 158562 56142
rect 163550 56194 163602 56206
rect 163550 56130 163602 56142
rect 169262 56194 169314 56206
rect 169262 56130 169314 56142
rect 169598 56194 169650 56206
rect 169598 56130 169650 56142
rect 174302 56194 174354 56206
rect 174302 56130 174354 56142
rect 179678 56194 179730 56206
rect 179678 56130 179730 56142
rect 180014 56194 180066 56206
rect 180014 56130 180066 56142
rect 185054 56194 185106 56206
rect 185054 56130 185106 56142
rect 189870 56194 189922 56206
rect 189870 56130 189922 56142
rect 191214 56194 191266 56206
rect 191214 56130 191266 56142
rect 195918 56194 195970 56206
rect 212258 56142 212270 56194
rect 212322 56142 212334 56194
rect 217298 56142 217310 56194
rect 217362 56142 217374 56194
rect 222674 56142 222686 56194
rect 222738 56142 222750 56194
rect 228050 56142 228062 56194
rect 228114 56142 228126 56194
rect 233986 56142 233998 56194
rect 234050 56142 234062 56194
rect 195918 56130 195970 56142
rect 85710 56082 85762 56094
rect 92430 56082 92482 56094
rect 107662 56082 107714 56094
rect 206894 56082 206946 56094
rect 283614 56082 283666 56094
rect 13346 56030 13358 56082
rect 13410 56030 13422 56082
rect 69346 56030 69358 56082
rect 69410 56030 69422 56082
rect 80434 56030 80446 56082
rect 80498 56030 80510 56082
rect 84914 56030 84926 56082
rect 84978 56030 84990 56082
rect 91858 56030 91870 56082
rect 91922 56030 91934 56082
rect 96226 56030 96238 56082
rect 96290 56030 96302 56082
rect 107090 56030 107102 56082
rect 107154 56030 107166 56082
rect 136882 56030 136894 56082
rect 136946 56030 136958 56082
rect 142818 56030 142830 56082
rect 142882 56030 142894 56082
rect 147634 56030 147646 56082
rect 147698 56030 147710 56082
rect 163762 56030 163774 56082
rect 163826 56030 163838 56082
rect 174514 56030 174526 56082
rect 174578 56030 174590 56082
rect 185266 56030 185278 56082
rect 185330 56030 185342 56082
rect 190866 56030 190878 56082
rect 190930 56030 190942 56082
rect 191426 56030 191438 56082
rect 191490 56030 191502 56082
rect 196130 56030 196142 56082
rect 196194 56030 196206 56082
rect 202962 56030 202974 56082
rect 203026 56030 203038 56082
rect 207330 56030 207342 56082
rect 207394 56030 207406 56082
rect 217522 56030 217534 56082
rect 217586 56030 217598 56082
rect 228274 56030 228286 56082
rect 228338 56030 228350 56082
rect 234210 56030 234222 56082
rect 234274 56030 234286 56082
rect 254930 56030 254942 56082
rect 254994 56030 255006 56082
rect 260754 56030 260766 56082
rect 260818 56030 260830 56082
rect 265682 56030 265694 56082
rect 265746 56030 265758 56082
rect 272178 56030 272190 56082
rect 272242 56030 272254 56082
rect 276434 56030 276446 56082
rect 276498 56030 276510 56082
rect 282706 56030 282718 56082
rect 282770 56030 282782 56082
rect 85710 56018 85762 56030
rect 92430 56018 92482 56030
rect 107662 56018 107714 56030
rect 206894 56018 206946 56030
rect 283614 56018 283666 56030
rect 25118 55970 25170 55982
rect 25118 55906 25170 55918
rect 29710 55970 29762 55982
rect 29710 55906 29762 55918
rect 35086 55970 35138 55982
rect 35086 55906 35138 55918
rect 40462 55970 40514 55982
rect 40462 55906 40514 55918
rect 45838 55970 45890 55982
rect 45838 55906 45890 55918
rect 51774 55970 51826 55982
rect 51774 55906 51826 55918
rect 56590 55970 56642 55982
rect 56590 55906 56642 55918
rect 61966 55970 62018 55982
rect 61966 55906 62018 55918
rect 67006 55970 67058 55982
rect 67006 55906 67058 55918
rect 70478 55970 70530 55982
rect 70478 55906 70530 55918
rect 78094 55970 78146 55982
rect 78094 55906 78146 55918
rect 81006 55970 81058 55982
rect 89518 55970 89570 55982
rect 82674 55918 82686 55970
rect 82738 55918 82750 55970
rect 81006 55906 81058 55918
rect 89518 55906 89570 55918
rect 93886 55970 93938 55982
rect 93886 55906 93938 55918
rect 97134 55970 97186 55982
rect 97134 55906 97186 55918
rect 104750 55970 104802 55982
rect 104750 55906 104802 55918
rect 110350 55970 110402 55982
rect 110350 55906 110402 55918
rect 116510 55970 116562 55982
rect 116510 55906 116562 55918
rect 121102 55970 121154 55982
rect 121102 55906 121154 55918
rect 187854 55970 187906 55982
rect 187854 55906 187906 55918
rect 188526 55970 188578 55982
rect 188526 55906 188578 55918
rect 189086 55970 189138 55982
rect 203758 55970 203810 55982
rect 244750 55970 244802 55982
rect 200946 55918 200958 55970
rect 201010 55918 201022 55970
rect 239250 55918 239262 55970
rect 239314 55918 239326 55970
rect 189086 55906 189138 55918
rect 203758 55906 203810 55918
rect 244750 55906 244802 55918
rect 250126 55970 250178 55982
rect 256050 55918 256062 55970
rect 256114 55918 256126 55970
rect 261762 55918 261774 55970
rect 261826 55918 261838 55970
rect 266354 55918 266366 55970
rect 266418 55918 266430 55970
rect 273186 55918 273198 55970
rect 273250 55918 273262 55970
rect 277218 55918 277230 55970
rect 277282 55918 277294 55970
rect 281810 55918 281822 55970
rect 281874 55918 281886 55970
rect 250126 55906 250178 55918
rect 288094 55858 288146 55870
rect 288094 55794 288146 55806
rect 293358 55858 293410 55870
rect 293358 55794 293410 55806
rect 1344 55690 298592 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 96638 55690
rect 96690 55638 96742 55690
rect 96794 55638 96846 55690
rect 96898 55638 127358 55690
rect 127410 55638 127462 55690
rect 127514 55638 127566 55690
rect 127618 55638 158078 55690
rect 158130 55638 158182 55690
rect 158234 55638 158286 55690
rect 158338 55638 188798 55690
rect 188850 55638 188902 55690
rect 188954 55638 189006 55690
rect 189058 55638 219518 55690
rect 219570 55638 219622 55690
rect 219674 55638 219726 55690
rect 219778 55638 250238 55690
rect 250290 55638 250342 55690
rect 250394 55638 250446 55690
rect 250498 55638 280958 55690
rect 281010 55638 281062 55690
rect 281114 55638 281166 55690
rect 281218 55638 298592 55690
rect 1344 55604 298592 55638
rect 72382 55410 72434 55422
rect 156270 55410 156322 55422
rect 100034 55358 100046 55410
rect 100098 55358 100110 55410
rect 141250 55358 141262 55410
rect 141314 55358 141326 55410
rect 72382 55346 72434 55358
rect 156270 55346 156322 55358
rect 161870 55410 161922 55422
rect 186174 55410 186226 55422
rect 180226 55358 180238 55410
rect 180290 55358 180302 55410
rect 182354 55358 182366 55410
rect 182418 55358 182430 55410
rect 161870 55346 161922 55358
rect 186174 55346 186226 55358
rect 186398 55410 186450 55422
rect 188290 55358 188302 55410
rect 188354 55358 188366 55410
rect 190418 55358 190430 55410
rect 190482 55358 190494 55410
rect 186398 55346 186450 55358
rect 138350 55298 138402 55310
rect 143838 55298 143890 55310
rect 170382 55298 170434 55310
rect 175534 55298 175586 55310
rect 186062 55298 186114 55310
rect 74722 55246 74734 55298
rect 74786 55246 74798 55298
rect 102274 55246 102286 55298
rect 102338 55246 102350 55298
rect 135090 55246 135102 55298
rect 135154 55246 135166 55298
rect 140466 55246 140478 55298
rect 140530 55246 140542 55298
rect 152674 55246 152686 55298
rect 152738 55246 152750 55298
rect 156706 55246 156718 55298
rect 156770 55246 156782 55298
rect 162418 55246 162430 55298
rect 162482 55246 162494 55298
rect 169698 55246 169710 55298
rect 169762 55246 169774 55298
rect 174962 55246 174974 55298
rect 175026 55246 175038 55298
rect 179442 55246 179454 55298
rect 179506 55246 179518 55298
rect 138350 55234 138402 55246
rect 143838 55234 143890 55246
rect 170382 55234 170434 55246
rect 175534 55234 175586 55246
rect 186062 55234 186114 55246
rect 187182 55298 187234 55310
rect 191202 55246 191214 55298
rect 191266 55246 191278 55298
rect 187182 55234 187234 55246
rect 186510 55186 186562 55198
rect 135762 55134 135774 55186
rect 135826 55134 135838 55186
rect 147858 55134 147870 55186
rect 147922 55134 147934 55186
rect 157378 55134 157390 55186
rect 157442 55134 157454 55186
rect 163202 55134 163214 55186
rect 163266 55134 163278 55186
rect 168914 55134 168926 55186
rect 168978 55134 168990 55186
rect 174290 55134 174302 55186
rect 174354 55134 174366 55186
rect 186510 55122 186562 55134
rect 186846 55186 186898 55198
rect 186846 55122 186898 55134
rect 186958 55186 187010 55198
rect 186958 55122 187010 55134
rect 187518 55186 187570 55198
rect 187518 55122 187570 55134
rect 75182 55074 75234 55086
rect 75182 55010 75234 55022
rect 102734 55074 102786 55086
rect 102734 55010 102786 55022
rect 153246 55074 153298 55086
rect 153246 55010 153298 55022
rect 182814 55074 182866 55086
rect 182814 55010 182866 55022
rect 187966 55074 188018 55086
rect 187966 55010 188018 55022
rect 1344 54906 298592 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 81278 54906
rect 81330 54854 81382 54906
rect 81434 54854 81486 54906
rect 81538 54854 111998 54906
rect 112050 54854 112102 54906
rect 112154 54854 112206 54906
rect 112258 54854 142718 54906
rect 142770 54854 142822 54906
rect 142874 54854 142926 54906
rect 142978 54854 173438 54906
rect 173490 54854 173542 54906
rect 173594 54854 173646 54906
rect 173698 54854 204158 54906
rect 204210 54854 204262 54906
rect 204314 54854 204366 54906
rect 204418 54854 234878 54906
rect 234930 54854 234982 54906
rect 235034 54854 235086 54906
rect 235138 54854 265598 54906
rect 265650 54854 265702 54906
rect 265754 54854 265806 54906
rect 265858 54854 296318 54906
rect 296370 54854 296422 54906
rect 296474 54854 296526 54906
rect 296578 54854 298592 54906
rect 1344 54820 298592 54854
rect 132974 54738 133026 54750
rect 132974 54674 133026 54686
rect 135774 54738 135826 54750
rect 135774 54674 135826 54686
rect 141038 54738 141090 54750
rect 141038 54674 141090 54686
rect 148654 54738 148706 54750
rect 148654 54674 148706 54686
rect 150110 54738 150162 54750
rect 150110 54674 150162 54686
rect 157166 54738 157218 54750
rect 157166 54674 157218 54686
rect 162318 54738 162370 54750
rect 162318 54674 162370 54686
rect 167918 54738 167970 54750
rect 167918 54674 167970 54686
rect 172734 54738 172786 54750
rect 172734 54674 172786 54686
rect 184034 54574 184046 54626
rect 184098 54574 184110 54626
rect 193890 54574 193902 54626
rect 193954 54574 193966 54626
rect 191438 54514 191490 54526
rect 132514 54462 132526 54514
rect 132578 54462 132590 54514
rect 148082 54462 148094 54514
rect 148146 54462 148158 54514
rect 153906 54462 153918 54514
rect 153970 54462 153982 54514
rect 183250 54462 183262 54514
rect 183314 54462 183326 54514
rect 194562 54462 194574 54514
rect 194626 54462 194638 54514
rect 191438 54450 191490 54462
rect 182926 54402 182978 54414
rect 131730 54350 131742 54402
rect 131794 54350 131806 54402
rect 147410 54350 147422 54402
rect 147474 54350 147486 54402
rect 153122 54350 153134 54402
rect 153186 54350 153198 54402
rect 186162 54350 186174 54402
rect 186226 54350 186238 54402
rect 191762 54350 191774 54402
rect 191826 54350 191838 54402
rect 182926 54338 182978 54350
rect 134990 54290 135042 54302
rect 134990 54226 135042 54238
rect 140254 54290 140306 54302
rect 140254 54226 140306 54238
rect 156382 54290 156434 54302
rect 156382 54226 156434 54238
rect 161534 54290 161586 54302
rect 161534 54226 161586 54238
rect 167134 54290 167186 54302
rect 167134 54226 167186 54238
rect 171950 54290 172002 54302
rect 171950 54226 172002 54238
rect 1344 54122 298592 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 96638 54122
rect 96690 54070 96742 54122
rect 96794 54070 96846 54122
rect 96898 54070 127358 54122
rect 127410 54070 127462 54122
rect 127514 54070 127566 54122
rect 127618 54070 158078 54122
rect 158130 54070 158182 54122
rect 158234 54070 158286 54122
rect 158338 54070 188798 54122
rect 188850 54070 188902 54122
rect 188954 54070 189006 54122
rect 189058 54070 219518 54122
rect 219570 54070 219622 54122
rect 219674 54070 219726 54122
rect 219778 54070 250238 54122
rect 250290 54070 250342 54122
rect 250394 54070 250446 54122
rect 250498 54070 280958 54122
rect 281010 54070 281062 54122
rect 281114 54070 281166 54122
rect 281218 54070 298592 54122
rect 1344 54036 298592 54070
rect 180114 53790 180126 53842
rect 180178 53790 180190 53842
rect 193218 53790 193230 53842
rect 193282 53790 193294 53842
rect 145966 53730 146018 53742
rect 130274 53678 130286 53730
rect 130338 53678 130350 53730
rect 145966 53666 146018 53678
rect 151566 53730 151618 53742
rect 151566 53666 151618 53678
rect 161982 53730 162034 53742
rect 189758 53730 189810 53742
rect 162418 53678 162430 53730
rect 162482 53678 162494 53730
rect 178098 53678 178110 53730
rect 178162 53678 178174 53730
rect 190418 53678 190430 53730
rect 190482 53678 190494 53730
rect 161982 53666 162034 53678
rect 189758 53666 189810 53678
rect 177662 53618 177714 53630
rect 129378 53566 129390 53618
rect 129442 53566 129454 53618
rect 167458 53566 167470 53618
rect 167522 53566 167534 53618
rect 191090 53566 191102 53618
rect 191154 53566 191166 53618
rect 177662 53554 177714 53566
rect 145182 53506 145234 53518
rect 145182 53442 145234 53454
rect 150782 53506 150834 53518
rect 150782 53442 150834 53454
rect 189422 53506 189474 53518
rect 189422 53442 189474 53454
rect 1344 53338 298592 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 81278 53338
rect 81330 53286 81382 53338
rect 81434 53286 81486 53338
rect 81538 53286 111998 53338
rect 112050 53286 112102 53338
rect 112154 53286 112206 53338
rect 112258 53286 142718 53338
rect 142770 53286 142822 53338
rect 142874 53286 142926 53338
rect 142978 53286 173438 53338
rect 173490 53286 173542 53338
rect 173594 53286 173646 53338
rect 173698 53286 204158 53338
rect 204210 53286 204262 53338
rect 204314 53286 204366 53338
rect 204418 53286 234878 53338
rect 234930 53286 234982 53338
rect 235034 53286 235086 53338
rect 235138 53286 265598 53338
rect 265650 53286 265702 53338
rect 265754 53286 265806 53338
rect 265858 53286 296318 53338
rect 296370 53286 296422 53338
rect 296474 53286 296526 53338
rect 296578 53286 298592 53338
rect 1344 53252 298592 53286
rect 182142 53170 182194 53182
rect 182142 53106 182194 53118
rect 185838 53170 185890 53182
rect 185838 53106 185890 53118
rect 182466 52894 182478 52946
rect 182530 52894 182542 52946
rect 186498 52894 186510 52946
rect 186562 52894 186574 52946
rect 181470 52834 181522 52846
rect 183250 52782 183262 52834
rect 183314 52782 183326 52834
rect 185378 52782 185390 52834
rect 185442 52782 185454 52834
rect 187170 52782 187182 52834
rect 187234 52782 187246 52834
rect 189298 52782 189310 52834
rect 189362 52782 189374 52834
rect 181470 52770 181522 52782
rect 1344 52554 298592 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 96638 52554
rect 96690 52502 96742 52554
rect 96794 52502 96846 52554
rect 96898 52502 127358 52554
rect 127410 52502 127462 52554
rect 127514 52502 127566 52554
rect 127618 52502 158078 52554
rect 158130 52502 158182 52554
rect 158234 52502 158286 52554
rect 158338 52502 188798 52554
rect 188850 52502 188902 52554
rect 188954 52502 189006 52554
rect 189058 52502 219518 52554
rect 219570 52502 219622 52554
rect 219674 52502 219726 52554
rect 219778 52502 250238 52554
rect 250290 52502 250342 52554
rect 250394 52502 250446 52554
rect 250498 52502 280958 52554
rect 281010 52502 281062 52554
rect 281114 52502 281166 52554
rect 281218 52502 298592 52554
rect 1344 52468 298592 52502
rect 186174 52274 186226 52286
rect 186174 52210 186226 52222
rect 1344 51770 298592 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 81278 51770
rect 81330 51718 81382 51770
rect 81434 51718 81486 51770
rect 81538 51718 111998 51770
rect 112050 51718 112102 51770
rect 112154 51718 112206 51770
rect 112258 51718 142718 51770
rect 142770 51718 142822 51770
rect 142874 51718 142926 51770
rect 142978 51718 173438 51770
rect 173490 51718 173542 51770
rect 173594 51718 173646 51770
rect 173698 51718 204158 51770
rect 204210 51718 204262 51770
rect 204314 51718 204366 51770
rect 204418 51718 234878 51770
rect 234930 51718 234982 51770
rect 235034 51718 235086 51770
rect 235138 51718 265598 51770
rect 265650 51718 265702 51770
rect 265754 51718 265806 51770
rect 265858 51718 296318 51770
rect 296370 51718 296422 51770
rect 296474 51718 296526 51770
rect 296578 51718 298592 51770
rect 1344 51684 298592 51718
rect 1344 50986 298592 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 96638 50986
rect 96690 50934 96742 50986
rect 96794 50934 96846 50986
rect 96898 50934 127358 50986
rect 127410 50934 127462 50986
rect 127514 50934 127566 50986
rect 127618 50934 158078 50986
rect 158130 50934 158182 50986
rect 158234 50934 158286 50986
rect 158338 50934 188798 50986
rect 188850 50934 188902 50986
rect 188954 50934 189006 50986
rect 189058 50934 219518 50986
rect 219570 50934 219622 50986
rect 219674 50934 219726 50986
rect 219778 50934 250238 50986
rect 250290 50934 250342 50986
rect 250394 50934 250446 50986
rect 250498 50934 280958 50986
rect 281010 50934 281062 50986
rect 281114 50934 281166 50986
rect 281218 50934 298592 50986
rect 1344 50900 298592 50934
rect 1344 50202 298592 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 81278 50202
rect 81330 50150 81382 50202
rect 81434 50150 81486 50202
rect 81538 50150 111998 50202
rect 112050 50150 112102 50202
rect 112154 50150 112206 50202
rect 112258 50150 142718 50202
rect 142770 50150 142822 50202
rect 142874 50150 142926 50202
rect 142978 50150 173438 50202
rect 173490 50150 173542 50202
rect 173594 50150 173646 50202
rect 173698 50150 204158 50202
rect 204210 50150 204262 50202
rect 204314 50150 204366 50202
rect 204418 50150 234878 50202
rect 234930 50150 234982 50202
rect 235034 50150 235086 50202
rect 235138 50150 265598 50202
rect 265650 50150 265702 50202
rect 265754 50150 265806 50202
rect 265858 50150 296318 50202
rect 296370 50150 296422 50202
rect 296474 50150 296526 50202
rect 296578 50150 298592 50202
rect 1344 50116 298592 50150
rect 1344 49418 298592 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 96638 49418
rect 96690 49366 96742 49418
rect 96794 49366 96846 49418
rect 96898 49366 127358 49418
rect 127410 49366 127462 49418
rect 127514 49366 127566 49418
rect 127618 49366 158078 49418
rect 158130 49366 158182 49418
rect 158234 49366 158286 49418
rect 158338 49366 188798 49418
rect 188850 49366 188902 49418
rect 188954 49366 189006 49418
rect 189058 49366 219518 49418
rect 219570 49366 219622 49418
rect 219674 49366 219726 49418
rect 219778 49366 250238 49418
rect 250290 49366 250342 49418
rect 250394 49366 250446 49418
rect 250498 49366 280958 49418
rect 281010 49366 281062 49418
rect 281114 49366 281166 49418
rect 281218 49366 298592 49418
rect 1344 49332 298592 49366
rect 1344 48634 298592 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 81278 48634
rect 81330 48582 81382 48634
rect 81434 48582 81486 48634
rect 81538 48582 111998 48634
rect 112050 48582 112102 48634
rect 112154 48582 112206 48634
rect 112258 48582 142718 48634
rect 142770 48582 142822 48634
rect 142874 48582 142926 48634
rect 142978 48582 173438 48634
rect 173490 48582 173542 48634
rect 173594 48582 173646 48634
rect 173698 48582 204158 48634
rect 204210 48582 204262 48634
rect 204314 48582 204366 48634
rect 204418 48582 234878 48634
rect 234930 48582 234982 48634
rect 235034 48582 235086 48634
rect 235138 48582 265598 48634
rect 265650 48582 265702 48634
rect 265754 48582 265806 48634
rect 265858 48582 296318 48634
rect 296370 48582 296422 48634
rect 296474 48582 296526 48634
rect 296578 48582 298592 48634
rect 1344 48548 298592 48582
rect 1344 47850 298592 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 96638 47850
rect 96690 47798 96742 47850
rect 96794 47798 96846 47850
rect 96898 47798 127358 47850
rect 127410 47798 127462 47850
rect 127514 47798 127566 47850
rect 127618 47798 158078 47850
rect 158130 47798 158182 47850
rect 158234 47798 158286 47850
rect 158338 47798 188798 47850
rect 188850 47798 188902 47850
rect 188954 47798 189006 47850
rect 189058 47798 219518 47850
rect 219570 47798 219622 47850
rect 219674 47798 219726 47850
rect 219778 47798 250238 47850
rect 250290 47798 250342 47850
rect 250394 47798 250446 47850
rect 250498 47798 280958 47850
rect 281010 47798 281062 47850
rect 281114 47798 281166 47850
rect 281218 47798 298592 47850
rect 1344 47764 298592 47798
rect 1344 47066 298592 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 81278 47066
rect 81330 47014 81382 47066
rect 81434 47014 81486 47066
rect 81538 47014 111998 47066
rect 112050 47014 112102 47066
rect 112154 47014 112206 47066
rect 112258 47014 142718 47066
rect 142770 47014 142822 47066
rect 142874 47014 142926 47066
rect 142978 47014 173438 47066
rect 173490 47014 173542 47066
rect 173594 47014 173646 47066
rect 173698 47014 204158 47066
rect 204210 47014 204262 47066
rect 204314 47014 204366 47066
rect 204418 47014 234878 47066
rect 234930 47014 234982 47066
rect 235034 47014 235086 47066
rect 235138 47014 265598 47066
rect 265650 47014 265702 47066
rect 265754 47014 265806 47066
rect 265858 47014 296318 47066
rect 296370 47014 296422 47066
rect 296474 47014 296526 47066
rect 296578 47014 298592 47066
rect 1344 46980 298592 47014
rect 1344 46282 298592 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 96638 46282
rect 96690 46230 96742 46282
rect 96794 46230 96846 46282
rect 96898 46230 127358 46282
rect 127410 46230 127462 46282
rect 127514 46230 127566 46282
rect 127618 46230 158078 46282
rect 158130 46230 158182 46282
rect 158234 46230 158286 46282
rect 158338 46230 188798 46282
rect 188850 46230 188902 46282
rect 188954 46230 189006 46282
rect 189058 46230 219518 46282
rect 219570 46230 219622 46282
rect 219674 46230 219726 46282
rect 219778 46230 250238 46282
rect 250290 46230 250342 46282
rect 250394 46230 250446 46282
rect 250498 46230 280958 46282
rect 281010 46230 281062 46282
rect 281114 46230 281166 46282
rect 281218 46230 298592 46282
rect 1344 46196 298592 46230
rect 1344 45498 298592 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 81278 45498
rect 81330 45446 81382 45498
rect 81434 45446 81486 45498
rect 81538 45446 111998 45498
rect 112050 45446 112102 45498
rect 112154 45446 112206 45498
rect 112258 45446 142718 45498
rect 142770 45446 142822 45498
rect 142874 45446 142926 45498
rect 142978 45446 173438 45498
rect 173490 45446 173542 45498
rect 173594 45446 173646 45498
rect 173698 45446 204158 45498
rect 204210 45446 204262 45498
rect 204314 45446 204366 45498
rect 204418 45446 234878 45498
rect 234930 45446 234982 45498
rect 235034 45446 235086 45498
rect 235138 45446 265598 45498
rect 265650 45446 265702 45498
rect 265754 45446 265806 45498
rect 265858 45446 296318 45498
rect 296370 45446 296422 45498
rect 296474 45446 296526 45498
rect 296578 45446 298592 45498
rect 1344 45412 298592 45446
rect 1344 44714 298592 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 96638 44714
rect 96690 44662 96742 44714
rect 96794 44662 96846 44714
rect 96898 44662 127358 44714
rect 127410 44662 127462 44714
rect 127514 44662 127566 44714
rect 127618 44662 158078 44714
rect 158130 44662 158182 44714
rect 158234 44662 158286 44714
rect 158338 44662 188798 44714
rect 188850 44662 188902 44714
rect 188954 44662 189006 44714
rect 189058 44662 219518 44714
rect 219570 44662 219622 44714
rect 219674 44662 219726 44714
rect 219778 44662 250238 44714
rect 250290 44662 250342 44714
rect 250394 44662 250446 44714
rect 250498 44662 280958 44714
rect 281010 44662 281062 44714
rect 281114 44662 281166 44714
rect 281218 44662 298592 44714
rect 1344 44628 298592 44662
rect 1344 43930 298592 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 81278 43930
rect 81330 43878 81382 43930
rect 81434 43878 81486 43930
rect 81538 43878 111998 43930
rect 112050 43878 112102 43930
rect 112154 43878 112206 43930
rect 112258 43878 142718 43930
rect 142770 43878 142822 43930
rect 142874 43878 142926 43930
rect 142978 43878 173438 43930
rect 173490 43878 173542 43930
rect 173594 43878 173646 43930
rect 173698 43878 204158 43930
rect 204210 43878 204262 43930
rect 204314 43878 204366 43930
rect 204418 43878 234878 43930
rect 234930 43878 234982 43930
rect 235034 43878 235086 43930
rect 235138 43878 265598 43930
rect 265650 43878 265702 43930
rect 265754 43878 265806 43930
rect 265858 43878 296318 43930
rect 296370 43878 296422 43930
rect 296474 43878 296526 43930
rect 296578 43878 298592 43930
rect 1344 43844 298592 43878
rect 1344 43146 298592 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 96638 43146
rect 96690 43094 96742 43146
rect 96794 43094 96846 43146
rect 96898 43094 127358 43146
rect 127410 43094 127462 43146
rect 127514 43094 127566 43146
rect 127618 43094 158078 43146
rect 158130 43094 158182 43146
rect 158234 43094 158286 43146
rect 158338 43094 188798 43146
rect 188850 43094 188902 43146
rect 188954 43094 189006 43146
rect 189058 43094 219518 43146
rect 219570 43094 219622 43146
rect 219674 43094 219726 43146
rect 219778 43094 250238 43146
rect 250290 43094 250342 43146
rect 250394 43094 250446 43146
rect 250498 43094 280958 43146
rect 281010 43094 281062 43146
rect 281114 43094 281166 43146
rect 281218 43094 298592 43146
rect 1344 43060 298592 43094
rect 1344 42362 298592 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 81278 42362
rect 81330 42310 81382 42362
rect 81434 42310 81486 42362
rect 81538 42310 111998 42362
rect 112050 42310 112102 42362
rect 112154 42310 112206 42362
rect 112258 42310 142718 42362
rect 142770 42310 142822 42362
rect 142874 42310 142926 42362
rect 142978 42310 173438 42362
rect 173490 42310 173542 42362
rect 173594 42310 173646 42362
rect 173698 42310 204158 42362
rect 204210 42310 204262 42362
rect 204314 42310 204366 42362
rect 204418 42310 234878 42362
rect 234930 42310 234982 42362
rect 235034 42310 235086 42362
rect 235138 42310 265598 42362
rect 265650 42310 265702 42362
rect 265754 42310 265806 42362
rect 265858 42310 296318 42362
rect 296370 42310 296422 42362
rect 296474 42310 296526 42362
rect 296578 42310 298592 42362
rect 1344 42276 298592 42310
rect 1344 41578 298592 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 96638 41578
rect 96690 41526 96742 41578
rect 96794 41526 96846 41578
rect 96898 41526 127358 41578
rect 127410 41526 127462 41578
rect 127514 41526 127566 41578
rect 127618 41526 158078 41578
rect 158130 41526 158182 41578
rect 158234 41526 158286 41578
rect 158338 41526 188798 41578
rect 188850 41526 188902 41578
rect 188954 41526 189006 41578
rect 189058 41526 219518 41578
rect 219570 41526 219622 41578
rect 219674 41526 219726 41578
rect 219778 41526 250238 41578
rect 250290 41526 250342 41578
rect 250394 41526 250446 41578
rect 250498 41526 280958 41578
rect 281010 41526 281062 41578
rect 281114 41526 281166 41578
rect 281218 41526 298592 41578
rect 1344 41492 298592 41526
rect 1344 40794 298592 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 81278 40794
rect 81330 40742 81382 40794
rect 81434 40742 81486 40794
rect 81538 40742 111998 40794
rect 112050 40742 112102 40794
rect 112154 40742 112206 40794
rect 112258 40742 142718 40794
rect 142770 40742 142822 40794
rect 142874 40742 142926 40794
rect 142978 40742 173438 40794
rect 173490 40742 173542 40794
rect 173594 40742 173646 40794
rect 173698 40742 204158 40794
rect 204210 40742 204262 40794
rect 204314 40742 204366 40794
rect 204418 40742 234878 40794
rect 234930 40742 234982 40794
rect 235034 40742 235086 40794
rect 235138 40742 265598 40794
rect 265650 40742 265702 40794
rect 265754 40742 265806 40794
rect 265858 40742 296318 40794
rect 296370 40742 296422 40794
rect 296474 40742 296526 40794
rect 296578 40742 298592 40794
rect 1344 40708 298592 40742
rect 1344 40010 298592 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 96638 40010
rect 96690 39958 96742 40010
rect 96794 39958 96846 40010
rect 96898 39958 127358 40010
rect 127410 39958 127462 40010
rect 127514 39958 127566 40010
rect 127618 39958 158078 40010
rect 158130 39958 158182 40010
rect 158234 39958 158286 40010
rect 158338 39958 188798 40010
rect 188850 39958 188902 40010
rect 188954 39958 189006 40010
rect 189058 39958 219518 40010
rect 219570 39958 219622 40010
rect 219674 39958 219726 40010
rect 219778 39958 250238 40010
rect 250290 39958 250342 40010
rect 250394 39958 250446 40010
rect 250498 39958 280958 40010
rect 281010 39958 281062 40010
rect 281114 39958 281166 40010
rect 281218 39958 298592 40010
rect 1344 39924 298592 39958
rect 1344 39226 298592 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 81278 39226
rect 81330 39174 81382 39226
rect 81434 39174 81486 39226
rect 81538 39174 111998 39226
rect 112050 39174 112102 39226
rect 112154 39174 112206 39226
rect 112258 39174 142718 39226
rect 142770 39174 142822 39226
rect 142874 39174 142926 39226
rect 142978 39174 173438 39226
rect 173490 39174 173542 39226
rect 173594 39174 173646 39226
rect 173698 39174 204158 39226
rect 204210 39174 204262 39226
rect 204314 39174 204366 39226
rect 204418 39174 234878 39226
rect 234930 39174 234982 39226
rect 235034 39174 235086 39226
rect 235138 39174 265598 39226
rect 265650 39174 265702 39226
rect 265754 39174 265806 39226
rect 265858 39174 296318 39226
rect 296370 39174 296422 39226
rect 296474 39174 296526 39226
rect 296578 39174 298592 39226
rect 1344 39140 298592 39174
rect 1344 38442 298592 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 96638 38442
rect 96690 38390 96742 38442
rect 96794 38390 96846 38442
rect 96898 38390 127358 38442
rect 127410 38390 127462 38442
rect 127514 38390 127566 38442
rect 127618 38390 158078 38442
rect 158130 38390 158182 38442
rect 158234 38390 158286 38442
rect 158338 38390 188798 38442
rect 188850 38390 188902 38442
rect 188954 38390 189006 38442
rect 189058 38390 219518 38442
rect 219570 38390 219622 38442
rect 219674 38390 219726 38442
rect 219778 38390 250238 38442
rect 250290 38390 250342 38442
rect 250394 38390 250446 38442
rect 250498 38390 280958 38442
rect 281010 38390 281062 38442
rect 281114 38390 281166 38442
rect 281218 38390 298592 38442
rect 1344 38356 298592 38390
rect 1344 37658 298592 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 81278 37658
rect 81330 37606 81382 37658
rect 81434 37606 81486 37658
rect 81538 37606 111998 37658
rect 112050 37606 112102 37658
rect 112154 37606 112206 37658
rect 112258 37606 142718 37658
rect 142770 37606 142822 37658
rect 142874 37606 142926 37658
rect 142978 37606 173438 37658
rect 173490 37606 173542 37658
rect 173594 37606 173646 37658
rect 173698 37606 204158 37658
rect 204210 37606 204262 37658
rect 204314 37606 204366 37658
rect 204418 37606 234878 37658
rect 234930 37606 234982 37658
rect 235034 37606 235086 37658
rect 235138 37606 265598 37658
rect 265650 37606 265702 37658
rect 265754 37606 265806 37658
rect 265858 37606 296318 37658
rect 296370 37606 296422 37658
rect 296474 37606 296526 37658
rect 296578 37606 298592 37658
rect 1344 37572 298592 37606
rect 1344 36874 298592 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 96638 36874
rect 96690 36822 96742 36874
rect 96794 36822 96846 36874
rect 96898 36822 127358 36874
rect 127410 36822 127462 36874
rect 127514 36822 127566 36874
rect 127618 36822 158078 36874
rect 158130 36822 158182 36874
rect 158234 36822 158286 36874
rect 158338 36822 188798 36874
rect 188850 36822 188902 36874
rect 188954 36822 189006 36874
rect 189058 36822 219518 36874
rect 219570 36822 219622 36874
rect 219674 36822 219726 36874
rect 219778 36822 250238 36874
rect 250290 36822 250342 36874
rect 250394 36822 250446 36874
rect 250498 36822 280958 36874
rect 281010 36822 281062 36874
rect 281114 36822 281166 36874
rect 281218 36822 298592 36874
rect 1344 36788 298592 36822
rect 1344 36090 298592 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 81278 36090
rect 81330 36038 81382 36090
rect 81434 36038 81486 36090
rect 81538 36038 111998 36090
rect 112050 36038 112102 36090
rect 112154 36038 112206 36090
rect 112258 36038 142718 36090
rect 142770 36038 142822 36090
rect 142874 36038 142926 36090
rect 142978 36038 173438 36090
rect 173490 36038 173542 36090
rect 173594 36038 173646 36090
rect 173698 36038 204158 36090
rect 204210 36038 204262 36090
rect 204314 36038 204366 36090
rect 204418 36038 234878 36090
rect 234930 36038 234982 36090
rect 235034 36038 235086 36090
rect 235138 36038 265598 36090
rect 265650 36038 265702 36090
rect 265754 36038 265806 36090
rect 265858 36038 296318 36090
rect 296370 36038 296422 36090
rect 296474 36038 296526 36090
rect 296578 36038 298592 36090
rect 1344 36004 298592 36038
rect 1344 35306 298592 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 96638 35306
rect 96690 35254 96742 35306
rect 96794 35254 96846 35306
rect 96898 35254 127358 35306
rect 127410 35254 127462 35306
rect 127514 35254 127566 35306
rect 127618 35254 158078 35306
rect 158130 35254 158182 35306
rect 158234 35254 158286 35306
rect 158338 35254 188798 35306
rect 188850 35254 188902 35306
rect 188954 35254 189006 35306
rect 189058 35254 219518 35306
rect 219570 35254 219622 35306
rect 219674 35254 219726 35306
rect 219778 35254 250238 35306
rect 250290 35254 250342 35306
rect 250394 35254 250446 35306
rect 250498 35254 280958 35306
rect 281010 35254 281062 35306
rect 281114 35254 281166 35306
rect 281218 35254 298592 35306
rect 1344 35220 298592 35254
rect 1344 34522 298592 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 81278 34522
rect 81330 34470 81382 34522
rect 81434 34470 81486 34522
rect 81538 34470 111998 34522
rect 112050 34470 112102 34522
rect 112154 34470 112206 34522
rect 112258 34470 142718 34522
rect 142770 34470 142822 34522
rect 142874 34470 142926 34522
rect 142978 34470 173438 34522
rect 173490 34470 173542 34522
rect 173594 34470 173646 34522
rect 173698 34470 204158 34522
rect 204210 34470 204262 34522
rect 204314 34470 204366 34522
rect 204418 34470 234878 34522
rect 234930 34470 234982 34522
rect 235034 34470 235086 34522
rect 235138 34470 265598 34522
rect 265650 34470 265702 34522
rect 265754 34470 265806 34522
rect 265858 34470 296318 34522
rect 296370 34470 296422 34522
rect 296474 34470 296526 34522
rect 296578 34470 298592 34522
rect 1344 34436 298592 34470
rect 1344 33738 298592 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 96638 33738
rect 96690 33686 96742 33738
rect 96794 33686 96846 33738
rect 96898 33686 127358 33738
rect 127410 33686 127462 33738
rect 127514 33686 127566 33738
rect 127618 33686 158078 33738
rect 158130 33686 158182 33738
rect 158234 33686 158286 33738
rect 158338 33686 188798 33738
rect 188850 33686 188902 33738
rect 188954 33686 189006 33738
rect 189058 33686 219518 33738
rect 219570 33686 219622 33738
rect 219674 33686 219726 33738
rect 219778 33686 250238 33738
rect 250290 33686 250342 33738
rect 250394 33686 250446 33738
rect 250498 33686 280958 33738
rect 281010 33686 281062 33738
rect 281114 33686 281166 33738
rect 281218 33686 298592 33738
rect 1344 33652 298592 33686
rect 1344 32954 298592 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 81278 32954
rect 81330 32902 81382 32954
rect 81434 32902 81486 32954
rect 81538 32902 111998 32954
rect 112050 32902 112102 32954
rect 112154 32902 112206 32954
rect 112258 32902 142718 32954
rect 142770 32902 142822 32954
rect 142874 32902 142926 32954
rect 142978 32902 173438 32954
rect 173490 32902 173542 32954
rect 173594 32902 173646 32954
rect 173698 32902 204158 32954
rect 204210 32902 204262 32954
rect 204314 32902 204366 32954
rect 204418 32902 234878 32954
rect 234930 32902 234982 32954
rect 235034 32902 235086 32954
rect 235138 32902 265598 32954
rect 265650 32902 265702 32954
rect 265754 32902 265806 32954
rect 265858 32902 296318 32954
rect 296370 32902 296422 32954
rect 296474 32902 296526 32954
rect 296578 32902 298592 32954
rect 1344 32868 298592 32902
rect 1344 32170 298592 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 96638 32170
rect 96690 32118 96742 32170
rect 96794 32118 96846 32170
rect 96898 32118 127358 32170
rect 127410 32118 127462 32170
rect 127514 32118 127566 32170
rect 127618 32118 158078 32170
rect 158130 32118 158182 32170
rect 158234 32118 158286 32170
rect 158338 32118 188798 32170
rect 188850 32118 188902 32170
rect 188954 32118 189006 32170
rect 189058 32118 219518 32170
rect 219570 32118 219622 32170
rect 219674 32118 219726 32170
rect 219778 32118 250238 32170
rect 250290 32118 250342 32170
rect 250394 32118 250446 32170
rect 250498 32118 280958 32170
rect 281010 32118 281062 32170
rect 281114 32118 281166 32170
rect 281218 32118 298592 32170
rect 1344 32084 298592 32118
rect 1344 31386 298592 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 81278 31386
rect 81330 31334 81382 31386
rect 81434 31334 81486 31386
rect 81538 31334 111998 31386
rect 112050 31334 112102 31386
rect 112154 31334 112206 31386
rect 112258 31334 142718 31386
rect 142770 31334 142822 31386
rect 142874 31334 142926 31386
rect 142978 31334 173438 31386
rect 173490 31334 173542 31386
rect 173594 31334 173646 31386
rect 173698 31334 204158 31386
rect 204210 31334 204262 31386
rect 204314 31334 204366 31386
rect 204418 31334 234878 31386
rect 234930 31334 234982 31386
rect 235034 31334 235086 31386
rect 235138 31334 265598 31386
rect 265650 31334 265702 31386
rect 265754 31334 265806 31386
rect 265858 31334 296318 31386
rect 296370 31334 296422 31386
rect 296474 31334 296526 31386
rect 296578 31334 298592 31386
rect 1344 31300 298592 31334
rect 1344 30602 298592 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 96638 30602
rect 96690 30550 96742 30602
rect 96794 30550 96846 30602
rect 96898 30550 127358 30602
rect 127410 30550 127462 30602
rect 127514 30550 127566 30602
rect 127618 30550 158078 30602
rect 158130 30550 158182 30602
rect 158234 30550 158286 30602
rect 158338 30550 188798 30602
rect 188850 30550 188902 30602
rect 188954 30550 189006 30602
rect 189058 30550 219518 30602
rect 219570 30550 219622 30602
rect 219674 30550 219726 30602
rect 219778 30550 250238 30602
rect 250290 30550 250342 30602
rect 250394 30550 250446 30602
rect 250498 30550 280958 30602
rect 281010 30550 281062 30602
rect 281114 30550 281166 30602
rect 281218 30550 298592 30602
rect 1344 30516 298592 30550
rect 1344 29818 298592 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 81278 29818
rect 81330 29766 81382 29818
rect 81434 29766 81486 29818
rect 81538 29766 111998 29818
rect 112050 29766 112102 29818
rect 112154 29766 112206 29818
rect 112258 29766 142718 29818
rect 142770 29766 142822 29818
rect 142874 29766 142926 29818
rect 142978 29766 173438 29818
rect 173490 29766 173542 29818
rect 173594 29766 173646 29818
rect 173698 29766 204158 29818
rect 204210 29766 204262 29818
rect 204314 29766 204366 29818
rect 204418 29766 234878 29818
rect 234930 29766 234982 29818
rect 235034 29766 235086 29818
rect 235138 29766 265598 29818
rect 265650 29766 265702 29818
rect 265754 29766 265806 29818
rect 265858 29766 296318 29818
rect 296370 29766 296422 29818
rect 296474 29766 296526 29818
rect 296578 29766 298592 29818
rect 1344 29732 298592 29766
rect 1344 29034 298592 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 96638 29034
rect 96690 28982 96742 29034
rect 96794 28982 96846 29034
rect 96898 28982 127358 29034
rect 127410 28982 127462 29034
rect 127514 28982 127566 29034
rect 127618 28982 158078 29034
rect 158130 28982 158182 29034
rect 158234 28982 158286 29034
rect 158338 28982 188798 29034
rect 188850 28982 188902 29034
rect 188954 28982 189006 29034
rect 189058 28982 219518 29034
rect 219570 28982 219622 29034
rect 219674 28982 219726 29034
rect 219778 28982 250238 29034
rect 250290 28982 250342 29034
rect 250394 28982 250446 29034
rect 250498 28982 280958 29034
rect 281010 28982 281062 29034
rect 281114 28982 281166 29034
rect 281218 28982 298592 29034
rect 1344 28948 298592 28982
rect 1344 28250 298592 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 81278 28250
rect 81330 28198 81382 28250
rect 81434 28198 81486 28250
rect 81538 28198 111998 28250
rect 112050 28198 112102 28250
rect 112154 28198 112206 28250
rect 112258 28198 142718 28250
rect 142770 28198 142822 28250
rect 142874 28198 142926 28250
rect 142978 28198 173438 28250
rect 173490 28198 173542 28250
rect 173594 28198 173646 28250
rect 173698 28198 204158 28250
rect 204210 28198 204262 28250
rect 204314 28198 204366 28250
rect 204418 28198 234878 28250
rect 234930 28198 234982 28250
rect 235034 28198 235086 28250
rect 235138 28198 265598 28250
rect 265650 28198 265702 28250
rect 265754 28198 265806 28250
rect 265858 28198 296318 28250
rect 296370 28198 296422 28250
rect 296474 28198 296526 28250
rect 296578 28198 298592 28250
rect 1344 28164 298592 28198
rect 1344 27466 298592 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 96638 27466
rect 96690 27414 96742 27466
rect 96794 27414 96846 27466
rect 96898 27414 127358 27466
rect 127410 27414 127462 27466
rect 127514 27414 127566 27466
rect 127618 27414 158078 27466
rect 158130 27414 158182 27466
rect 158234 27414 158286 27466
rect 158338 27414 188798 27466
rect 188850 27414 188902 27466
rect 188954 27414 189006 27466
rect 189058 27414 219518 27466
rect 219570 27414 219622 27466
rect 219674 27414 219726 27466
rect 219778 27414 250238 27466
rect 250290 27414 250342 27466
rect 250394 27414 250446 27466
rect 250498 27414 280958 27466
rect 281010 27414 281062 27466
rect 281114 27414 281166 27466
rect 281218 27414 298592 27466
rect 1344 27380 298592 27414
rect 1344 26682 298592 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 81278 26682
rect 81330 26630 81382 26682
rect 81434 26630 81486 26682
rect 81538 26630 111998 26682
rect 112050 26630 112102 26682
rect 112154 26630 112206 26682
rect 112258 26630 142718 26682
rect 142770 26630 142822 26682
rect 142874 26630 142926 26682
rect 142978 26630 173438 26682
rect 173490 26630 173542 26682
rect 173594 26630 173646 26682
rect 173698 26630 204158 26682
rect 204210 26630 204262 26682
rect 204314 26630 204366 26682
rect 204418 26630 234878 26682
rect 234930 26630 234982 26682
rect 235034 26630 235086 26682
rect 235138 26630 265598 26682
rect 265650 26630 265702 26682
rect 265754 26630 265806 26682
rect 265858 26630 296318 26682
rect 296370 26630 296422 26682
rect 296474 26630 296526 26682
rect 296578 26630 298592 26682
rect 1344 26596 298592 26630
rect 1344 25898 298592 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 96638 25898
rect 96690 25846 96742 25898
rect 96794 25846 96846 25898
rect 96898 25846 127358 25898
rect 127410 25846 127462 25898
rect 127514 25846 127566 25898
rect 127618 25846 158078 25898
rect 158130 25846 158182 25898
rect 158234 25846 158286 25898
rect 158338 25846 188798 25898
rect 188850 25846 188902 25898
rect 188954 25846 189006 25898
rect 189058 25846 219518 25898
rect 219570 25846 219622 25898
rect 219674 25846 219726 25898
rect 219778 25846 250238 25898
rect 250290 25846 250342 25898
rect 250394 25846 250446 25898
rect 250498 25846 280958 25898
rect 281010 25846 281062 25898
rect 281114 25846 281166 25898
rect 281218 25846 298592 25898
rect 1344 25812 298592 25846
rect 1344 25114 298592 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 81278 25114
rect 81330 25062 81382 25114
rect 81434 25062 81486 25114
rect 81538 25062 111998 25114
rect 112050 25062 112102 25114
rect 112154 25062 112206 25114
rect 112258 25062 142718 25114
rect 142770 25062 142822 25114
rect 142874 25062 142926 25114
rect 142978 25062 173438 25114
rect 173490 25062 173542 25114
rect 173594 25062 173646 25114
rect 173698 25062 204158 25114
rect 204210 25062 204262 25114
rect 204314 25062 204366 25114
rect 204418 25062 234878 25114
rect 234930 25062 234982 25114
rect 235034 25062 235086 25114
rect 235138 25062 265598 25114
rect 265650 25062 265702 25114
rect 265754 25062 265806 25114
rect 265858 25062 296318 25114
rect 296370 25062 296422 25114
rect 296474 25062 296526 25114
rect 296578 25062 298592 25114
rect 1344 25028 298592 25062
rect 1344 24330 298592 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 96638 24330
rect 96690 24278 96742 24330
rect 96794 24278 96846 24330
rect 96898 24278 127358 24330
rect 127410 24278 127462 24330
rect 127514 24278 127566 24330
rect 127618 24278 158078 24330
rect 158130 24278 158182 24330
rect 158234 24278 158286 24330
rect 158338 24278 188798 24330
rect 188850 24278 188902 24330
rect 188954 24278 189006 24330
rect 189058 24278 219518 24330
rect 219570 24278 219622 24330
rect 219674 24278 219726 24330
rect 219778 24278 250238 24330
rect 250290 24278 250342 24330
rect 250394 24278 250446 24330
rect 250498 24278 280958 24330
rect 281010 24278 281062 24330
rect 281114 24278 281166 24330
rect 281218 24278 298592 24330
rect 1344 24244 298592 24278
rect 1344 23546 298592 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 81278 23546
rect 81330 23494 81382 23546
rect 81434 23494 81486 23546
rect 81538 23494 111998 23546
rect 112050 23494 112102 23546
rect 112154 23494 112206 23546
rect 112258 23494 142718 23546
rect 142770 23494 142822 23546
rect 142874 23494 142926 23546
rect 142978 23494 173438 23546
rect 173490 23494 173542 23546
rect 173594 23494 173646 23546
rect 173698 23494 204158 23546
rect 204210 23494 204262 23546
rect 204314 23494 204366 23546
rect 204418 23494 234878 23546
rect 234930 23494 234982 23546
rect 235034 23494 235086 23546
rect 235138 23494 265598 23546
rect 265650 23494 265702 23546
rect 265754 23494 265806 23546
rect 265858 23494 296318 23546
rect 296370 23494 296422 23546
rect 296474 23494 296526 23546
rect 296578 23494 298592 23546
rect 1344 23460 298592 23494
rect 1344 22762 298592 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 96638 22762
rect 96690 22710 96742 22762
rect 96794 22710 96846 22762
rect 96898 22710 127358 22762
rect 127410 22710 127462 22762
rect 127514 22710 127566 22762
rect 127618 22710 158078 22762
rect 158130 22710 158182 22762
rect 158234 22710 158286 22762
rect 158338 22710 188798 22762
rect 188850 22710 188902 22762
rect 188954 22710 189006 22762
rect 189058 22710 219518 22762
rect 219570 22710 219622 22762
rect 219674 22710 219726 22762
rect 219778 22710 250238 22762
rect 250290 22710 250342 22762
rect 250394 22710 250446 22762
rect 250498 22710 280958 22762
rect 281010 22710 281062 22762
rect 281114 22710 281166 22762
rect 281218 22710 298592 22762
rect 1344 22676 298592 22710
rect 1344 21978 298592 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 81278 21978
rect 81330 21926 81382 21978
rect 81434 21926 81486 21978
rect 81538 21926 111998 21978
rect 112050 21926 112102 21978
rect 112154 21926 112206 21978
rect 112258 21926 142718 21978
rect 142770 21926 142822 21978
rect 142874 21926 142926 21978
rect 142978 21926 173438 21978
rect 173490 21926 173542 21978
rect 173594 21926 173646 21978
rect 173698 21926 204158 21978
rect 204210 21926 204262 21978
rect 204314 21926 204366 21978
rect 204418 21926 234878 21978
rect 234930 21926 234982 21978
rect 235034 21926 235086 21978
rect 235138 21926 265598 21978
rect 265650 21926 265702 21978
rect 265754 21926 265806 21978
rect 265858 21926 296318 21978
rect 296370 21926 296422 21978
rect 296474 21926 296526 21978
rect 296578 21926 298592 21978
rect 1344 21892 298592 21926
rect 1344 21194 298592 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 96638 21194
rect 96690 21142 96742 21194
rect 96794 21142 96846 21194
rect 96898 21142 127358 21194
rect 127410 21142 127462 21194
rect 127514 21142 127566 21194
rect 127618 21142 158078 21194
rect 158130 21142 158182 21194
rect 158234 21142 158286 21194
rect 158338 21142 188798 21194
rect 188850 21142 188902 21194
rect 188954 21142 189006 21194
rect 189058 21142 219518 21194
rect 219570 21142 219622 21194
rect 219674 21142 219726 21194
rect 219778 21142 250238 21194
rect 250290 21142 250342 21194
rect 250394 21142 250446 21194
rect 250498 21142 280958 21194
rect 281010 21142 281062 21194
rect 281114 21142 281166 21194
rect 281218 21142 298592 21194
rect 1344 21108 298592 21142
rect 1344 20410 298592 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 81278 20410
rect 81330 20358 81382 20410
rect 81434 20358 81486 20410
rect 81538 20358 111998 20410
rect 112050 20358 112102 20410
rect 112154 20358 112206 20410
rect 112258 20358 142718 20410
rect 142770 20358 142822 20410
rect 142874 20358 142926 20410
rect 142978 20358 173438 20410
rect 173490 20358 173542 20410
rect 173594 20358 173646 20410
rect 173698 20358 204158 20410
rect 204210 20358 204262 20410
rect 204314 20358 204366 20410
rect 204418 20358 234878 20410
rect 234930 20358 234982 20410
rect 235034 20358 235086 20410
rect 235138 20358 265598 20410
rect 265650 20358 265702 20410
rect 265754 20358 265806 20410
rect 265858 20358 296318 20410
rect 296370 20358 296422 20410
rect 296474 20358 296526 20410
rect 296578 20358 298592 20410
rect 1344 20324 298592 20358
rect 1344 19626 298592 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 96638 19626
rect 96690 19574 96742 19626
rect 96794 19574 96846 19626
rect 96898 19574 127358 19626
rect 127410 19574 127462 19626
rect 127514 19574 127566 19626
rect 127618 19574 158078 19626
rect 158130 19574 158182 19626
rect 158234 19574 158286 19626
rect 158338 19574 188798 19626
rect 188850 19574 188902 19626
rect 188954 19574 189006 19626
rect 189058 19574 219518 19626
rect 219570 19574 219622 19626
rect 219674 19574 219726 19626
rect 219778 19574 250238 19626
rect 250290 19574 250342 19626
rect 250394 19574 250446 19626
rect 250498 19574 280958 19626
rect 281010 19574 281062 19626
rect 281114 19574 281166 19626
rect 281218 19574 298592 19626
rect 1344 19540 298592 19574
rect 1344 18842 298592 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 81278 18842
rect 81330 18790 81382 18842
rect 81434 18790 81486 18842
rect 81538 18790 111998 18842
rect 112050 18790 112102 18842
rect 112154 18790 112206 18842
rect 112258 18790 142718 18842
rect 142770 18790 142822 18842
rect 142874 18790 142926 18842
rect 142978 18790 173438 18842
rect 173490 18790 173542 18842
rect 173594 18790 173646 18842
rect 173698 18790 204158 18842
rect 204210 18790 204262 18842
rect 204314 18790 204366 18842
rect 204418 18790 234878 18842
rect 234930 18790 234982 18842
rect 235034 18790 235086 18842
rect 235138 18790 265598 18842
rect 265650 18790 265702 18842
rect 265754 18790 265806 18842
rect 265858 18790 296318 18842
rect 296370 18790 296422 18842
rect 296474 18790 296526 18842
rect 296578 18790 298592 18842
rect 1344 18756 298592 18790
rect 1344 18058 298592 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 96638 18058
rect 96690 18006 96742 18058
rect 96794 18006 96846 18058
rect 96898 18006 127358 18058
rect 127410 18006 127462 18058
rect 127514 18006 127566 18058
rect 127618 18006 158078 18058
rect 158130 18006 158182 18058
rect 158234 18006 158286 18058
rect 158338 18006 188798 18058
rect 188850 18006 188902 18058
rect 188954 18006 189006 18058
rect 189058 18006 219518 18058
rect 219570 18006 219622 18058
rect 219674 18006 219726 18058
rect 219778 18006 250238 18058
rect 250290 18006 250342 18058
rect 250394 18006 250446 18058
rect 250498 18006 280958 18058
rect 281010 18006 281062 18058
rect 281114 18006 281166 18058
rect 281218 18006 298592 18058
rect 1344 17972 298592 18006
rect 1344 17274 298592 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 81278 17274
rect 81330 17222 81382 17274
rect 81434 17222 81486 17274
rect 81538 17222 111998 17274
rect 112050 17222 112102 17274
rect 112154 17222 112206 17274
rect 112258 17222 142718 17274
rect 142770 17222 142822 17274
rect 142874 17222 142926 17274
rect 142978 17222 173438 17274
rect 173490 17222 173542 17274
rect 173594 17222 173646 17274
rect 173698 17222 204158 17274
rect 204210 17222 204262 17274
rect 204314 17222 204366 17274
rect 204418 17222 234878 17274
rect 234930 17222 234982 17274
rect 235034 17222 235086 17274
rect 235138 17222 265598 17274
rect 265650 17222 265702 17274
rect 265754 17222 265806 17274
rect 265858 17222 296318 17274
rect 296370 17222 296422 17274
rect 296474 17222 296526 17274
rect 296578 17222 298592 17274
rect 1344 17188 298592 17222
rect 1344 16490 298592 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 96638 16490
rect 96690 16438 96742 16490
rect 96794 16438 96846 16490
rect 96898 16438 127358 16490
rect 127410 16438 127462 16490
rect 127514 16438 127566 16490
rect 127618 16438 158078 16490
rect 158130 16438 158182 16490
rect 158234 16438 158286 16490
rect 158338 16438 188798 16490
rect 188850 16438 188902 16490
rect 188954 16438 189006 16490
rect 189058 16438 219518 16490
rect 219570 16438 219622 16490
rect 219674 16438 219726 16490
rect 219778 16438 250238 16490
rect 250290 16438 250342 16490
rect 250394 16438 250446 16490
rect 250498 16438 280958 16490
rect 281010 16438 281062 16490
rect 281114 16438 281166 16490
rect 281218 16438 298592 16490
rect 1344 16404 298592 16438
rect 1344 15706 298592 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 81278 15706
rect 81330 15654 81382 15706
rect 81434 15654 81486 15706
rect 81538 15654 111998 15706
rect 112050 15654 112102 15706
rect 112154 15654 112206 15706
rect 112258 15654 142718 15706
rect 142770 15654 142822 15706
rect 142874 15654 142926 15706
rect 142978 15654 173438 15706
rect 173490 15654 173542 15706
rect 173594 15654 173646 15706
rect 173698 15654 204158 15706
rect 204210 15654 204262 15706
rect 204314 15654 204366 15706
rect 204418 15654 234878 15706
rect 234930 15654 234982 15706
rect 235034 15654 235086 15706
rect 235138 15654 265598 15706
rect 265650 15654 265702 15706
rect 265754 15654 265806 15706
rect 265858 15654 296318 15706
rect 296370 15654 296422 15706
rect 296474 15654 296526 15706
rect 296578 15654 298592 15706
rect 1344 15620 298592 15654
rect 1344 14922 298592 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 96638 14922
rect 96690 14870 96742 14922
rect 96794 14870 96846 14922
rect 96898 14870 127358 14922
rect 127410 14870 127462 14922
rect 127514 14870 127566 14922
rect 127618 14870 158078 14922
rect 158130 14870 158182 14922
rect 158234 14870 158286 14922
rect 158338 14870 188798 14922
rect 188850 14870 188902 14922
rect 188954 14870 189006 14922
rect 189058 14870 219518 14922
rect 219570 14870 219622 14922
rect 219674 14870 219726 14922
rect 219778 14870 250238 14922
rect 250290 14870 250342 14922
rect 250394 14870 250446 14922
rect 250498 14870 280958 14922
rect 281010 14870 281062 14922
rect 281114 14870 281166 14922
rect 281218 14870 298592 14922
rect 1344 14836 298592 14870
rect 1344 14138 298592 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 81278 14138
rect 81330 14086 81382 14138
rect 81434 14086 81486 14138
rect 81538 14086 111998 14138
rect 112050 14086 112102 14138
rect 112154 14086 112206 14138
rect 112258 14086 142718 14138
rect 142770 14086 142822 14138
rect 142874 14086 142926 14138
rect 142978 14086 173438 14138
rect 173490 14086 173542 14138
rect 173594 14086 173646 14138
rect 173698 14086 204158 14138
rect 204210 14086 204262 14138
rect 204314 14086 204366 14138
rect 204418 14086 234878 14138
rect 234930 14086 234982 14138
rect 235034 14086 235086 14138
rect 235138 14086 265598 14138
rect 265650 14086 265702 14138
rect 265754 14086 265806 14138
rect 265858 14086 296318 14138
rect 296370 14086 296422 14138
rect 296474 14086 296526 14138
rect 296578 14086 298592 14138
rect 1344 14052 298592 14086
rect 1344 13354 298592 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 96638 13354
rect 96690 13302 96742 13354
rect 96794 13302 96846 13354
rect 96898 13302 127358 13354
rect 127410 13302 127462 13354
rect 127514 13302 127566 13354
rect 127618 13302 158078 13354
rect 158130 13302 158182 13354
rect 158234 13302 158286 13354
rect 158338 13302 188798 13354
rect 188850 13302 188902 13354
rect 188954 13302 189006 13354
rect 189058 13302 219518 13354
rect 219570 13302 219622 13354
rect 219674 13302 219726 13354
rect 219778 13302 250238 13354
rect 250290 13302 250342 13354
rect 250394 13302 250446 13354
rect 250498 13302 280958 13354
rect 281010 13302 281062 13354
rect 281114 13302 281166 13354
rect 281218 13302 298592 13354
rect 1344 13268 298592 13302
rect 1344 12570 298592 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 81278 12570
rect 81330 12518 81382 12570
rect 81434 12518 81486 12570
rect 81538 12518 111998 12570
rect 112050 12518 112102 12570
rect 112154 12518 112206 12570
rect 112258 12518 142718 12570
rect 142770 12518 142822 12570
rect 142874 12518 142926 12570
rect 142978 12518 173438 12570
rect 173490 12518 173542 12570
rect 173594 12518 173646 12570
rect 173698 12518 204158 12570
rect 204210 12518 204262 12570
rect 204314 12518 204366 12570
rect 204418 12518 234878 12570
rect 234930 12518 234982 12570
rect 235034 12518 235086 12570
rect 235138 12518 265598 12570
rect 265650 12518 265702 12570
rect 265754 12518 265806 12570
rect 265858 12518 296318 12570
rect 296370 12518 296422 12570
rect 296474 12518 296526 12570
rect 296578 12518 298592 12570
rect 1344 12484 298592 12518
rect 1344 11786 298592 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 96638 11786
rect 96690 11734 96742 11786
rect 96794 11734 96846 11786
rect 96898 11734 127358 11786
rect 127410 11734 127462 11786
rect 127514 11734 127566 11786
rect 127618 11734 158078 11786
rect 158130 11734 158182 11786
rect 158234 11734 158286 11786
rect 158338 11734 188798 11786
rect 188850 11734 188902 11786
rect 188954 11734 189006 11786
rect 189058 11734 219518 11786
rect 219570 11734 219622 11786
rect 219674 11734 219726 11786
rect 219778 11734 250238 11786
rect 250290 11734 250342 11786
rect 250394 11734 250446 11786
rect 250498 11734 280958 11786
rect 281010 11734 281062 11786
rect 281114 11734 281166 11786
rect 281218 11734 298592 11786
rect 1344 11700 298592 11734
rect 1344 11002 298592 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 81278 11002
rect 81330 10950 81382 11002
rect 81434 10950 81486 11002
rect 81538 10950 111998 11002
rect 112050 10950 112102 11002
rect 112154 10950 112206 11002
rect 112258 10950 142718 11002
rect 142770 10950 142822 11002
rect 142874 10950 142926 11002
rect 142978 10950 173438 11002
rect 173490 10950 173542 11002
rect 173594 10950 173646 11002
rect 173698 10950 204158 11002
rect 204210 10950 204262 11002
rect 204314 10950 204366 11002
rect 204418 10950 234878 11002
rect 234930 10950 234982 11002
rect 235034 10950 235086 11002
rect 235138 10950 265598 11002
rect 265650 10950 265702 11002
rect 265754 10950 265806 11002
rect 265858 10950 296318 11002
rect 296370 10950 296422 11002
rect 296474 10950 296526 11002
rect 296578 10950 298592 11002
rect 1344 10916 298592 10950
rect 211934 10834 211986 10846
rect 211934 10770 211986 10782
rect 1344 10218 298592 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 96638 10218
rect 96690 10166 96742 10218
rect 96794 10166 96846 10218
rect 96898 10166 127358 10218
rect 127410 10166 127462 10218
rect 127514 10166 127566 10218
rect 127618 10166 158078 10218
rect 158130 10166 158182 10218
rect 158234 10166 158286 10218
rect 158338 10166 188798 10218
rect 188850 10166 188902 10218
rect 188954 10166 189006 10218
rect 189058 10166 219518 10218
rect 219570 10166 219622 10218
rect 219674 10166 219726 10218
rect 219778 10166 250238 10218
rect 250290 10166 250342 10218
rect 250394 10166 250446 10218
rect 250498 10166 280958 10218
rect 281010 10166 281062 10218
rect 281114 10166 281166 10218
rect 281218 10166 298592 10218
rect 1344 10132 298592 10166
rect 199166 9938 199218 9950
rect 199166 9874 199218 9886
rect 200062 9938 200114 9950
rect 200062 9874 200114 9886
rect 217422 9938 217474 9950
rect 217422 9874 217474 9886
rect 220894 9938 220946 9950
rect 220894 9874 220946 9886
rect 211486 9826 211538 9838
rect 211486 9762 211538 9774
rect 211710 9826 211762 9838
rect 211710 9762 211762 9774
rect 212046 9826 212098 9838
rect 212482 9774 212494 9826
rect 212546 9774 212558 9826
rect 212046 9762 212098 9774
rect 211038 9714 211090 9726
rect 211038 9650 211090 9662
rect 200958 9602 201010 9614
rect 200958 9538 201010 9550
rect 210926 9602 210978 9614
rect 210926 9538 210978 9550
rect 211262 9602 211314 9614
rect 211262 9538 211314 9550
rect 1344 9434 298592 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 81278 9434
rect 81330 9382 81382 9434
rect 81434 9382 81486 9434
rect 81538 9382 111998 9434
rect 112050 9382 112102 9434
rect 112154 9382 112206 9434
rect 112258 9382 142718 9434
rect 142770 9382 142822 9434
rect 142874 9382 142926 9434
rect 142978 9382 173438 9434
rect 173490 9382 173542 9434
rect 173594 9382 173646 9434
rect 173698 9382 204158 9434
rect 204210 9382 204262 9434
rect 204314 9382 204366 9434
rect 204418 9382 234878 9434
rect 234930 9382 234982 9434
rect 235034 9382 235086 9434
rect 235138 9382 265598 9434
rect 265650 9382 265702 9434
rect 265754 9382 265806 9434
rect 265858 9382 296318 9434
rect 296370 9382 296422 9434
rect 296474 9382 296526 9434
rect 296578 9382 298592 9434
rect 1344 9348 298592 9382
rect 188862 9266 188914 9278
rect 188862 9202 188914 9214
rect 196030 9266 196082 9278
rect 196030 9202 196082 9214
rect 198494 9266 198546 9278
rect 198494 9202 198546 9214
rect 198830 9266 198882 9278
rect 198830 9202 198882 9214
rect 201294 9266 201346 9278
rect 201294 9202 201346 9214
rect 202302 9266 202354 9278
rect 202302 9202 202354 9214
rect 203086 9266 203138 9278
rect 203086 9202 203138 9214
rect 203646 9266 203698 9278
rect 203646 9202 203698 9214
rect 216750 9266 216802 9278
rect 216750 9202 216802 9214
rect 219102 9266 219154 9278
rect 219102 9202 219154 9214
rect 219550 9266 219602 9278
rect 219550 9202 219602 9214
rect 220446 9266 220498 9278
rect 220446 9202 220498 9214
rect 222350 9266 222402 9278
rect 222350 9202 222402 9214
rect 200398 9154 200450 9166
rect 217198 9154 217250 9166
rect 195570 9102 195582 9154
rect 195634 9102 195646 9154
rect 199154 9102 199166 9154
rect 199218 9102 199230 9154
rect 208114 9102 208126 9154
rect 208178 9102 208190 9154
rect 210130 9102 210142 9154
rect 210194 9102 210206 9154
rect 211250 9102 211262 9154
rect 211314 9102 211326 9154
rect 200398 9090 200450 9102
rect 217198 9090 217250 9102
rect 217758 9154 217810 9166
rect 217758 9090 217810 9102
rect 218430 9154 218482 9166
rect 218430 9090 218482 9102
rect 219998 9154 220050 9166
rect 219998 9090 220050 9102
rect 220670 9154 220722 9166
rect 220670 9090 220722 9102
rect 221230 9154 221282 9166
rect 221230 9090 221282 9102
rect 221902 9154 221954 9166
rect 221902 9090 221954 9102
rect 192670 9042 192722 9054
rect 193678 9042 193730 9054
rect 199726 9042 199778 9054
rect 192994 8990 193006 9042
rect 193058 8990 193070 9042
rect 195346 8990 195358 9042
rect 195410 8990 195422 9042
rect 192670 8978 192722 8990
rect 193678 8978 193730 8990
rect 199726 8978 199778 8990
rect 205774 9042 205826 9054
rect 205774 8978 205826 8990
rect 207790 9042 207842 9054
rect 212718 9042 212770 9054
rect 210802 8990 210814 9042
rect 210866 8990 210878 9042
rect 207790 8978 207842 8990
rect 212718 8978 212770 8990
rect 213390 9042 213442 9054
rect 216526 9042 216578 9054
rect 213826 8990 213838 9042
rect 213890 8990 213902 9042
rect 213390 8978 213442 8990
rect 216526 8978 216578 8990
rect 216974 9042 217026 9054
rect 216974 8978 217026 8990
rect 217982 9042 218034 9054
rect 217982 8978 218034 8990
rect 218206 9042 218258 9054
rect 218206 8978 218258 8990
rect 218766 9042 218818 9054
rect 218766 8978 218818 8990
rect 220222 9042 220274 9054
rect 220222 8978 220274 8990
rect 221454 9042 221506 9054
rect 221454 8978 221506 8990
rect 221678 9042 221730 9054
rect 221678 8978 221730 8990
rect 189422 8930 189474 8942
rect 189422 8866 189474 8878
rect 199502 8930 199554 8942
rect 199502 8866 199554 8878
rect 200958 8930 201010 8942
rect 200958 8866 201010 8878
rect 201854 8930 201906 8942
rect 201854 8866 201906 8878
rect 203198 8930 203250 8942
rect 203198 8866 203250 8878
rect 206334 8930 206386 8942
rect 206334 8866 206386 8878
rect 209246 8930 209298 8942
rect 216414 8930 216466 8942
rect 210018 8878 210030 8930
rect 210082 8878 210094 8930
rect 209246 8866 209298 8878
rect 216414 8866 216466 8878
rect 217870 8818 217922 8830
rect 200050 8766 200062 8818
rect 200114 8766 200126 8818
rect 217870 8754 217922 8766
rect 220558 8818 220610 8830
rect 220558 8754 220610 8766
rect 221790 8818 221842 8830
rect 221790 8754 221842 8766
rect 1344 8650 298592 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 96638 8650
rect 96690 8598 96742 8650
rect 96794 8598 96846 8650
rect 96898 8598 127358 8650
rect 127410 8598 127462 8650
rect 127514 8598 127566 8650
rect 127618 8598 158078 8650
rect 158130 8598 158182 8650
rect 158234 8598 158286 8650
rect 158338 8598 188798 8650
rect 188850 8598 188902 8650
rect 188954 8598 189006 8650
rect 189058 8598 219518 8650
rect 219570 8598 219622 8650
rect 219674 8598 219726 8650
rect 219778 8598 250238 8650
rect 250290 8598 250342 8650
rect 250394 8598 250446 8650
rect 250498 8598 280958 8650
rect 281010 8598 281062 8650
rect 281114 8598 281166 8650
rect 281218 8598 298592 8650
rect 1344 8564 298592 8598
rect 212270 8482 212322 8494
rect 212270 8418 212322 8430
rect 221342 8482 221394 8494
rect 221342 8418 221394 8430
rect 199054 8370 199106 8382
rect 187618 8318 187630 8370
rect 187682 8318 187694 8370
rect 189746 8318 189758 8370
rect 189810 8318 189822 8370
rect 199054 8306 199106 8318
rect 199614 8370 199666 8382
rect 199614 8306 199666 8318
rect 207678 8370 207730 8382
rect 207678 8306 207730 8318
rect 222014 8370 222066 8382
rect 222014 8306 222066 8318
rect 189086 8258 189138 8270
rect 188626 8206 188638 8258
rect 188690 8206 188702 8258
rect 189086 8194 189138 8206
rect 190766 8258 190818 8270
rect 190766 8194 190818 8206
rect 199950 8258 200002 8270
rect 203422 8258 203474 8270
rect 205102 8258 205154 8270
rect 210702 8258 210754 8270
rect 200834 8206 200846 8258
rect 200898 8206 200910 8258
rect 203186 8206 203198 8258
rect 203250 8206 203262 8258
rect 204642 8206 204654 8258
rect 204706 8206 204718 8258
rect 205874 8206 205886 8258
rect 205938 8206 205950 8258
rect 199950 8194 200002 8206
rect 203422 8194 203474 8206
rect 205102 8194 205154 8206
rect 210702 8194 210754 8206
rect 211150 8258 211202 8270
rect 211150 8194 211202 8206
rect 211710 8258 211762 8270
rect 211710 8194 211762 8206
rect 212382 8258 212434 8270
rect 212382 8194 212434 8206
rect 213390 8258 213442 8270
rect 220782 8258 220834 8270
rect 217522 8206 217534 8258
rect 217586 8206 217598 8258
rect 213390 8194 213442 8206
rect 220782 8194 220834 8206
rect 221454 8258 221506 8270
rect 221454 8194 221506 8206
rect 200062 8146 200114 8158
rect 200062 8082 200114 8094
rect 202190 8146 202242 8158
rect 202190 8082 202242 8094
rect 206894 8146 206946 8158
rect 206894 8082 206946 8094
rect 210366 8146 210418 8158
rect 210366 8082 210418 8094
rect 211374 8146 211426 8158
rect 211374 8082 211426 8094
rect 212830 8146 212882 8158
rect 212830 8082 212882 8094
rect 217758 8146 217810 8158
rect 217758 8082 217810 8094
rect 221006 8146 221058 8158
rect 221006 8082 221058 8094
rect 190430 8034 190482 8046
rect 190430 7970 190482 7982
rect 201070 8034 201122 8046
rect 201070 7970 201122 7982
rect 203086 8034 203138 8046
rect 203086 7970 203138 7982
rect 205662 8034 205714 8046
rect 205662 7970 205714 7982
rect 205998 8034 206050 8046
rect 205998 7970 206050 7982
rect 209806 8034 209858 8046
rect 209806 7970 209858 7982
rect 210590 8034 210642 8046
rect 210590 7970 210642 7982
rect 210926 8034 210978 8046
rect 210926 7970 210978 7982
rect 211934 8034 211986 8046
rect 211934 7970 211986 7982
rect 212158 8034 212210 8046
rect 212158 7970 212210 7982
rect 221230 8034 221282 8046
rect 221230 7970 221282 7982
rect 1344 7866 298592 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 81278 7866
rect 81330 7814 81382 7866
rect 81434 7814 81486 7866
rect 81538 7814 111998 7866
rect 112050 7814 112102 7866
rect 112154 7814 112206 7866
rect 112258 7814 142718 7866
rect 142770 7814 142822 7866
rect 142874 7814 142926 7866
rect 142978 7814 173438 7866
rect 173490 7814 173542 7866
rect 173594 7814 173646 7866
rect 173698 7814 204158 7866
rect 204210 7814 204262 7866
rect 204314 7814 204366 7866
rect 204418 7814 234878 7866
rect 234930 7814 234982 7866
rect 235034 7814 235086 7866
rect 235138 7814 265598 7866
rect 265650 7814 265702 7866
rect 265754 7814 265806 7866
rect 265858 7814 296318 7866
rect 296370 7814 296422 7866
rect 296474 7814 296526 7866
rect 296578 7814 298592 7866
rect 1344 7780 298592 7814
rect 196030 7698 196082 7710
rect 196030 7634 196082 7646
rect 202862 7698 202914 7710
rect 202862 7634 202914 7646
rect 204878 7698 204930 7710
rect 204878 7634 204930 7646
rect 207342 7698 207394 7710
rect 207342 7634 207394 7646
rect 215742 7698 215794 7710
rect 215742 7634 215794 7646
rect 185390 7586 185442 7598
rect 191102 7586 191154 7598
rect 186274 7534 186286 7586
rect 186338 7534 186350 7586
rect 188066 7534 188078 7586
rect 188130 7534 188142 7586
rect 188738 7534 188750 7586
rect 188802 7534 188814 7586
rect 189298 7534 189310 7586
rect 189362 7534 189374 7586
rect 185390 7522 185442 7534
rect 191102 7522 191154 7534
rect 192670 7586 192722 7598
rect 202414 7586 202466 7598
rect 195570 7534 195582 7586
rect 195634 7534 195646 7586
rect 201058 7534 201070 7586
rect 201122 7534 201134 7586
rect 192670 7522 192722 7534
rect 202414 7522 202466 7534
rect 204654 7586 204706 7598
rect 209906 7534 209918 7586
rect 209970 7534 209982 7586
rect 211586 7534 211598 7586
rect 211650 7534 211662 7586
rect 204654 7522 204706 7534
rect 190654 7474 190706 7486
rect 198494 7474 198546 7486
rect 185602 7422 185614 7474
rect 185666 7422 185678 7474
rect 187842 7422 187854 7474
rect 187906 7422 187918 7474
rect 189186 7422 189198 7474
rect 189250 7422 189262 7474
rect 192882 7422 192894 7474
rect 192946 7422 192958 7474
rect 193778 7422 193790 7474
rect 193842 7422 193854 7474
rect 195122 7422 195134 7474
rect 195186 7422 195198 7474
rect 190654 7410 190706 7422
rect 198494 7410 198546 7422
rect 200398 7474 200450 7486
rect 214062 7474 214114 7486
rect 216414 7474 216466 7486
rect 200834 7422 200846 7474
rect 200898 7422 200910 7474
rect 202962 7422 202974 7474
rect 203026 7422 203038 7474
rect 205762 7422 205774 7474
rect 205826 7422 205838 7474
rect 210354 7422 210366 7474
rect 210418 7422 210430 7474
rect 210914 7422 210926 7474
rect 210978 7422 210990 7474
rect 214498 7422 214510 7474
rect 214562 7422 214574 7474
rect 216178 7422 216190 7474
rect 216242 7422 216254 7474
rect 200398 7410 200450 7422
rect 214062 7410 214114 7422
rect 216414 7410 216466 7422
rect 216526 7474 216578 7486
rect 216526 7410 216578 7422
rect 191662 7362 191714 7374
rect 191662 7298 191714 7310
rect 199166 7362 199218 7374
rect 199166 7298 199218 7310
rect 199614 7362 199666 7374
rect 199614 7298 199666 7310
rect 203198 7362 203250 7374
rect 206334 7362 206386 7374
rect 209470 7362 209522 7374
rect 204866 7310 204878 7362
rect 204930 7310 204942 7362
rect 205538 7310 205550 7362
rect 205602 7310 205614 7362
rect 206882 7310 206894 7362
rect 206946 7310 206958 7362
rect 203198 7298 203250 7310
rect 206334 7298 206386 7310
rect 209470 7298 209522 7310
rect 216750 7362 216802 7374
rect 216750 7298 216802 7310
rect 189870 7250 189922 7262
rect 189870 7186 189922 7198
rect 197710 7250 197762 7262
rect 200174 7250 200226 7262
rect 199826 7198 199838 7250
rect 199890 7198 199902 7250
rect 197710 7186 197762 7198
rect 200174 7186 200226 7198
rect 1344 7082 298592 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 96638 7082
rect 96690 7030 96742 7082
rect 96794 7030 96846 7082
rect 96898 7030 127358 7082
rect 127410 7030 127462 7082
rect 127514 7030 127566 7082
rect 127618 7030 158078 7082
rect 158130 7030 158182 7082
rect 158234 7030 158286 7082
rect 158338 7030 188798 7082
rect 188850 7030 188902 7082
rect 188954 7030 189006 7082
rect 189058 7030 219518 7082
rect 219570 7030 219622 7082
rect 219674 7030 219726 7082
rect 219778 7030 250238 7082
rect 250290 7030 250342 7082
rect 250394 7030 250446 7082
rect 250498 7030 280958 7082
rect 281010 7030 281062 7082
rect 281114 7030 281166 7082
rect 281218 7030 298592 7082
rect 1344 6996 298592 7030
rect 199390 6802 199442 6814
rect 199390 6738 199442 6750
rect 217758 6802 217810 6814
rect 217758 6738 217810 6750
rect 184494 6690 184546 6702
rect 184494 6626 184546 6638
rect 186734 6690 186786 6702
rect 193230 6690 193282 6702
rect 187730 6638 187742 6690
rect 187794 6638 187806 6690
rect 190306 6638 190318 6690
rect 190370 6638 190382 6690
rect 190642 6638 190654 6690
rect 190706 6638 190718 6690
rect 190978 6638 190990 6690
rect 191042 6638 191054 6690
rect 192322 6638 192334 6690
rect 192386 6638 192398 6690
rect 186734 6626 186786 6638
rect 193230 6626 193282 6638
rect 193902 6690 193954 6702
rect 193902 6626 193954 6638
rect 195918 6690 195970 6702
rect 207454 6690 207506 6702
rect 217198 6690 217250 6702
rect 196802 6638 196814 6690
rect 196866 6638 196878 6690
rect 197586 6638 197598 6690
rect 197650 6638 197662 6690
rect 197922 6638 197934 6690
rect 197986 6638 197998 6690
rect 198594 6638 198606 6690
rect 198658 6638 198670 6690
rect 201058 6638 201070 6690
rect 201122 6638 201134 6690
rect 201618 6638 201630 6690
rect 201682 6638 201694 6690
rect 203074 6638 203086 6690
rect 203138 6638 203150 6690
rect 204642 6638 204654 6690
rect 204706 6638 204718 6690
rect 206322 6638 206334 6690
rect 206386 6638 206398 6690
rect 213826 6638 213838 6690
rect 213890 6638 213902 6690
rect 195918 6626 195970 6638
rect 207454 6626 207506 6638
rect 217198 6626 217250 6638
rect 218206 6690 218258 6702
rect 218206 6626 218258 6638
rect 184382 6578 184434 6590
rect 188290 6526 188302 6578
rect 188354 6526 188366 6578
rect 199602 6526 199614 6578
rect 199666 6526 199678 6578
rect 204754 6526 204766 6578
rect 204818 6526 204830 6578
rect 205090 6526 205102 6578
rect 205154 6526 205166 6578
rect 184382 6514 184434 6526
rect 184046 6466 184098 6478
rect 192782 6466 192834 6478
rect 187394 6414 187406 6466
rect 187458 6414 187470 6466
rect 184046 6402 184098 6414
rect 192782 6402 192834 6414
rect 194350 6466 194402 6478
rect 207006 6466 207058 6478
rect 204642 6414 204654 6466
rect 204706 6414 204718 6466
rect 194350 6402 194402 6414
rect 207006 6402 207058 6414
rect 207902 6466 207954 6478
rect 217646 6466 217698 6478
rect 213602 6414 213614 6466
rect 213666 6414 213678 6466
rect 207902 6402 207954 6414
rect 217646 6402 217698 6414
rect 217870 6466 217922 6478
rect 219102 6466 219154 6478
rect 218530 6414 218542 6466
rect 218594 6414 218606 6466
rect 217870 6402 217922 6414
rect 219102 6402 219154 6414
rect 1344 6298 298592 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 81278 6298
rect 81330 6246 81382 6298
rect 81434 6246 81486 6298
rect 81538 6246 111998 6298
rect 112050 6246 112102 6298
rect 112154 6246 112206 6298
rect 112258 6246 142718 6298
rect 142770 6246 142822 6298
rect 142874 6246 142926 6298
rect 142978 6246 173438 6298
rect 173490 6246 173542 6298
rect 173594 6246 173646 6298
rect 173698 6246 204158 6298
rect 204210 6246 204262 6298
rect 204314 6246 204366 6298
rect 204418 6246 234878 6298
rect 234930 6246 234982 6298
rect 235034 6246 235086 6298
rect 235138 6246 265598 6298
rect 265650 6246 265702 6298
rect 265754 6246 265806 6298
rect 265858 6246 296318 6298
rect 296370 6246 296422 6298
rect 296474 6246 296526 6298
rect 296578 6246 298592 6298
rect 1344 6212 298592 6246
rect 187518 6130 187570 6142
rect 203534 6130 203586 6142
rect 185266 6078 185278 6130
rect 185330 6078 185342 6130
rect 193554 6078 193566 6130
rect 193618 6078 193630 6130
rect 197698 6078 197710 6130
rect 197762 6078 197774 6130
rect 187518 6066 187570 6078
rect 203534 6066 203586 6078
rect 209470 6130 209522 6142
rect 209470 6066 209522 6078
rect 214622 6130 214674 6142
rect 214622 6066 214674 6078
rect 187966 6018 188018 6030
rect 186386 5966 186398 6018
rect 186450 5966 186462 6018
rect 187966 5954 188018 5966
rect 191662 6018 191714 6030
rect 191662 5954 191714 5966
rect 191774 6018 191826 6030
rect 205550 6018 205602 6030
rect 216638 6018 216690 6030
rect 195570 5966 195582 6018
rect 195634 5966 195646 6018
rect 199154 5966 199166 6018
rect 199218 5966 199230 6018
rect 199490 5966 199502 6018
rect 199554 5966 199566 6018
rect 214946 5966 214958 6018
rect 215010 5966 215022 6018
rect 191774 5954 191826 5966
rect 205550 5954 205602 5966
rect 216638 5954 216690 5966
rect 186734 5906 186786 5918
rect 183698 5854 183710 5906
rect 183762 5854 183774 5906
rect 184594 5854 184606 5906
rect 184658 5854 184670 5906
rect 186162 5854 186174 5906
rect 186226 5854 186238 5906
rect 186734 5842 186786 5854
rect 189310 5906 189362 5918
rect 196030 5906 196082 5918
rect 205774 5906 205826 5918
rect 191090 5854 191102 5906
rect 191154 5854 191166 5906
rect 192882 5854 192894 5906
rect 192946 5854 192958 5906
rect 193778 5854 193790 5906
rect 193842 5854 193854 5906
rect 195346 5854 195358 5906
rect 195410 5854 195422 5906
rect 198034 5854 198046 5906
rect 198098 5854 198110 5906
rect 200610 5854 200622 5906
rect 200674 5854 200686 5906
rect 201282 5854 201294 5906
rect 201346 5854 201358 5906
rect 201842 5854 201854 5906
rect 201906 5854 201918 5906
rect 204530 5854 204542 5906
rect 204594 5854 204606 5906
rect 189310 5842 189362 5854
rect 196030 5842 196082 5854
rect 205774 5842 205826 5854
rect 205998 5906 206050 5918
rect 205998 5842 206050 5854
rect 206222 5906 206274 5918
rect 206222 5842 206274 5854
rect 206558 5906 206610 5918
rect 206558 5842 206610 5854
rect 210366 5906 210418 5918
rect 210366 5842 210418 5854
rect 210814 5906 210866 5918
rect 210814 5842 210866 5854
rect 211262 5906 211314 5918
rect 211262 5842 211314 5854
rect 211374 5906 211426 5918
rect 216178 5854 216190 5906
rect 216242 5854 216254 5906
rect 216402 5854 216414 5906
rect 216466 5854 216478 5906
rect 211374 5842 211426 5854
rect 203982 5794 204034 5806
rect 188850 5742 188862 5794
rect 188914 5742 188926 5794
rect 190418 5742 190430 5794
rect 190482 5742 190494 5794
rect 203074 5742 203086 5794
rect 203138 5742 203150 5794
rect 203982 5730 204034 5742
rect 204990 5794 205042 5806
rect 207566 5794 207618 5806
rect 206994 5742 207006 5794
rect 207058 5742 207070 5794
rect 204990 5730 205042 5742
rect 207566 5730 207618 5742
rect 208014 5794 208066 5806
rect 208014 5730 208066 5742
rect 208462 5794 208514 5806
rect 208462 5730 208514 5742
rect 208910 5794 208962 5806
rect 208910 5730 208962 5742
rect 209806 5794 209858 5806
rect 209806 5730 209858 5742
rect 211598 5794 211650 5806
rect 211598 5730 211650 5742
rect 215854 5794 215906 5806
rect 217086 5794 217138 5806
rect 216514 5742 216526 5794
rect 216578 5742 216590 5794
rect 215854 5730 215906 5742
rect 217086 5730 217138 5742
rect 219550 5794 219602 5806
rect 219550 5730 219602 5742
rect 223582 5794 223634 5806
rect 223582 5730 223634 5742
rect 196814 5682 196866 5694
rect 196814 5618 196866 5630
rect 206110 5682 206162 5694
rect 210590 5682 210642 5694
rect 207442 5630 207454 5682
rect 207506 5679 207518 5682
rect 208002 5679 208014 5682
rect 207506 5633 208014 5679
rect 207506 5630 207518 5633
rect 208002 5630 208014 5633
rect 208066 5630 208078 5682
rect 206110 5618 206162 5630
rect 210590 5618 210642 5630
rect 1344 5514 298592 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 96638 5514
rect 96690 5462 96742 5514
rect 96794 5462 96846 5514
rect 96898 5462 127358 5514
rect 127410 5462 127462 5514
rect 127514 5462 127566 5514
rect 127618 5462 158078 5514
rect 158130 5462 158182 5514
rect 158234 5462 158286 5514
rect 158338 5462 188798 5514
rect 188850 5462 188902 5514
rect 188954 5462 189006 5514
rect 189058 5462 219518 5514
rect 219570 5462 219622 5514
rect 219674 5462 219726 5514
rect 219778 5462 250238 5514
rect 250290 5462 250342 5514
rect 250394 5462 250446 5514
rect 250498 5462 280958 5514
rect 281010 5462 281062 5514
rect 281114 5462 281166 5514
rect 281218 5462 298592 5514
rect 1344 5428 298592 5462
rect 192782 5346 192834 5358
rect 192782 5282 192834 5294
rect 204094 5346 204146 5358
rect 204094 5282 204146 5294
rect 207342 5346 207394 5358
rect 207342 5282 207394 5294
rect 210478 5346 210530 5358
rect 210478 5282 210530 5294
rect 218318 5346 218370 5358
rect 218318 5282 218370 5294
rect 220782 5346 220834 5358
rect 220782 5282 220834 5294
rect 220894 5346 220946 5358
rect 220894 5282 220946 5294
rect 93550 5234 93602 5246
rect 192670 5234 192722 5246
rect 185938 5182 185950 5234
rect 186002 5182 186014 5234
rect 93550 5170 93602 5182
rect 192670 5170 192722 5182
rect 193230 5234 193282 5246
rect 193230 5170 193282 5182
rect 195022 5234 195074 5246
rect 195022 5170 195074 5182
rect 195470 5234 195522 5246
rect 195470 5170 195522 5182
rect 206558 5234 206610 5246
rect 206558 5170 206610 5182
rect 215294 5234 215346 5246
rect 215294 5170 215346 5182
rect 217310 5234 217362 5246
rect 217310 5170 217362 5182
rect 185390 5122 185442 5134
rect 187070 5122 187122 5134
rect 194574 5122 194626 5134
rect 204094 5122 204146 5134
rect 182690 5070 182702 5122
rect 182754 5070 182766 5122
rect 183586 5070 183598 5122
rect 183650 5070 183662 5122
rect 184706 5070 184718 5122
rect 184770 5070 184782 5122
rect 186386 5070 186398 5122
rect 186450 5070 186462 5122
rect 187506 5070 187518 5122
rect 187570 5070 187582 5122
rect 190306 5070 190318 5122
rect 190370 5070 190382 5122
rect 190642 5070 190654 5122
rect 190706 5070 190718 5122
rect 190978 5070 190990 5122
rect 191042 5070 191054 5122
rect 192322 5070 192334 5122
rect 192386 5070 192398 5122
rect 196242 5070 196254 5122
rect 196306 5070 196318 5122
rect 199042 5070 199054 5122
rect 199106 5070 199118 5122
rect 199714 5070 199726 5122
rect 199778 5070 199790 5122
rect 201058 5070 201070 5122
rect 201122 5070 201134 5122
rect 201730 5070 201742 5122
rect 201794 5070 201806 5122
rect 202514 5070 202526 5122
rect 202578 5070 202590 5122
rect 202962 5070 202974 5122
rect 203026 5070 203038 5122
rect 185390 5058 185442 5070
rect 187070 5058 187122 5070
rect 194574 5058 194626 5070
rect 204094 5058 204146 5070
rect 204542 5122 204594 5134
rect 204542 5058 204594 5070
rect 205102 5122 205154 5134
rect 205102 5058 205154 5070
rect 205774 5122 205826 5134
rect 205774 5058 205826 5070
rect 206446 5122 206498 5134
rect 206446 5058 206498 5070
rect 206782 5122 206834 5134
rect 206782 5058 206834 5070
rect 207454 5122 207506 5134
rect 207454 5058 207506 5070
rect 208014 5122 208066 5134
rect 209470 5122 209522 5134
rect 208786 5070 208798 5122
rect 208850 5070 208862 5122
rect 208014 5058 208066 5070
rect 209470 5058 209522 5070
rect 210254 5122 210306 5134
rect 210254 5058 210306 5070
rect 210702 5122 210754 5134
rect 210702 5058 210754 5070
rect 212270 5122 212322 5134
rect 214734 5122 214786 5134
rect 214274 5070 214286 5122
rect 214338 5070 214350 5122
rect 212270 5058 212322 5070
rect 214734 5058 214786 5070
rect 215182 5122 215234 5134
rect 215182 5058 215234 5070
rect 215630 5122 215682 5134
rect 215630 5058 215682 5070
rect 216190 5122 216242 5134
rect 216190 5058 216242 5070
rect 216862 5122 216914 5134
rect 218990 5122 219042 5134
rect 217970 5070 217982 5122
rect 218034 5070 218046 5122
rect 218530 5070 218542 5122
rect 218594 5070 218606 5122
rect 216862 5058 216914 5070
rect 218990 5058 219042 5070
rect 219774 5122 219826 5134
rect 219774 5058 219826 5070
rect 220558 5122 220610 5134
rect 220558 5058 220610 5070
rect 221118 5122 221170 5134
rect 221118 5058 221170 5070
rect 221566 5122 221618 5134
rect 221566 5058 221618 5070
rect 221790 5122 221842 5134
rect 221790 5058 221842 5070
rect 222574 5122 222626 5134
rect 222574 5058 222626 5070
rect 223470 5122 223522 5134
rect 223470 5058 223522 5070
rect 224030 5122 224082 5134
rect 224030 5058 224082 5070
rect 201966 5010 202018 5022
rect 186610 4958 186622 5010
rect 186674 4958 186686 5010
rect 188850 4958 188862 5010
rect 188914 4958 188926 5010
rect 197586 4958 197598 5010
rect 197650 4958 197662 5010
rect 197922 4958 197934 5010
rect 197986 4958 197998 5010
rect 201966 4946 202018 4958
rect 203534 5010 203586 5022
rect 203534 4946 203586 4958
rect 203982 5010 204034 5022
rect 203982 4946 204034 4958
rect 205998 5010 206050 5022
rect 205998 4946 206050 4958
rect 207230 5010 207282 5022
rect 207230 4946 207282 4958
rect 208350 5010 208402 5022
rect 212382 5010 212434 5022
rect 209570 4958 209582 5010
rect 209634 4958 209646 5010
rect 209906 4958 209918 5010
rect 209970 4958 209982 5010
rect 208350 4946 208402 4958
rect 212382 4946 212434 4958
rect 212606 5010 212658 5022
rect 212606 4946 212658 4958
rect 212830 5010 212882 5022
rect 212830 4946 212882 4958
rect 216078 5010 216130 5022
rect 218878 5010 218930 5022
rect 217410 4958 217422 5010
rect 217474 4958 217486 5010
rect 217746 4958 217758 5010
rect 217810 4958 217822 5010
rect 216078 4946 216130 4958
rect 218878 4946 218930 4958
rect 219998 5010 220050 5022
rect 221678 5010 221730 5022
rect 220210 4958 220222 5010
rect 220274 4958 220286 5010
rect 219998 4946 220050 4958
rect 221678 4946 221730 4958
rect 193118 4898 193170 4910
rect 183362 4846 183374 4898
rect 183426 4846 183438 4898
rect 187394 4846 187406 4898
rect 187458 4846 187470 4898
rect 193118 4834 193170 4846
rect 193790 4898 193842 4910
rect 203086 4898 203138 4910
rect 196130 4846 196142 4898
rect 196194 4846 196206 4898
rect 193790 4834 193842 4846
rect 203086 4834 203138 4846
rect 203758 4898 203810 4910
rect 203758 4834 203810 4846
rect 206222 4898 206274 4910
rect 206222 4834 206274 4846
rect 207006 4898 207058 4910
rect 215406 4898 215458 4910
rect 211026 4846 211038 4898
rect 211090 4846 211102 4898
rect 211810 4846 211822 4898
rect 211874 4846 211886 4898
rect 214498 4846 214510 4898
rect 214562 4846 214574 4898
rect 207006 4834 207058 4846
rect 215406 4834 215458 4846
rect 216302 4898 216354 4910
rect 216302 4834 216354 4846
rect 219102 4898 219154 4910
rect 219102 4834 219154 4846
rect 223022 4898 223074 4910
rect 223022 4834 223074 4846
rect 223134 4898 223186 4910
rect 223134 4834 223186 4846
rect 223246 4898 223298 4910
rect 223246 4834 223298 4846
rect 223918 4898 223970 4910
rect 223918 4834 223970 4846
rect 224142 4898 224194 4910
rect 224142 4834 224194 4846
rect 224702 4898 224754 4910
rect 224702 4834 224754 4846
rect 1344 4730 298592 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 81278 4730
rect 81330 4678 81382 4730
rect 81434 4678 81486 4730
rect 81538 4678 111998 4730
rect 112050 4678 112102 4730
rect 112154 4678 112206 4730
rect 112258 4678 142718 4730
rect 142770 4678 142822 4730
rect 142874 4678 142926 4730
rect 142978 4678 173438 4730
rect 173490 4678 173542 4730
rect 173594 4678 173646 4730
rect 173698 4678 204158 4730
rect 204210 4678 204262 4730
rect 204314 4678 204366 4730
rect 204418 4678 234878 4730
rect 234930 4678 234982 4730
rect 235034 4678 235086 4730
rect 235138 4678 265598 4730
rect 265650 4678 265702 4730
rect 265754 4678 265806 4730
rect 265858 4678 296318 4730
rect 296370 4678 296422 4730
rect 296474 4678 296526 4730
rect 296578 4678 298592 4730
rect 1344 4644 298592 4678
rect 12462 4562 12514 4574
rect 12462 4498 12514 4510
rect 54350 4562 54402 4574
rect 54350 4498 54402 4510
rect 71150 4562 71202 4574
rect 71150 4498 71202 4510
rect 74846 4562 74898 4574
rect 74846 4498 74898 4510
rect 96238 4562 96290 4574
rect 96238 4498 96290 4510
rect 122558 4562 122610 4574
rect 122558 4498 122610 4510
rect 182366 4562 182418 4574
rect 189310 4562 189362 4574
rect 195358 4562 195410 4574
rect 184706 4510 184718 4562
rect 184770 4510 184782 4562
rect 189858 4510 189870 4562
rect 189922 4510 189934 4562
rect 182366 4498 182418 4510
rect 189310 4498 189362 4510
rect 195358 4498 195410 4510
rect 196366 4562 196418 4574
rect 196366 4498 196418 4510
rect 197150 4562 197202 4574
rect 204878 4562 204930 4574
rect 197698 4510 197710 4562
rect 197762 4510 197774 4562
rect 197150 4498 197202 4510
rect 204878 4498 204930 4510
rect 212494 4562 212546 4574
rect 212494 4498 212546 4510
rect 212606 4562 212658 4574
rect 212606 4498 212658 4510
rect 215294 4562 215346 4574
rect 215294 4498 215346 4510
rect 215406 4562 215458 4574
rect 215406 4498 215458 4510
rect 215966 4562 216018 4574
rect 215966 4498 216018 4510
rect 217086 4562 217138 4574
rect 217086 4498 217138 4510
rect 217310 4562 217362 4574
rect 217310 4498 217362 4510
rect 220110 4562 220162 4574
rect 220110 4498 220162 4510
rect 11566 4450 11618 4462
rect 11566 4386 11618 4398
rect 11902 4450 11954 4462
rect 11902 4386 11954 4398
rect 71374 4450 71426 4462
rect 71374 4386 71426 4398
rect 71710 4450 71762 4462
rect 71710 4386 71762 4398
rect 75070 4450 75122 4462
rect 75070 4386 75122 4398
rect 75406 4450 75458 4462
rect 75406 4386 75458 4398
rect 83134 4450 83186 4462
rect 83134 4386 83186 4398
rect 83470 4450 83522 4462
rect 83470 4386 83522 4398
rect 86718 4450 86770 4462
rect 86718 4386 86770 4398
rect 87054 4450 87106 4462
rect 87054 4386 87106 4398
rect 93886 4450 93938 4462
rect 93886 4386 93938 4398
rect 94222 4450 94274 4462
rect 94222 4386 94274 4398
rect 96462 4450 96514 4462
rect 96462 4386 96514 4398
rect 96798 4450 96850 4462
rect 216750 4450 216802 4462
rect 187954 4398 187966 4450
rect 188018 4398 188030 4450
rect 190530 4398 190542 4450
rect 190594 4398 190606 4450
rect 191650 4398 191662 4450
rect 191714 4398 191726 4450
rect 199154 4398 199166 4450
rect 199218 4398 199230 4450
rect 199490 4398 199502 4450
rect 199554 4398 199566 4450
rect 202962 4398 202974 4450
rect 203026 4398 203038 4450
rect 206994 4398 207006 4450
rect 207058 4398 207070 4450
rect 208226 4398 208238 4450
rect 208290 4398 208302 4450
rect 210802 4398 210814 4450
rect 210866 4398 210878 4450
rect 96798 4386 96850 4398
rect 216750 4386 216802 4398
rect 217534 4450 217586 4462
rect 217534 4386 217586 4398
rect 220670 4450 220722 4462
rect 220670 4386 220722 4398
rect 221790 4450 221842 4462
rect 221790 4386 221842 4398
rect 182814 4338 182866 4350
rect 186398 4338 186450 4350
rect 211934 4338 211986 4350
rect 214846 4338 214898 4350
rect 76626 4286 76638 4338
rect 76690 4286 76702 4338
rect 80210 4286 80222 4338
rect 80274 4286 80286 4338
rect 83794 4286 83806 4338
rect 83858 4286 83870 4338
rect 87938 4286 87950 4338
rect 88002 4286 88014 4338
rect 90962 4286 90974 4338
rect 91026 4286 91038 4338
rect 183698 4286 183710 4338
rect 183762 4286 183774 4338
rect 184594 4286 184606 4338
rect 184658 4286 184670 4338
rect 186162 4286 186174 4338
rect 186226 4286 186238 4338
rect 186722 4286 186734 4338
rect 186786 4286 186798 4338
rect 189858 4286 189870 4338
rect 189922 4286 189934 4338
rect 192770 4286 192782 4338
rect 192834 4286 192846 4338
rect 193442 4286 193454 4338
rect 193506 4286 193518 4338
rect 193666 4286 193678 4338
rect 193730 4286 193742 4338
rect 197698 4286 197710 4338
rect 197762 4286 197774 4338
rect 200610 4286 200622 4338
rect 200674 4286 200686 4338
rect 201282 4286 201294 4338
rect 201346 4286 201358 4338
rect 201842 4286 201854 4338
rect 201906 4286 201918 4338
rect 203186 4286 203198 4338
rect 203250 4286 203262 4338
rect 203746 4286 203758 4338
rect 203810 4286 203822 4338
rect 204194 4286 204206 4338
rect 204258 4286 204270 4338
rect 205538 4286 205550 4338
rect 205602 4286 205614 4338
rect 208786 4286 208798 4338
rect 208850 4286 208862 4338
rect 210018 4286 210030 4338
rect 210082 4286 210094 4338
rect 210242 4286 210254 4338
rect 210306 4286 210318 4338
rect 212258 4286 212270 4338
rect 212322 4286 212334 4338
rect 182814 4274 182866 4286
rect 186398 4274 186450 4286
rect 211934 4274 211986 4286
rect 214846 4274 214898 4286
rect 215518 4338 215570 4350
rect 217982 4338 218034 4350
rect 216514 4286 216526 4338
rect 216578 4286 216590 4338
rect 215518 4274 215570 4286
rect 217982 4274 218034 4286
rect 219550 4338 219602 4350
rect 221342 4338 221394 4350
rect 219874 4286 219886 4338
rect 219938 4286 219950 4338
rect 219550 4274 219602 4286
rect 221342 4274 221394 4286
rect 221902 4338 221954 4350
rect 221902 4274 221954 4286
rect 222014 4338 222066 4350
rect 222014 4274 222066 4286
rect 222574 4338 222626 4350
rect 222574 4274 222626 4286
rect 223022 4338 223074 4350
rect 223022 4274 223074 4286
rect 223246 4338 223298 4350
rect 223246 4274 223298 4286
rect 223694 4338 223746 4350
rect 223694 4274 223746 4286
rect 50766 4226 50818 4238
rect 111806 4226 111858 4238
rect 89058 4174 89070 4226
rect 89122 4174 89134 4226
rect 50766 4162 50818 4174
rect 111806 4162 111858 4174
rect 115390 4226 115442 4238
rect 115390 4162 115442 4174
rect 181582 4226 181634 4238
rect 181582 4162 181634 4174
rect 182254 4226 182306 4238
rect 182254 4162 182306 4174
rect 182702 4226 182754 4238
rect 182702 4162 182754 4174
rect 195806 4226 195858 4238
rect 217422 4226 217474 4238
rect 206882 4174 206894 4226
rect 206946 4174 206958 4226
rect 210354 4174 210366 4226
rect 210418 4174 210430 4226
rect 195806 4162 195858 4174
rect 217422 4162 217474 4174
rect 219326 4226 219378 4238
rect 223134 4226 223186 4238
rect 219986 4174 219998 4226
rect 220050 4174 220062 4226
rect 219326 4162 219378 4174
rect 223134 4162 223186 4174
rect 77646 4114 77698 4126
rect 77646 4050 77698 4062
rect 81230 4114 81282 4126
rect 81230 4050 81282 4062
rect 84814 4114 84866 4126
rect 84814 4050 84866 4062
rect 91982 4114 92034 4126
rect 204542 4114 204594 4126
rect 186834 4062 186846 4114
rect 186898 4062 186910 4114
rect 91982 4050 92034 4062
rect 204542 4050 204594 4062
rect 221118 4114 221170 4126
rect 221118 4050 221170 4062
rect 1344 3946 298592 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 96638 3946
rect 96690 3894 96742 3946
rect 96794 3894 96846 3946
rect 96898 3894 127358 3946
rect 127410 3894 127462 3946
rect 127514 3894 127566 3946
rect 127618 3894 158078 3946
rect 158130 3894 158182 3946
rect 158234 3894 158286 3946
rect 158338 3894 188798 3946
rect 188850 3894 188902 3946
rect 188954 3894 189006 3946
rect 189058 3894 219518 3946
rect 219570 3894 219622 3946
rect 219674 3894 219726 3946
rect 219778 3894 250238 3946
rect 250290 3894 250342 3946
rect 250394 3894 250446 3946
rect 250498 3894 280958 3946
rect 281010 3894 281062 3946
rect 281114 3894 281166 3946
rect 281218 3894 298592 3946
rect 1344 3860 298592 3894
rect 182366 3778 182418 3790
rect 220782 3778 220834 3790
rect 208226 3726 208238 3778
rect 208290 3775 208302 3778
rect 208674 3775 208686 3778
rect 208290 3729 208686 3775
rect 208290 3726 208302 3729
rect 208674 3726 208686 3729
rect 208738 3726 208750 3778
rect 215394 3726 215406 3778
rect 215458 3775 215470 3778
rect 216178 3775 216190 3778
rect 215458 3729 216190 3775
rect 215458 3726 215470 3729
rect 216178 3726 216190 3729
rect 216242 3726 216254 3778
rect 182366 3714 182418 3726
rect 220782 3714 220834 3726
rect 221566 3778 221618 3790
rect 221566 3714 221618 3726
rect 40686 3666 40738 3678
rect 40686 3602 40738 3614
rect 43822 3666 43874 3678
rect 43822 3602 43874 3614
rect 44494 3666 44546 3678
rect 44494 3602 44546 3614
rect 47630 3666 47682 3678
rect 47630 3602 47682 3614
rect 48190 3666 48242 3678
rect 48190 3602 48242 3614
rect 51774 3666 51826 3678
rect 51774 3602 51826 3614
rect 55358 3666 55410 3678
rect 55358 3602 55410 3614
rect 58270 3666 58322 3678
rect 58270 3602 58322 3614
rect 59054 3666 59106 3678
rect 59054 3602 59106 3614
rect 61966 3666 62018 3678
rect 61966 3602 62018 3614
rect 62862 3666 62914 3678
rect 62862 3602 62914 3614
rect 65774 3666 65826 3678
rect 65774 3602 65826 3614
rect 66670 3666 66722 3678
rect 66670 3602 66722 3614
rect 69582 3666 69634 3678
rect 69582 3602 69634 3614
rect 70478 3666 70530 3678
rect 70478 3602 70530 3614
rect 73390 3666 73442 3678
rect 73390 3602 73442 3614
rect 78318 3666 78370 3678
rect 78318 3602 78370 3614
rect 82910 3666 82962 3678
rect 82910 3602 82962 3614
rect 86494 3666 86546 3678
rect 86494 3602 86546 3614
rect 88734 3666 88786 3678
rect 88734 3602 88786 3614
rect 101614 3666 101666 3678
rect 101614 3602 101666 3614
rect 105422 3666 105474 3678
rect 105422 3602 105474 3614
rect 109118 3666 109170 3678
rect 109118 3602 109170 3614
rect 112702 3666 112754 3678
rect 112702 3602 112754 3614
rect 116286 3666 116338 3678
rect 116286 3602 116338 3614
rect 119198 3666 119250 3678
rect 119198 3602 119250 3614
rect 119982 3666 120034 3678
rect 119982 3602 120034 3614
rect 182030 3666 182082 3678
rect 182030 3602 182082 3614
rect 182254 3666 182306 3678
rect 182254 3602 182306 3614
rect 196814 3666 196866 3678
rect 196814 3602 196866 3614
rect 198158 3666 198210 3678
rect 198158 3602 198210 3614
rect 204542 3666 204594 3678
rect 204542 3602 204594 3614
rect 205662 3666 205714 3678
rect 205662 3602 205714 3614
rect 206670 3666 206722 3678
rect 206670 3602 206722 3614
rect 208686 3666 208738 3678
rect 215406 3666 215458 3678
rect 209122 3614 209134 3666
rect 209186 3614 209198 3666
rect 211362 3614 211374 3666
rect 211426 3614 211438 3666
rect 208686 3602 208738 3614
rect 215406 3602 215458 3614
rect 222014 3666 222066 3678
rect 267026 3614 267038 3666
rect 267090 3614 267102 3666
rect 270610 3614 270622 3666
rect 270674 3614 270686 3666
rect 281362 3614 281374 3666
rect 281426 3614 281438 3666
rect 288530 3614 288542 3666
rect 288594 3614 288606 3666
rect 292114 3614 292126 3666
rect 292178 3614 292190 3666
rect 222014 3602 222066 3614
rect 78654 3554 78706 3566
rect 182814 3554 182866 3566
rect 195358 3554 195410 3566
rect 203534 3554 203586 3566
rect 205102 3554 205154 3566
rect 11554 3502 11566 3554
rect 11618 3502 11630 3554
rect 43026 3502 43038 3554
rect 43090 3502 43102 3554
rect 46834 3502 46846 3554
rect 46898 3502 46910 3554
rect 50530 3502 50542 3554
rect 50594 3502 50606 3554
rect 54114 3502 54126 3554
rect 54178 3502 54190 3554
rect 57250 3502 57262 3554
rect 57314 3502 57326 3554
rect 60946 3502 60958 3554
rect 61010 3502 61022 3554
rect 65202 3502 65214 3554
rect 65266 3502 65278 3554
rect 68898 3502 68910 3554
rect 68962 3502 68974 3554
rect 72818 3502 72830 3554
rect 72882 3502 72894 3554
rect 74050 3502 74062 3554
rect 74114 3502 74126 3554
rect 89394 3502 89406 3554
rect 89458 3502 89470 3554
rect 94210 3502 94222 3554
rect 94274 3502 94286 3554
rect 97570 3502 97582 3554
rect 97634 3502 97646 3554
rect 103954 3502 103966 3554
rect 104018 3502 104030 3554
rect 107762 3502 107774 3554
rect 107826 3502 107838 3554
rect 111458 3502 111470 3554
rect 111522 3502 111534 3554
rect 115042 3502 115054 3554
rect 115106 3502 115118 3554
rect 118626 3502 118638 3554
rect 118690 3502 118702 3554
rect 122322 3502 122334 3554
rect 122386 3502 122398 3554
rect 183698 3502 183710 3554
rect 183762 3502 183774 3554
rect 185938 3502 185950 3554
rect 186002 3502 186014 3554
rect 188514 3502 188526 3554
rect 188578 3502 188590 3554
rect 193106 3502 193118 3554
rect 193170 3502 193182 3554
rect 193554 3502 193566 3554
rect 193618 3502 193630 3554
rect 194786 3502 194798 3554
rect 194850 3502 194862 3554
rect 201618 3502 201630 3554
rect 201682 3502 201694 3554
rect 202402 3502 202414 3554
rect 202466 3502 202478 3554
rect 202738 3502 202750 3554
rect 202802 3502 202814 3554
rect 203970 3502 203982 3554
rect 204034 3502 204046 3554
rect 78654 3490 78706 3502
rect 182814 3490 182866 3502
rect 195358 3490 195410 3502
rect 203534 3490 203586 3502
rect 205102 3490 205154 3502
rect 205326 3554 205378 3566
rect 205326 3490 205378 3502
rect 205550 3554 205602 3566
rect 208238 3554 208290 3566
rect 210590 3554 210642 3566
rect 212046 3554 212098 3566
rect 220894 3554 220946 3566
rect 285070 3554 285122 3566
rect 206098 3502 206110 3554
rect 206162 3502 206174 3554
rect 207554 3502 207566 3554
rect 207618 3502 207630 3554
rect 209458 3502 209470 3554
rect 209522 3502 209534 3554
rect 210018 3502 210030 3554
rect 210082 3502 210094 3554
rect 211586 3502 211598 3554
rect 211650 3502 211662 3554
rect 213042 3502 213054 3554
rect 213106 3502 213118 3554
rect 216626 3502 216638 3554
rect 216690 3502 216702 3554
rect 220210 3502 220222 3554
rect 220274 3502 220286 3554
rect 223794 3502 223806 3554
rect 223858 3502 223870 3554
rect 227378 3502 227390 3554
rect 227442 3502 227454 3554
rect 230962 3502 230974 3554
rect 231026 3502 231038 3554
rect 234546 3502 234558 3554
rect 234610 3502 234622 3554
rect 238130 3502 238142 3554
rect 238194 3502 238206 3554
rect 241826 3502 241838 3554
rect 241890 3502 241902 3554
rect 245634 3502 245646 3554
rect 245698 3502 245710 3554
rect 249442 3502 249454 3554
rect 249506 3502 249518 3554
rect 253250 3502 253262 3554
rect 253314 3502 253326 3554
rect 256050 3502 256062 3554
rect 256114 3502 256126 3554
rect 259634 3502 259646 3554
rect 259698 3502 259710 3554
rect 263218 3502 263230 3554
rect 263282 3502 263294 3554
rect 205550 3490 205602 3502
rect 208238 3490 208290 3502
rect 210590 3490 210642 3502
rect 212046 3490 212098 3502
rect 220894 3490 220946 3502
rect 285070 3490 285122 3502
rect 78990 3442 79042 3454
rect 10098 3390 10110 3442
rect 10162 3390 10174 3442
rect 75618 3390 75630 3442
rect 75682 3390 75694 3442
rect 78990 3378 79042 3390
rect 89630 3442 89682 3454
rect 89630 3378 89682 3390
rect 104750 3442 104802 3454
rect 104750 3378 104802 3390
rect 108558 3442 108610 3454
rect 108558 3378 108610 3390
rect 123118 3442 123170 3454
rect 123118 3378 123170 3390
rect 123566 3442 123618 3454
rect 126926 3442 126978 3454
rect 123890 3390 123902 3442
rect 123954 3390 123966 3442
rect 123566 3378 123618 3390
rect 126926 3378 126978 3390
rect 127374 3442 127426 3454
rect 130734 3442 130786 3454
rect 127698 3390 127710 3442
rect 127762 3390 127774 3442
rect 127374 3378 127426 3390
rect 130734 3378 130786 3390
rect 131182 3442 131234 3454
rect 133758 3442 133810 3454
rect 131506 3390 131518 3442
rect 131570 3390 131582 3442
rect 131182 3378 131234 3390
rect 133758 3378 133810 3390
rect 133982 3442 134034 3454
rect 137342 3442 137394 3454
rect 134306 3390 134318 3442
rect 134370 3390 134382 3442
rect 133982 3378 134034 3390
rect 137342 3378 137394 3390
rect 137566 3442 137618 3454
rect 140926 3442 140978 3454
rect 137890 3390 137902 3442
rect 137954 3390 137966 3442
rect 137566 3378 137618 3390
rect 140926 3378 140978 3390
rect 141150 3442 141202 3454
rect 144510 3442 144562 3454
rect 141474 3390 141486 3442
rect 141538 3390 141550 3442
rect 141150 3378 141202 3390
rect 144510 3378 144562 3390
rect 144734 3442 144786 3454
rect 148094 3442 148146 3454
rect 145058 3390 145070 3442
rect 145122 3390 145134 3442
rect 144734 3378 144786 3390
rect 148094 3378 148146 3390
rect 148318 3442 148370 3454
rect 148318 3378 148370 3390
rect 148654 3442 148706 3454
rect 148654 3378 148706 3390
rect 151678 3442 151730 3454
rect 151678 3378 151730 3390
rect 151902 3442 151954 3454
rect 155262 3442 155314 3454
rect 152226 3390 152238 3442
rect 152290 3390 152302 3442
rect 151902 3378 151954 3390
rect 155262 3378 155314 3390
rect 155486 3442 155538 3454
rect 158846 3442 158898 3454
rect 155810 3390 155822 3442
rect 155874 3390 155886 3442
rect 155486 3378 155538 3390
rect 158846 3378 158898 3390
rect 159070 3442 159122 3454
rect 162430 3442 162482 3454
rect 159394 3390 159406 3442
rect 159458 3390 159470 3442
rect 159070 3378 159122 3390
rect 162430 3378 162482 3390
rect 162654 3442 162706 3454
rect 162654 3378 162706 3390
rect 166014 3442 166066 3454
rect 166014 3378 166066 3390
rect 166238 3442 166290 3454
rect 169598 3442 169650 3454
rect 166562 3390 166574 3442
rect 166626 3390 166638 3442
rect 166238 3378 166290 3390
rect 169598 3378 169650 3390
rect 169822 3442 169874 3454
rect 172622 3442 172674 3454
rect 170146 3390 170158 3442
rect 170210 3390 170222 3442
rect 169822 3378 169874 3390
rect 172622 3378 172674 3390
rect 173406 3442 173458 3454
rect 173406 3378 173458 3390
rect 173742 3442 173794 3454
rect 173742 3378 173794 3390
rect 176430 3442 176482 3454
rect 176430 3378 176482 3390
rect 176990 3442 177042 3454
rect 176990 3378 177042 3390
rect 180238 3442 180290 3454
rect 180238 3378 180290 3390
rect 180686 3442 180738 3454
rect 183374 3442 183426 3454
rect 187854 3442 187906 3454
rect 190094 3442 190146 3454
rect 181010 3390 181022 3442
rect 181074 3390 181086 3442
rect 183922 3390 183934 3442
rect 183986 3390 183998 3442
rect 184706 3390 184718 3442
rect 184770 3390 184782 3442
rect 188290 3390 188302 3442
rect 188354 3390 188366 3442
rect 180686 3378 180738 3390
rect 183374 3378 183426 3390
rect 187854 3378 187906 3390
rect 190094 3378 190146 3390
rect 190542 3442 190594 3454
rect 190542 3378 190594 3390
rect 190766 3442 190818 3454
rect 190766 3378 190818 3390
rect 190878 3442 190930 3454
rect 190878 3378 190930 3390
rect 191214 3442 191266 3454
rect 195918 3442 195970 3454
rect 197150 3442 197202 3454
rect 191538 3390 191550 3442
rect 191602 3390 191614 3442
rect 196242 3390 196254 3442
rect 196306 3390 196318 3442
rect 191214 3378 191266 3390
rect 195918 3378 195970 3390
rect 197150 3378 197202 3390
rect 197598 3442 197650 3454
rect 197598 3378 197650 3390
rect 198494 3442 198546 3454
rect 198494 3378 198546 3390
rect 198830 3442 198882 3454
rect 198830 3378 198882 3390
rect 199838 3442 199890 3454
rect 199838 3378 199890 3390
rect 200398 3442 200450 3454
rect 200398 3378 200450 3390
rect 200846 3442 200898 3454
rect 200846 3378 200898 3390
rect 201294 3442 201346 3454
rect 201294 3378 201346 3390
rect 201742 3442 201794 3454
rect 201742 3378 201794 3390
rect 203086 3442 203138 3454
rect 203086 3378 203138 3390
rect 204878 3442 204930 3454
rect 207342 3442 207394 3454
rect 205874 3390 205886 3442
rect 205938 3390 205950 3442
rect 204878 3378 204930 3390
rect 207342 3378 207394 3390
rect 209022 3442 209074 3454
rect 209022 3378 209074 3390
rect 209246 3442 209298 3454
rect 209246 3378 209298 3390
rect 209806 3442 209858 3454
rect 209806 3378 209858 3390
rect 211150 3442 211202 3454
rect 211150 3378 211202 3390
rect 211374 3442 211426 3454
rect 211374 3378 211426 3390
rect 212606 3442 212658 3454
rect 212606 3378 212658 3390
rect 212830 3442 212882 3454
rect 212830 3378 212882 3390
rect 219326 3442 219378 3454
rect 219326 3378 219378 3390
rect 219550 3442 219602 3454
rect 219550 3378 219602 3390
rect 219886 3442 219938 3454
rect 219886 3378 219938 3390
rect 220446 3442 220498 3454
rect 220446 3378 220498 3390
rect 220670 3442 220722 3454
rect 220670 3378 220722 3390
rect 221230 3442 221282 3454
rect 221230 3378 221282 3390
rect 221454 3442 221506 3454
rect 221454 3378 221506 3390
rect 223358 3442 223410 3454
rect 223358 3378 223410 3390
rect 226942 3442 226994 3454
rect 226942 3378 226994 3390
rect 230526 3442 230578 3454
rect 230526 3378 230578 3390
rect 233550 3442 233602 3454
rect 233550 3378 233602 3390
rect 237358 3442 237410 3454
rect 237358 3378 237410 3390
rect 241166 3442 241218 3454
rect 241166 3378 241218 3390
rect 244974 3442 245026 3454
rect 244974 3378 245026 3390
rect 245422 3442 245474 3454
rect 245422 3378 245474 3390
rect 248782 3442 248834 3454
rect 248782 3378 248834 3390
rect 249230 3442 249282 3454
rect 249230 3378 249282 3390
rect 252590 3442 252642 3454
rect 252590 3378 252642 3390
rect 255614 3442 255666 3454
rect 255614 3378 255666 3390
rect 259198 3442 259250 3454
rect 259198 3378 259250 3390
rect 262782 3442 262834 3454
rect 262782 3378 262834 3390
rect 266366 3442 266418 3454
rect 266366 3378 266418 3390
rect 266590 3442 266642 3454
rect 266590 3378 266642 3390
rect 269950 3442 270002 3454
rect 269950 3378 270002 3390
rect 270174 3442 270226 3454
rect 270174 3378 270226 3390
rect 273534 3442 273586 3454
rect 273534 3378 273586 3390
rect 273758 3442 273810 3454
rect 273758 3378 273810 3390
rect 274318 3442 274370 3454
rect 274318 3378 274370 3390
rect 277118 3442 277170 3454
rect 277118 3378 277170 3390
rect 277342 3442 277394 3454
rect 277342 3378 277394 3390
rect 277902 3442 277954 3454
rect 277902 3378 277954 3390
rect 280702 3442 280754 3454
rect 280702 3378 280754 3390
rect 280926 3442 280978 3454
rect 280926 3378 280978 3390
rect 284286 3442 284338 3454
rect 284286 3378 284338 3390
rect 284510 3442 284562 3454
rect 284510 3378 284562 3390
rect 287870 3442 287922 3454
rect 287870 3378 287922 3390
rect 288094 3442 288146 3454
rect 288094 3378 288146 3390
rect 291454 3442 291506 3454
rect 291454 3378 291506 3390
rect 291678 3442 291730 3454
rect 291678 3378 291730 3390
rect 12238 3330 12290 3342
rect 12238 3266 12290 3278
rect 15710 3330 15762 3342
rect 15710 3266 15762 3278
rect 19294 3330 19346 3342
rect 19294 3266 19346 3278
rect 22878 3330 22930 3342
rect 22878 3266 22930 3278
rect 26462 3330 26514 3342
rect 26462 3266 26514 3278
rect 30046 3330 30098 3342
rect 30046 3266 30098 3278
rect 33630 3330 33682 3342
rect 33630 3266 33682 3278
rect 37214 3330 37266 3342
rect 37214 3266 37266 3278
rect 94782 3330 94834 3342
rect 94782 3266 94834 3278
rect 98590 3330 98642 3342
rect 177326 3330 177378 3342
rect 186734 3330 186786 3342
rect 215854 3330 215906 3342
rect 162978 3278 162990 3330
rect 163042 3278 163054 3330
rect 184818 3278 184830 3330
rect 184882 3278 184894 3330
rect 193330 3278 193342 3330
rect 193394 3278 193406 3330
rect 98590 3266 98642 3278
rect 177326 3266 177378 3278
rect 186734 3266 186786 3278
rect 215854 3266 215906 3278
rect 216414 3330 216466 3342
rect 216414 3266 216466 3278
rect 223582 3330 223634 3342
rect 223582 3266 223634 3278
rect 227166 3330 227218 3342
rect 227166 3266 227218 3278
rect 230750 3330 230802 3342
rect 230750 3266 230802 3278
rect 234334 3330 234386 3342
rect 234334 3266 234386 3278
rect 237918 3330 237970 3342
rect 237918 3266 237970 3278
rect 241614 3330 241666 3342
rect 241614 3266 241666 3278
rect 253038 3330 253090 3342
rect 253038 3266 253090 3278
rect 255838 3330 255890 3342
rect 259410 3278 259422 3330
rect 259474 3278 259486 3330
rect 262994 3278 263006 3330
rect 263058 3278 263070 3330
rect 255838 3266 255890 3278
rect 1344 3162 298592 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 81278 3162
rect 81330 3110 81382 3162
rect 81434 3110 81486 3162
rect 81538 3110 111998 3162
rect 112050 3110 112102 3162
rect 112154 3110 112206 3162
rect 112258 3110 142718 3162
rect 142770 3110 142822 3162
rect 142874 3110 142926 3162
rect 142978 3110 173438 3162
rect 173490 3110 173542 3162
rect 173594 3110 173646 3162
rect 173698 3110 204158 3162
rect 204210 3110 204262 3162
rect 204314 3110 204366 3162
rect 204418 3110 234878 3162
rect 234930 3110 234982 3162
rect 235034 3110 235086 3162
rect 235138 3110 265598 3162
rect 265650 3110 265702 3162
rect 265754 3110 265806 3162
rect 265858 3110 296318 3162
rect 296370 3110 296422 3162
rect 296474 3110 296526 3162
rect 296578 3110 298592 3162
rect 1344 3076 298592 3110
<< via1 >>
rect 77310 57038 77362 57090
rect 78094 57038 78146 57090
rect 157390 57038 157442 57090
rect 157950 57038 158002 57090
rect 158510 57038 158562 57090
rect 270846 57038 270898 57090
rect 271518 57038 271570 57090
rect 11902 56590 11954 56642
rect 13134 56590 13186 56642
rect 23550 56590 23602 56642
rect 24110 56590 24162 56642
rect 24558 56590 24610 56642
rect 114942 56590 114994 56642
rect 115502 56590 115554 56642
rect 115950 56590 116002 56642
rect 168702 56590 168754 56642
rect 169598 56590 169650 56642
rect 190206 56590 190258 56642
rect 191438 56590 191490 56642
rect 192222 56590 192274 56642
rect 222126 56590 222178 56642
rect 223022 56590 223074 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 81278 56422 81330 56474
rect 81382 56422 81434 56474
rect 81486 56422 81538 56474
rect 111998 56422 112050 56474
rect 112102 56422 112154 56474
rect 112206 56422 112258 56474
rect 142718 56422 142770 56474
rect 142822 56422 142874 56474
rect 142926 56422 142978 56474
rect 173438 56422 173490 56474
rect 173542 56422 173594 56474
rect 173646 56422 173698 56474
rect 204158 56422 204210 56474
rect 204262 56422 204314 56474
rect 204366 56422 204418 56474
rect 234878 56422 234930 56474
rect 234982 56422 235034 56474
rect 235086 56422 235138 56474
rect 265598 56422 265650 56474
rect 265702 56422 265754 56474
rect 265806 56422 265858 56474
rect 296318 56422 296370 56474
rect 296422 56422 296474 56474
rect 296526 56422 296578 56474
rect 12686 56254 12738 56306
rect 18174 56254 18226 56306
rect 18398 56254 18450 56306
rect 19182 56254 19234 56306
rect 24110 56254 24162 56306
rect 24558 56254 24610 56306
rect 28926 56254 28978 56306
rect 29150 56254 29202 56306
rect 34302 56254 34354 56306
rect 34526 56254 34578 56306
rect 39342 56254 39394 56306
rect 39902 56254 39954 56306
rect 45054 56254 45106 56306
rect 45278 56254 45330 56306
rect 50766 56254 50818 56306
rect 51214 56254 51266 56306
rect 55806 56254 55858 56306
rect 56030 56254 56082 56306
rect 61182 56254 61234 56306
rect 61406 56254 61458 56306
rect 109566 56254 109618 56306
rect 109790 56254 109842 56306
rect 115502 56254 115554 56306
rect 115950 56254 116002 56306
rect 120318 56254 120370 56306
rect 120542 56254 120594 56306
rect 125694 56254 125746 56306
rect 125918 56254 125970 56306
rect 130734 56254 130786 56306
rect 136446 56254 136498 56306
rect 142158 56254 142210 56306
rect 147198 56254 147250 56306
rect 152574 56254 152626 56306
rect 157390 56254 157442 56306
rect 163326 56254 163378 56306
rect 168814 56254 168866 56306
rect 174078 56254 174130 56306
rect 179454 56254 179506 56306
rect 184830 56254 184882 56306
rect 192222 56254 192274 56306
rect 195470 56254 195522 56306
rect 208350 56254 208402 56306
rect 211710 56254 211762 56306
rect 211934 56254 211986 56306
rect 217086 56254 217138 56306
rect 222126 56254 222178 56306
rect 223022 56254 223074 56306
rect 227838 56254 227890 56306
rect 233550 56254 233602 56306
rect 238590 56254 238642 56306
rect 238814 56254 238866 56306
rect 243966 56254 244018 56306
rect 244190 56254 244242 56306
rect 248782 56254 248834 56306
rect 249566 56254 249618 56306
rect 254718 56254 254770 56306
rect 260094 56254 260146 56306
rect 265470 56254 265522 56306
rect 271518 56254 271570 56306
rect 276222 56254 276274 56306
rect 286862 56254 286914 56306
rect 287310 56254 287362 56306
rect 292350 56254 292402 56306
rect 292574 56254 292626 56306
rect 13134 56142 13186 56194
rect 126254 56142 126306 56194
rect 131294 56142 131346 56194
rect 131630 56142 131682 56194
rect 136670 56142 136722 56194
rect 142606 56142 142658 56194
rect 147422 56142 147474 56194
rect 152798 56142 152850 56194
rect 153134 56142 153186 56194
rect 158174 56142 158226 56194
rect 158510 56142 158562 56194
rect 163550 56142 163602 56194
rect 169262 56142 169314 56194
rect 169598 56142 169650 56194
rect 174302 56142 174354 56194
rect 179678 56142 179730 56194
rect 180014 56142 180066 56194
rect 185054 56142 185106 56194
rect 189870 56142 189922 56194
rect 191214 56142 191266 56194
rect 195918 56142 195970 56194
rect 212270 56142 212322 56194
rect 217310 56142 217362 56194
rect 222686 56142 222738 56194
rect 228062 56142 228114 56194
rect 233998 56142 234050 56194
rect 13358 56030 13410 56082
rect 69358 56030 69410 56082
rect 80446 56030 80498 56082
rect 84926 56030 84978 56082
rect 85710 56030 85762 56082
rect 91870 56030 91922 56082
rect 92430 56030 92482 56082
rect 96238 56030 96290 56082
rect 107102 56030 107154 56082
rect 107662 56030 107714 56082
rect 136894 56030 136946 56082
rect 142830 56030 142882 56082
rect 147646 56030 147698 56082
rect 163774 56030 163826 56082
rect 174526 56030 174578 56082
rect 185278 56030 185330 56082
rect 190878 56030 190930 56082
rect 191438 56030 191490 56082
rect 196142 56030 196194 56082
rect 202974 56030 203026 56082
rect 206894 56030 206946 56082
rect 207342 56030 207394 56082
rect 217534 56030 217586 56082
rect 228286 56030 228338 56082
rect 234222 56030 234274 56082
rect 254942 56030 254994 56082
rect 260766 56030 260818 56082
rect 265694 56030 265746 56082
rect 272190 56030 272242 56082
rect 276446 56030 276498 56082
rect 282718 56030 282770 56082
rect 283614 56030 283666 56082
rect 25118 55918 25170 55970
rect 29710 55918 29762 55970
rect 35086 55918 35138 55970
rect 40462 55918 40514 55970
rect 45838 55918 45890 55970
rect 51774 55918 51826 55970
rect 56590 55918 56642 55970
rect 61966 55918 62018 55970
rect 67006 55918 67058 55970
rect 70478 55918 70530 55970
rect 78094 55918 78146 55970
rect 81006 55918 81058 55970
rect 82686 55918 82738 55970
rect 89518 55918 89570 55970
rect 93886 55918 93938 55970
rect 97134 55918 97186 55970
rect 104750 55918 104802 55970
rect 110350 55918 110402 55970
rect 116510 55918 116562 55970
rect 121102 55918 121154 55970
rect 187854 55918 187906 55970
rect 188526 55918 188578 55970
rect 189086 55918 189138 55970
rect 200958 55918 201010 55970
rect 203758 55918 203810 55970
rect 239262 55918 239314 55970
rect 244750 55918 244802 55970
rect 250126 55918 250178 55970
rect 256062 55918 256114 55970
rect 261774 55918 261826 55970
rect 266366 55918 266418 55970
rect 273198 55918 273250 55970
rect 277230 55918 277282 55970
rect 281822 55918 281874 55970
rect 288094 55806 288146 55858
rect 293358 55806 293410 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 96638 55638 96690 55690
rect 96742 55638 96794 55690
rect 96846 55638 96898 55690
rect 127358 55638 127410 55690
rect 127462 55638 127514 55690
rect 127566 55638 127618 55690
rect 158078 55638 158130 55690
rect 158182 55638 158234 55690
rect 158286 55638 158338 55690
rect 188798 55638 188850 55690
rect 188902 55638 188954 55690
rect 189006 55638 189058 55690
rect 219518 55638 219570 55690
rect 219622 55638 219674 55690
rect 219726 55638 219778 55690
rect 250238 55638 250290 55690
rect 250342 55638 250394 55690
rect 250446 55638 250498 55690
rect 280958 55638 281010 55690
rect 281062 55638 281114 55690
rect 281166 55638 281218 55690
rect 72382 55358 72434 55410
rect 100046 55358 100098 55410
rect 141262 55358 141314 55410
rect 156270 55358 156322 55410
rect 161870 55358 161922 55410
rect 180238 55358 180290 55410
rect 182366 55358 182418 55410
rect 186174 55358 186226 55410
rect 186398 55358 186450 55410
rect 188302 55358 188354 55410
rect 190430 55358 190482 55410
rect 74734 55246 74786 55298
rect 102286 55246 102338 55298
rect 135102 55246 135154 55298
rect 138350 55246 138402 55298
rect 140478 55246 140530 55298
rect 143838 55246 143890 55298
rect 152686 55246 152738 55298
rect 156718 55246 156770 55298
rect 162430 55246 162482 55298
rect 169710 55246 169762 55298
rect 170382 55246 170434 55298
rect 174974 55246 175026 55298
rect 175534 55246 175586 55298
rect 179454 55246 179506 55298
rect 186062 55246 186114 55298
rect 187182 55246 187234 55298
rect 191214 55246 191266 55298
rect 135774 55134 135826 55186
rect 147870 55134 147922 55186
rect 157390 55134 157442 55186
rect 163214 55134 163266 55186
rect 168926 55134 168978 55186
rect 174302 55134 174354 55186
rect 186510 55134 186562 55186
rect 186846 55134 186898 55186
rect 186958 55134 187010 55186
rect 187518 55134 187570 55186
rect 75182 55022 75234 55074
rect 102734 55022 102786 55074
rect 153246 55022 153298 55074
rect 182814 55022 182866 55074
rect 187966 55022 188018 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 81278 54854 81330 54906
rect 81382 54854 81434 54906
rect 81486 54854 81538 54906
rect 111998 54854 112050 54906
rect 112102 54854 112154 54906
rect 112206 54854 112258 54906
rect 142718 54854 142770 54906
rect 142822 54854 142874 54906
rect 142926 54854 142978 54906
rect 173438 54854 173490 54906
rect 173542 54854 173594 54906
rect 173646 54854 173698 54906
rect 204158 54854 204210 54906
rect 204262 54854 204314 54906
rect 204366 54854 204418 54906
rect 234878 54854 234930 54906
rect 234982 54854 235034 54906
rect 235086 54854 235138 54906
rect 265598 54854 265650 54906
rect 265702 54854 265754 54906
rect 265806 54854 265858 54906
rect 296318 54854 296370 54906
rect 296422 54854 296474 54906
rect 296526 54854 296578 54906
rect 132974 54686 133026 54738
rect 135774 54686 135826 54738
rect 141038 54686 141090 54738
rect 148654 54686 148706 54738
rect 150110 54686 150162 54738
rect 157166 54686 157218 54738
rect 162318 54686 162370 54738
rect 167918 54686 167970 54738
rect 172734 54686 172786 54738
rect 184046 54574 184098 54626
rect 193902 54574 193954 54626
rect 132526 54462 132578 54514
rect 148094 54462 148146 54514
rect 153918 54462 153970 54514
rect 183262 54462 183314 54514
rect 191438 54462 191490 54514
rect 194574 54462 194626 54514
rect 131742 54350 131794 54402
rect 147422 54350 147474 54402
rect 153134 54350 153186 54402
rect 182926 54350 182978 54402
rect 186174 54350 186226 54402
rect 191774 54350 191826 54402
rect 134990 54238 135042 54290
rect 140254 54238 140306 54290
rect 156382 54238 156434 54290
rect 161534 54238 161586 54290
rect 167134 54238 167186 54290
rect 171950 54238 172002 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 96638 54070 96690 54122
rect 96742 54070 96794 54122
rect 96846 54070 96898 54122
rect 127358 54070 127410 54122
rect 127462 54070 127514 54122
rect 127566 54070 127618 54122
rect 158078 54070 158130 54122
rect 158182 54070 158234 54122
rect 158286 54070 158338 54122
rect 188798 54070 188850 54122
rect 188902 54070 188954 54122
rect 189006 54070 189058 54122
rect 219518 54070 219570 54122
rect 219622 54070 219674 54122
rect 219726 54070 219778 54122
rect 250238 54070 250290 54122
rect 250342 54070 250394 54122
rect 250446 54070 250498 54122
rect 280958 54070 281010 54122
rect 281062 54070 281114 54122
rect 281166 54070 281218 54122
rect 180126 53790 180178 53842
rect 193230 53790 193282 53842
rect 130286 53678 130338 53730
rect 145966 53678 146018 53730
rect 151566 53678 151618 53730
rect 161982 53678 162034 53730
rect 162430 53678 162482 53730
rect 178110 53678 178162 53730
rect 189758 53678 189810 53730
rect 190430 53678 190482 53730
rect 129390 53566 129442 53618
rect 167470 53566 167522 53618
rect 177662 53566 177714 53618
rect 191102 53566 191154 53618
rect 145182 53454 145234 53506
rect 150782 53454 150834 53506
rect 189422 53454 189474 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 81278 53286 81330 53338
rect 81382 53286 81434 53338
rect 81486 53286 81538 53338
rect 111998 53286 112050 53338
rect 112102 53286 112154 53338
rect 112206 53286 112258 53338
rect 142718 53286 142770 53338
rect 142822 53286 142874 53338
rect 142926 53286 142978 53338
rect 173438 53286 173490 53338
rect 173542 53286 173594 53338
rect 173646 53286 173698 53338
rect 204158 53286 204210 53338
rect 204262 53286 204314 53338
rect 204366 53286 204418 53338
rect 234878 53286 234930 53338
rect 234982 53286 235034 53338
rect 235086 53286 235138 53338
rect 265598 53286 265650 53338
rect 265702 53286 265754 53338
rect 265806 53286 265858 53338
rect 296318 53286 296370 53338
rect 296422 53286 296474 53338
rect 296526 53286 296578 53338
rect 182142 53118 182194 53170
rect 185838 53118 185890 53170
rect 182478 52894 182530 52946
rect 186510 52894 186562 52946
rect 181470 52782 181522 52834
rect 183262 52782 183314 52834
rect 185390 52782 185442 52834
rect 187182 52782 187234 52834
rect 189310 52782 189362 52834
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 96638 52502 96690 52554
rect 96742 52502 96794 52554
rect 96846 52502 96898 52554
rect 127358 52502 127410 52554
rect 127462 52502 127514 52554
rect 127566 52502 127618 52554
rect 158078 52502 158130 52554
rect 158182 52502 158234 52554
rect 158286 52502 158338 52554
rect 188798 52502 188850 52554
rect 188902 52502 188954 52554
rect 189006 52502 189058 52554
rect 219518 52502 219570 52554
rect 219622 52502 219674 52554
rect 219726 52502 219778 52554
rect 250238 52502 250290 52554
rect 250342 52502 250394 52554
rect 250446 52502 250498 52554
rect 280958 52502 281010 52554
rect 281062 52502 281114 52554
rect 281166 52502 281218 52554
rect 186174 52222 186226 52274
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 81278 51718 81330 51770
rect 81382 51718 81434 51770
rect 81486 51718 81538 51770
rect 111998 51718 112050 51770
rect 112102 51718 112154 51770
rect 112206 51718 112258 51770
rect 142718 51718 142770 51770
rect 142822 51718 142874 51770
rect 142926 51718 142978 51770
rect 173438 51718 173490 51770
rect 173542 51718 173594 51770
rect 173646 51718 173698 51770
rect 204158 51718 204210 51770
rect 204262 51718 204314 51770
rect 204366 51718 204418 51770
rect 234878 51718 234930 51770
rect 234982 51718 235034 51770
rect 235086 51718 235138 51770
rect 265598 51718 265650 51770
rect 265702 51718 265754 51770
rect 265806 51718 265858 51770
rect 296318 51718 296370 51770
rect 296422 51718 296474 51770
rect 296526 51718 296578 51770
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 96638 50934 96690 50986
rect 96742 50934 96794 50986
rect 96846 50934 96898 50986
rect 127358 50934 127410 50986
rect 127462 50934 127514 50986
rect 127566 50934 127618 50986
rect 158078 50934 158130 50986
rect 158182 50934 158234 50986
rect 158286 50934 158338 50986
rect 188798 50934 188850 50986
rect 188902 50934 188954 50986
rect 189006 50934 189058 50986
rect 219518 50934 219570 50986
rect 219622 50934 219674 50986
rect 219726 50934 219778 50986
rect 250238 50934 250290 50986
rect 250342 50934 250394 50986
rect 250446 50934 250498 50986
rect 280958 50934 281010 50986
rect 281062 50934 281114 50986
rect 281166 50934 281218 50986
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 81278 50150 81330 50202
rect 81382 50150 81434 50202
rect 81486 50150 81538 50202
rect 111998 50150 112050 50202
rect 112102 50150 112154 50202
rect 112206 50150 112258 50202
rect 142718 50150 142770 50202
rect 142822 50150 142874 50202
rect 142926 50150 142978 50202
rect 173438 50150 173490 50202
rect 173542 50150 173594 50202
rect 173646 50150 173698 50202
rect 204158 50150 204210 50202
rect 204262 50150 204314 50202
rect 204366 50150 204418 50202
rect 234878 50150 234930 50202
rect 234982 50150 235034 50202
rect 235086 50150 235138 50202
rect 265598 50150 265650 50202
rect 265702 50150 265754 50202
rect 265806 50150 265858 50202
rect 296318 50150 296370 50202
rect 296422 50150 296474 50202
rect 296526 50150 296578 50202
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 96638 49366 96690 49418
rect 96742 49366 96794 49418
rect 96846 49366 96898 49418
rect 127358 49366 127410 49418
rect 127462 49366 127514 49418
rect 127566 49366 127618 49418
rect 158078 49366 158130 49418
rect 158182 49366 158234 49418
rect 158286 49366 158338 49418
rect 188798 49366 188850 49418
rect 188902 49366 188954 49418
rect 189006 49366 189058 49418
rect 219518 49366 219570 49418
rect 219622 49366 219674 49418
rect 219726 49366 219778 49418
rect 250238 49366 250290 49418
rect 250342 49366 250394 49418
rect 250446 49366 250498 49418
rect 280958 49366 281010 49418
rect 281062 49366 281114 49418
rect 281166 49366 281218 49418
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 81278 48582 81330 48634
rect 81382 48582 81434 48634
rect 81486 48582 81538 48634
rect 111998 48582 112050 48634
rect 112102 48582 112154 48634
rect 112206 48582 112258 48634
rect 142718 48582 142770 48634
rect 142822 48582 142874 48634
rect 142926 48582 142978 48634
rect 173438 48582 173490 48634
rect 173542 48582 173594 48634
rect 173646 48582 173698 48634
rect 204158 48582 204210 48634
rect 204262 48582 204314 48634
rect 204366 48582 204418 48634
rect 234878 48582 234930 48634
rect 234982 48582 235034 48634
rect 235086 48582 235138 48634
rect 265598 48582 265650 48634
rect 265702 48582 265754 48634
rect 265806 48582 265858 48634
rect 296318 48582 296370 48634
rect 296422 48582 296474 48634
rect 296526 48582 296578 48634
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 96638 47798 96690 47850
rect 96742 47798 96794 47850
rect 96846 47798 96898 47850
rect 127358 47798 127410 47850
rect 127462 47798 127514 47850
rect 127566 47798 127618 47850
rect 158078 47798 158130 47850
rect 158182 47798 158234 47850
rect 158286 47798 158338 47850
rect 188798 47798 188850 47850
rect 188902 47798 188954 47850
rect 189006 47798 189058 47850
rect 219518 47798 219570 47850
rect 219622 47798 219674 47850
rect 219726 47798 219778 47850
rect 250238 47798 250290 47850
rect 250342 47798 250394 47850
rect 250446 47798 250498 47850
rect 280958 47798 281010 47850
rect 281062 47798 281114 47850
rect 281166 47798 281218 47850
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 81278 47014 81330 47066
rect 81382 47014 81434 47066
rect 81486 47014 81538 47066
rect 111998 47014 112050 47066
rect 112102 47014 112154 47066
rect 112206 47014 112258 47066
rect 142718 47014 142770 47066
rect 142822 47014 142874 47066
rect 142926 47014 142978 47066
rect 173438 47014 173490 47066
rect 173542 47014 173594 47066
rect 173646 47014 173698 47066
rect 204158 47014 204210 47066
rect 204262 47014 204314 47066
rect 204366 47014 204418 47066
rect 234878 47014 234930 47066
rect 234982 47014 235034 47066
rect 235086 47014 235138 47066
rect 265598 47014 265650 47066
rect 265702 47014 265754 47066
rect 265806 47014 265858 47066
rect 296318 47014 296370 47066
rect 296422 47014 296474 47066
rect 296526 47014 296578 47066
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 96638 46230 96690 46282
rect 96742 46230 96794 46282
rect 96846 46230 96898 46282
rect 127358 46230 127410 46282
rect 127462 46230 127514 46282
rect 127566 46230 127618 46282
rect 158078 46230 158130 46282
rect 158182 46230 158234 46282
rect 158286 46230 158338 46282
rect 188798 46230 188850 46282
rect 188902 46230 188954 46282
rect 189006 46230 189058 46282
rect 219518 46230 219570 46282
rect 219622 46230 219674 46282
rect 219726 46230 219778 46282
rect 250238 46230 250290 46282
rect 250342 46230 250394 46282
rect 250446 46230 250498 46282
rect 280958 46230 281010 46282
rect 281062 46230 281114 46282
rect 281166 46230 281218 46282
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 81278 45446 81330 45498
rect 81382 45446 81434 45498
rect 81486 45446 81538 45498
rect 111998 45446 112050 45498
rect 112102 45446 112154 45498
rect 112206 45446 112258 45498
rect 142718 45446 142770 45498
rect 142822 45446 142874 45498
rect 142926 45446 142978 45498
rect 173438 45446 173490 45498
rect 173542 45446 173594 45498
rect 173646 45446 173698 45498
rect 204158 45446 204210 45498
rect 204262 45446 204314 45498
rect 204366 45446 204418 45498
rect 234878 45446 234930 45498
rect 234982 45446 235034 45498
rect 235086 45446 235138 45498
rect 265598 45446 265650 45498
rect 265702 45446 265754 45498
rect 265806 45446 265858 45498
rect 296318 45446 296370 45498
rect 296422 45446 296474 45498
rect 296526 45446 296578 45498
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 96638 44662 96690 44714
rect 96742 44662 96794 44714
rect 96846 44662 96898 44714
rect 127358 44662 127410 44714
rect 127462 44662 127514 44714
rect 127566 44662 127618 44714
rect 158078 44662 158130 44714
rect 158182 44662 158234 44714
rect 158286 44662 158338 44714
rect 188798 44662 188850 44714
rect 188902 44662 188954 44714
rect 189006 44662 189058 44714
rect 219518 44662 219570 44714
rect 219622 44662 219674 44714
rect 219726 44662 219778 44714
rect 250238 44662 250290 44714
rect 250342 44662 250394 44714
rect 250446 44662 250498 44714
rect 280958 44662 281010 44714
rect 281062 44662 281114 44714
rect 281166 44662 281218 44714
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 81278 43878 81330 43930
rect 81382 43878 81434 43930
rect 81486 43878 81538 43930
rect 111998 43878 112050 43930
rect 112102 43878 112154 43930
rect 112206 43878 112258 43930
rect 142718 43878 142770 43930
rect 142822 43878 142874 43930
rect 142926 43878 142978 43930
rect 173438 43878 173490 43930
rect 173542 43878 173594 43930
rect 173646 43878 173698 43930
rect 204158 43878 204210 43930
rect 204262 43878 204314 43930
rect 204366 43878 204418 43930
rect 234878 43878 234930 43930
rect 234982 43878 235034 43930
rect 235086 43878 235138 43930
rect 265598 43878 265650 43930
rect 265702 43878 265754 43930
rect 265806 43878 265858 43930
rect 296318 43878 296370 43930
rect 296422 43878 296474 43930
rect 296526 43878 296578 43930
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 96638 43094 96690 43146
rect 96742 43094 96794 43146
rect 96846 43094 96898 43146
rect 127358 43094 127410 43146
rect 127462 43094 127514 43146
rect 127566 43094 127618 43146
rect 158078 43094 158130 43146
rect 158182 43094 158234 43146
rect 158286 43094 158338 43146
rect 188798 43094 188850 43146
rect 188902 43094 188954 43146
rect 189006 43094 189058 43146
rect 219518 43094 219570 43146
rect 219622 43094 219674 43146
rect 219726 43094 219778 43146
rect 250238 43094 250290 43146
rect 250342 43094 250394 43146
rect 250446 43094 250498 43146
rect 280958 43094 281010 43146
rect 281062 43094 281114 43146
rect 281166 43094 281218 43146
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 81278 42310 81330 42362
rect 81382 42310 81434 42362
rect 81486 42310 81538 42362
rect 111998 42310 112050 42362
rect 112102 42310 112154 42362
rect 112206 42310 112258 42362
rect 142718 42310 142770 42362
rect 142822 42310 142874 42362
rect 142926 42310 142978 42362
rect 173438 42310 173490 42362
rect 173542 42310 173594 42362
rect 173646 42310 173698 42362
rect 204158 42310 204210 42362
rect 204262 42310 204314 42362
rect 204366 42310 204418 42362
rect 234878 42310 234930 42362
rect 234982 42310 235034 42362
rect 235086 42310 235138 42362
rect 265598 42310 265650 42362
rect 265702 42310 265754 42362
rect 265806 42310 265858 42362
rect 296318 42310 296370 42362
rect 296422 42310 296474 42362
rect 296526 42310 296578 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 96638 41526 96690 41578
rect 96742 41526 96794 41578
rect 96846 41526 96898 41578
rect 127358 41526 127410 41578
rect 127462 41526 127514 41578
rect 127566 41526 127618 41578
rect 158078 41526 158130 41578
rect 158182 41526 158234 41578
rect 158286 41526 158338 41578
rect 188798 41526 188850 41578
rect 188902 41526 188954 41578
rect 189006 41526 189058 41578
rect 219518 41526 219570 41578
rect 219622 41526 219674 41578
rect 219726 41526 219778 41578
rect 250238 41526 250290 41578
rect 250342 41526 250394 41578
rect 250446 41526 250498 41578
rect 280958 41526 281010 41578
rect 281062 41526 281114 41578
rect 281166 41526 281218 41578
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 81278 40742 81330 40794
rect 81382 40742 81434 40794
rect 81486 40742 81538 40794
rect 111998 40742 112050 40794
rect 112102 40742 112154 40794
rect 112206 40742 112258 40794
rect 142718 40742 142770 40794
rect 142822 40742 142874 40794
rect 142926 40742 142978 40794
rect 173438 40742 173490 40794
rect 173542 40742 173594 40794
rect 173646 40742 173698 40794
rect 204158 40742 204210 40794
rect 204262 40742 204314 40794
rect 204366 40742 204418 40794
rect 234878 40742 234930 40794
rect 234982 40742 235034 40794
rect 235086 40742 235138 40794
rect 265598 40742 265650 40794
rect 265702 40742 265754 40794
rect 265806 40742 265858 40794
rect 296318 40742 296370 40794
rect 296422 40742 296474 40794
rect 296526 40742 296578 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 96638 39958 96690 40010
rect 96742 39958 96794 40010
rect 96846 39958 96898 40010
rect 127358 39958 127410 40010
rect 127462 39958 127514 40010
rect 127566 39958 127618 40010
rect 158078 39958 158130 40010
rect 158182 39958 158234 40010
rect 158286 39958 158338 40010
rect 188798 39958 188850 40010
rect 188902 39958 188954 40010
rect 189006 39958 189058 40010
rect 219518 39958 219570 40010
rect 219622 39958 219674 40010
rect 219726 39958 219778 40010
rect 250238 39958 250290 40010
rect 250342 39958 250394 40010
rect 250446 39958 250498 40010
rect 280958 39958 281010 40010
rect 281062 39958 281114 40010
rect 281166 39958 281218 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 81278 39174 81330 39226
rect 81382 39174 81434 39226
rect 81486 39174 81538 39226
rect 111998 39174 112050 39226
rect 112102 39174 112154 39226
rect 112206 39174 112258 39226
rect 142718 39174 142770 39226
rect 142822 39174 142874 39226
rect 142926 39174 142978 39226
rect 173438 39174 173490 39226
rect 173542 39174 173594 39226
rect 173646 39174 173698 39226
rect 204158 39174 204210 39226
rect 204262 39174 204314 39226
rect 204366 39174 204418 39226
rect 234878 39174 234930 39226
rect 234982 39174 235034 39226
rect 235086 39174 235138 39226
rect 265598 39174 265650 39226
rect 265702 39174 265754 39226
rect 265806 39174 265858 39226
rect 296318 39174 296370 39226
rect 296422 39174 296474 39226
rect 296526 39174 296578 39226
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 96638 38390 96690 38442
rect 96742 38390 96794 38442
rect 96846 38390 96898 38442
rect 127358 38390 127410 38442
rect 127462 38390 127514 38442
rect 127566 38390 127618 38442
rect 158078 38390 158130 38442
rect 158182 38390 158234 38442
rect 158286 38390 158338 38442
rect 188798 38390 188850 38442
rect 188902 38390 188954 38442
rect 189006 38390 189058 38442
rect 219518 38390 219570 38442
rect 219622 38390 219674 38442
rect 219726 38390 219778 38442
rect 250238 38390 250290 38442
rect 250342 38390 250394 38442
rect 250446 38390 250498 38442
rect 280958 38390 281010 38442
rect 281062 38390 281114 38442
rect 281166 38390 281218 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 81278 37606 81330 37658
rect 81382 37606 81434 37658
rect 81486 37606 81538 37658
rect 111998 37606 112050 37658
rect 112102 37606 112154 37658
rect 112206 37606 112258 37658
rect 142718 37606 142770 37658
rect 142822 37606 142874 37658
rect 142926 37606 142978 37658
rect 173438 37606 173490 37658
rect 173542 37606 173594 37658
rect 173646 37606 173698 37658
rect 204158 37606 204210 37658
rect 204262 37606 204314 37658
rect 204366 37606 204418 37658
rect 234878 37606 234930 37658
rect 234982 37606 235034 37658
rect 235086 37606 235138 37658
rect 265598 37606 265650 37658
rect 265702 37606 265754 37658
rect 265806 37606 265858 37658
rect 296318 37606 296370 37658
rect 296422 37606 296474 37658
rect 296526 37606 296578 37658
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 96638 36822 96690 36874
rect 96742 36822 96794 36874
rect 96846 36822 96898 36874
rect 127358 36822 127410 36874
rect 127462 36822 127514 36874
rect 127566 36822 127618 36874
rect 158078 36822 158130 36874
rect 158182 36822 158234 36874
rect 158286 36822 158338 36874
rect 188798 36822 188850 36874
rect 188902 36822 188954 36874
rect 189006 36822 189058 36874
rect 219518 36822 219570 36874
rect 219622 36822 219674 36874
rect 219726 36822 219778 36874
rect 250238 36822 250290 36874
rect 250342 36822 250394 36874
rect 250446 36822 250498 36874
rect 280958 36822 281010 36874
rect 281062 36822 281114 36874
rect 281166 36822 281218 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 81278 36038 81330 36090
rect 81382 36038 81434 36090
rect 81486 36038 81538 36090
rect 111998 36038 112050 36090
rect 112102 36038 112154 36090
rect 112206 36038 112258 36090
rect 142718 36038 142770 36090
rect 142822 36038 142874 36090
rect 142926 36038 142978 36090
rect 173438 36038 173490 36090
rect 173542 36038 173594 36090
rect 173646 36038 173698 36090
rect 204158 36038 204210 36090
rect 204262 36038 204314 36090
rect 204366 36038 204418 36090
rect 234878 36038 234930 36090
rect 234982 36038 235034 36090
rect 235086 36038 235138 36090
rect 265598 36038 265650 36090
rect 265702 36038 265754 36090
rect 265806 36038 265858 36090
rect 296318 36038 296370 36090
rect 296422 36038 296474 36090
rect 296526 36038 296578 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 96638 35254 96690 35306
rect 96742 35254 96794 35306
rect 96846 35254 96898 35306
rect 127358 35254 127410 35306
rect 127462 35254 127514 35306
rect 127566 35254 127618 35306
rect 158078 35254 158130 35306
rect 158182 35254 158234 35306
rect 158286 35254 158338 35306
rect 188798 35254 188850 35306
rect 188902 35254 188954 35306
rect 189006 35254 189058 35306
rect 219518 35254 219570 35306
rect 219622 35254 219674 35306
rect 219726 35254 219778 35306
rect 250238 35254 250290 35306
rect 250342 35254 250394 35306
rect 250446 35254 250498 35306
rect 280958 35254 281010 35306
rect 281062 35254 281114 35306
rect 281166 35254 281218 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 81278 34470 81330 34522
rect 81382 34470 81434 34522
rect 81486 34470 81538 34522
rect 111998 34470 112050 34522
rect 112102 34470 112154 34522
rect 112206 34470 112258 34522
rect 142718 34470 142770 34522
rect 142822 34470 142874 34522
rect 142926 34470 142978 34522
rect 173438 34470 173490 34522
rect 173542 34470 173594 34522
rect 173646 34470 173698 34522
rect 204158 34470 204210 34522
rect 204262 34470 204314 34522
rect 204366 34470 204418 34522
rect 234878 34470 234930 34522
rect 234982 34470 235034 34522
rect 235086 34470 235138 34522
rect 265598 34470 265650 34522
rect 265702 34470 265754 34522
rect 265806 34470 265858 34522
rect 296318 34470 296370 34522
rect 296422 34470 296474 34522
rect 296526 34470 296578 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 96638 33686 96690 33738
rect 96742 33686 96794 33738
rect 96846 33686 96898 33738
rect 127358 33686 127410 33738
rect 127462 33686 127514 33738
rect 127566 33686 127618 33738
rect 158078 33686 158130 33738
rect 158182 33686 158234 33738
rect 158286 33686 158338 33738
rect 188798 33686 188850 33738
rect 188902 33686 188954 33738
rect 189006 33686 189058 33738
rect 219518 33686 219570 33738
rect 219622 33686 219674 33738
rect 219726 33686 219778 33738
rect 250238 33686 250290 33738
rect 250342 33686 250394 33738
rect 250446 33686 250498 33738
rect 280958 33686 281010 33738
rect 281062 33686 281114 33738
rect 281166 33686 281218 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 81278 32902 81330 32954
rect 81382 32902 81434 32954
rect 81486 32902 81538 32954
rect 111998 32902 112050 32954
rect 112102 32902 112154 32954
rect 112206 32902 112258 32954
rect 142718 32902 142770 32954
rect 142822 32902 142874 32954
rect 142926 32902 142978 32954
rect 173438 32902 173490 32954
rect 173542 32902 173594 32954
rect 173646 32902 173698 32954
rect 204158 32902 204210 32954
rect 204262 32902 204314 32954
rect 204366 32902 204418 32954
rect 234878 32902 234930 32954
rect 234982 32902 235034 32954
rect 235086 32902 235138 32954
rect 265598 32902 265650 32954
rect 265702 32902 265754 32954
rect 265806 32902 265858 32954
rect 296318 32902 296370 32954
rect 296422 32902 296474 32954
rect 296526 32902 296578 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 96638 32118 96690 32170
rect 96742 32118 96794 32170
rect 96846 32118 96898 32170
rect 127358 32118 127410 32170
rect 127462 32118 127514 32170
rect 127566 32118 127618 32170
rect 158078 32118 158130 32170
rect 158182 32118 158234 32170
rect 158286 32118 158338 32170
rect 188798 32118 188850 32170
rect 188902 32118 188954 32170
rect 189006 32118 189058 32170
rect 219518 32118 219570 32170
rect 219622 32118 219674 32170
rect 219726 32118 219778 32170
rect 250238 32118 250290 32170
rect 250342 32118 250394 32170
rect 250446 32118 250498 32170
rect 280958 32118 281010 32170
rect 281062 32118 281114 32170
rect 281166 32118 281218 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 81278 31334 81330 31386
rect 81382 31334 81434 31386
rect 81486 31334 81538 31386
rect 111998 31334 112050 31386
rect 112102 31334 112154 31386
rect 112206 31334 112258 31386
rect 142718 31334 142770 31386
rect 142822 31334 142874 31386
rect 142926 31334 142978 31386
rect 173438 31334 173490 31386
rect 173542 31334 173594 31386
rect 173646 31334 173698 31386
rect 204158 31334 204210 31386
rect 204262 31334 204314 31386
rect 204366 31334 204418 31386
rect 234878 31334 234930 31386
rect 234982 31334 235034 31386
rect 235086 31334 235138 31386
rect 265598 31334 265650 31386
rect 265702 31334 265754 31386
rect 265806 31334 265858 31386
rect 296318 31334 296370 31386
rect 296422 31334 296474 31386
rect 296526 31334 296578 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 96638 30550 96690 30602
rect 96742 30550 96794 30602
rect 96846 30550 96898 30602
rect 127358 30550 127410 30602
rect 127462 30550 127514 30602
rect 127566 30550 127618 30602
rect 158078 30550 158130 30602
rect 158182 30550 158234 30602
rect 158286 30550 158338 30602
rect 188798 30550 188850 30602
rect 188902 30550 188954 30602
rect 189006 30550 189058 30602
rect 219518 30550 219570 30602
rect 219622 30550 219674 30602
rect 219726 30550 219778 30602
rect 250238 30550 250290 30602
rect 250342 30550 250394 30602
rect 250446 30550 250498 30602
rect 280958 30550 281010 30602
rect 281062 30550 281114 30602
rect 281166 30550 281218 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 81278 29766 81330 29818
rect 81382 29766 81434 29818
rect 81486 29766 81538 29818
rect 111998 29766 112050 29818
rect 112102 29766 112154 29818
rect 112206 29766 112258 29818
rect 142718 29766 142770 29818
rect 142822 29766 142874 29818
rect 142926 29766 142978 29818
rect 173438 29766 173490 29818
rect 173542 29766 173594 29818
rect 173646 29766 173698 29818
rect 204158 29766 204210 29818
rect 204262 29766 204314 29818
rect 204366 29766 204418 29818
rect 234878 29766 234930 29818
rect 234982 29766 235034 29818
rect 235086 29766 235138 29818
rect 265598 29766 265650 29818
rect 265702 29766 265754 29818
rect 265806 29766 265858 29818
rect 296318 29766 296370 29818
rect 296422 29766 296474 29818
rect 296526 29766 296578 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 96638 28982 96690 29034
rect 96742 28982 96794 29034
rect 96846 28982 96898 29034
rect 127358 28982 127410 29034
rect 127462 28982 127514 29034
rect 127566 28982 127618 29034
rect 158078 28982 158130 29034
rect 158182 28982 158234 29034
rect 158286 28982 158338 29034
rect 188798 28982 188850 29034
rect 188902 28982 188954 29034
rect 189006 28982 189058 29034
rect 219518 28982 219570 29034
rect 219622 28982 219674 29034
rect 219726 28982 219778 29034
rect 250238 28982 250290 29034
rect 250342 28982 250394 29034
rect 250446 28982 250498 29034
rect 280958 28982 281010 29034
rect 281062 28982 281114 29034
rect 281166 28982 281218 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 81278 28198 81330 28250
rect 81382 28198 81434 28250
rect 81486 28198 81538 28250
rect 111998 28198 112050 28250
rect 112102 28198 112154 28250
rect 112206 28198 112258 28250
rect 142718 28198 142770 28250
rect 142822 28198 142874 28250
rect 142926 28198 142978 28250
rect 173438 28198 173490 28250
rect 173542 28198 173594 28250
rect 173646 28198 173698 28250
rect 204158 28198 204210 28250
rect 204262 28198 204314 28250
rect 204366 28198 204418 28250
rect 234878 28198 234930 28250
rect 234982 28198 235034 28250
rect 235086 28198 235138 28250
rect 265598 28198 265650 28250
rect 265702 28198 265754 28250
rect 265806 28198 265858 28250
rect 296318 28198 296370 28250
rect 296422 28198 296474 28250
rect 296526 28198 296578 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 96638 27414 96690 27466
rect 96742 27414 96794 27466
rect 96846 27414 96898 27466
rect 127358 27414 127410 27466
rect 127462 27414 127514 27466
rect 127566 27414 127618 27466
rect 158078 27414 158130 27466
rect 158182 27414 158234 27466
rect 158286 27414 158338 27466
rect 188798 27414 188850 27466
rect 188902 27414 188954 27466
rect 189006 27414 189058 27466
rect 219518 27414 219570 27466
rect 219622 27414 219674 27466
rect 219726 27414 219778 27466
rect 250238 27414 250290 27466
rect 250342 27414 250394 27466
rect 250446 27414 250498 27466
rect 280958 27414 281010 27466
rect 281062 27414 281114 27466
rect 281166 27414 281218 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 81278 26630 81330 26682
rect 81382 26630 81434 26682
rect 81486 26630 81538 26682
rect 111998 26630 112050 26682
rect 112102 26630 112154 26682
rect 112206 26630 112258 26682
rect 142718 26630 142770 26682
rect 142822 26630 142874 26682
rect 142926 26630 142978 26682
rect 173438 26630 173490 26682
rect 173542 26630 173594 26682
rect 173646 26630 173698 26682
rect 204158 26630 204210 26682
rect 204262 26630 204314 26682
rect 204366 26630 204418 26682
rect 234878 26630 234930 26682
rect 234982 26630 235034 26682
rect 235086 26630 235138 26682
rect 265598 26630 265650 26682
rect 265702 26630 265754 26682
rect 265806 26630 265858 26682
rect 296318 26630 296370 26682
rect 296422 26630 296474 26682
rect 296526 26630 296578 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 96638 25846 96690 25898
rect 96742 25846 96794 25898
rect 96846 25846 96898 25898
rect 127358 25846 127410 25898
rect 127462 25846 127514 25898
rect 127566 25846 127618 25898
rect 158078 25846 158130 25898
rect 158182 25846 158234 25898
rect 158286 25846 158338 25898
rect 188798 25846 188850 25898
rect 188902 25846 188954 25898
rect 189006 25846 189058 25898
rect 219518 25846 219570 25898
rect 219622 25846 219674 25898
rect 219726 25846 219778 25898
rect 250238 25846 250290 25898
rect 250342 25846 250394 25898
rect 250446 25846 250498 25898
rect 280958 25846 281010 25898
rect 281062 25846 281114 25898
rect 281166 25846 281218 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 81278 25062 81330 25114
rect 81382 25062 81434 25114
rect 81486 25062 81538 25114
rect 111998 25062 112050 25114
rect 112102 25062 112154 25114
rect 112206 25062 112258 25114
rect 142718 25062 142770 25114
rect 142822 25062 142874 25114
rect 142926 25062 142978 25114
rect 173438 25062 173490 25114
rect 173542 25062 173594 25114
rect 173646 25062 173698 25114
rect 204158 25062 204210 25114
rect 204262 25062 204314 25114
rect 204366 25062 204418 25114
rect 234878 25062 234930 25114
rect 234982 25062 235034 25114
rect 235086 25062 235138 25114
rect 265598 25062 265650 25114
rect 265702 25062 265754 25114
rect 265806 25062 265858 25114
rect 296318 25062 296370 25114
rect 296422 25062 296474 25114
rect 296526 25062 296578 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 96638 24278 96690 24330
rect 96742 24278 96794 24330
rect 96846 24278 96898 24330
rect 127358 24278 127410 24330
rect 127462 24278 127514 24330
rect 127566 24278 127618 24330
rect 158078 24278 158130 24330
rect 158182 24278 158234 24330
rect 158286 24278 158338 24330
rect 188798 24278 188850 24330
rect 188902 24278 188954 24330
rect 189006 24278 189058 24330
rect 219518 24278 219570 24330
rect 219622 24278 219674 24330
rect 219726 24278 219778 24330
rect 250238 24278 250290 24330
rect 250342 24278 250394 24330
rect 250446 24278 250498 24330
rect 280958 24278 281010 24330
rect 281062 24278 281114 24330
rect 281166 24278 281218 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 81278 23494 81330 23546
rect 81382 23494 81434 23546
rect 81486 23494 81538 23546
rect 111998 23494 112050 23546
rect 112102 23494 112154 23546
rect 112206 23494 112258 23546
rect 142718 23494 142770 23546
rect 142822 23494 142874 23546
rect 142926 23494 142978 23546
rect 173438 23494 173490 23546
rect 173542 23494 173594 23546
rect 173646 23494 173698 23546
rect 204158 23494 204210 23546
rect 204262 23494 204314 23546
rect 204366 23494 204418 23546
rect 234878 23494 234930 23546
rect 234982 23494 235034 23546
rect 235086 23494 235138 23546
rect 265598 23494 265650 23546
rect 265702 23494 265754 23546
rect 265806 23494 265858 23546
rect 296318 23494 296370 23546
rect 296422 23494 296474 23546
rect 296526 23494 296578 23546
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 96638 22710 96690 22762
rect 96742 22710 96794 22762
rect 96846 22710 96898 22762
rect 127358 22710 127410 22762
rect 127462 22710 127514 22762
rect 127566 22710 127618 22762
rect 158078 22710 158130 22762
rect 158182 22710 158234 22762
rect 158286 22710 158338 22762
rect 188798 22710 188850 22762
rect 188902 22710 188954 22762
rect 189006 22710 189058 22762
rect 219518 22710 219570 22762
rect 219622 22710 219674 22762
rect 219726 22710 219778 22762
rect 250238 22710 250290 22762
rect 250342 22710 250394 22762
rect 250446 22710 250498 22762
rect 280958 22710 281010 22762
rect 281062 22710 281114 22762
rect 281166 22710 281218 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 81278 21926 81330 21978
rect 81382 21926 81434 21978
rect 81486 21926 81538 21978
rect 111998 21926 112050 21978
rect 112102 21926 112154 21978
rect 112206 21926 112258 21978
rect 142718 21926 142770 21978
rect 142822 21926 142874 21978
rect 142926 21926 142978 21978
rect 173438 21926 173490 21978
rect 173542 21926 173594 21978
rect 173646 21926 173698 21978
rect 204158 21926 204210 21978
rect 204262 21926 204314 21978
rect 204366 21926 204418 21978
rect 234878 21926 234930 21978
rect 234982 21926 235034 21978
rect 235086 21926 235138 21978
rect 265598 21926 265650 21978
rect 265702 21926 265754 21978
rect 265806 21926 265858 21978
rect 296318 21926 296370 21978
rect 296422 21926 296474 21978
rect 296526 21926 296578 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 96638 21142 96690 21194
rect 96742 21142 96794 21194
rect 96846 21142 96898 21194
rect 127358 21142 127410 21194
rect 127462 21142 127514 21194
rect 127566 21142 127618 21194
rect 158078 21142 158130 21194
rect 158182 21142 158234 21194
rect 158286 21142 158338 21194
rect 188798 21142 188850 21194
rect 188902 21142 188954 21194
rect 189006 21142 189058 21194
rect 219518 21142 219570 21194
rect 219622 21142 219674 21194
rect 219726 21142 219778 21194
rect 250238 21142 250290 21194
rect 250342 21142 250394 21194
rect 250446 21142 250498 21194
rect 280958 21142 281010 21194
rect 281062 21142 281114 21194
rect 281166 21142 281218 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 81278 20358 81330 20410
rect 81382 20358 81434 20410
rect 81486 20358 81538 20410
rect 111998 20358 112050 20410
rect 112102 20358 112154 20410
rect 112206 20358 112258 20410
rect 142718 20358 142770 20410
rect 142822 20358 142874 20410
rect 142926 20358 142978 20410
rect 173438 20358 173490 20410
rect 173542 20358 173594 20410
rect 173646 20358 173698 20410
rect 204158 20358 204210 20410
rect 204262 20358 204314 20410
rect 204366 20358 204418 20410
rect 234878 20358 234930 20410
rect 234982 20358 235034 20410
rect 235086 20358 235138 20410
rect 265598 20358 265650 20410
rect 265702 20358 265754 20410
rect 265806 20358 265858 20410
rect 296318 20358 296370 20410
rect 296422 20358 296474 20410
rect 296526 20358 296578 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 96638 19574 96690 19626
rect 96742 19574 96794 19626
rect 96846 19574 96898 19626
rect 127358 19574 127410 19626
rect 127462 19574 127514 19626
rect 127566 19574 127618 19626
rect 158078 19574 158130 19626
rect 158182 19574 158234 19626
rect 158286 19574 158338 19626
rect 188798 19574 188850 19626
rect 188902 19574 188954 19626
rect 189006 19574 189058 19626
rect 219518 19574 219570 19626
rect 219622 19574 219674 19626
rect 219726 19574 219778 19626
rect 250238 19574 250290 19626
rect 250342 19574 250394 19626
rect 250446 19574 250498 19626
rect 280958 19574 281010 19626
rect 281062 19574 281114 19626
rect 281166 19574 281218 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 81278 18790 81330 18842
rect 81382 18790 81434 18842
rect 81486 18790 81538 18842
rect 111998 18790 112050 18842
rect 112102 18790 112154 18842
rect 112206 18790 112258 18842
rect 142718 18790 142770 18842
rect 142822 18790 142874 18842
rect 142926 18790 142978 18842
rect 173438 18790 173490 18842
rect 173542 18790 173594 18842
rect 173646 18790 173698 18842
rect 204158 18790 204210 18842
rect 204262 18790 204314 18842
rect 204366 18790 204418 18842
rect 234878 18790 234930 18842
rect 234982 18790 235034 18842
rect 235086 18790 235138 18842
rect 265598 18790 265650 18842
rect 265702 18790 265754 18842
rect 265806 18790 265858 18842
rect 296318 18790 296370 18842
rect 296422 18790 296474 18842
rect 296526 18790 296578 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 96638 18006 96690 18058
rect 96742 18006 96794 18058
rect 96846 18006 96898 18058
rect 127358 18006 127410 18058
rect 127462 18006 127514 18058
rect 127566 18006 127618 18058
rect 158078 18006 158130 18058
rect 158182 18006 158234 18058
rect 158286 18006 158338 18058
rect 188798 18006 188850 18058
rect 188902 18006 188954 18058
rect 189006 18006 189058 18058
rect 219518 18006 219570 18058
rect 219622 18006 219674 18058
rect 219726 18006 219778 18058
rect 250238 18006 250290 18058
rect 250342 18006 250394 18058
rect 250446 18006 250498 18058
rect 280958 18006 281010 18058
rect 281062 18006 281114 18058
rect 281166 18006 281218 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 81278 17222 81330 17274
rect 81382 17222 81434 17274
rect 81486 17222 81538 17274
rect 111998 17222 112050 17274
rect 112102 17222 112154 17274
rect 112206 17222 112258 17274
rect 142718 17222 142770 17274
rect 142822 17222 142874 17274
rect 142926 17222 142978 17274
rect 173438 17222 173490 17274
rect 173542 17222 173594 17274
rect 173646 17222 173698 17274
rect 204158 17222 204210 17274
rect 204262 17222 204314 17274
rect 204366 17222 204418 17274
rect 234878 17222 234930 17274
rect 234982 17222 235034 17274
rect 235086 17222 235138 17274
rect 265598 17222 265650 17274
rect 265702 17222 265754 17274
rect 265806 17222 265858 17274
rect 296318 17222 296370 17274
rect 296422 17222 296474 17274
rect 296526 17222 296578 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 96638 16438 96690 16490
rect 96742 16438 96794 16490
rect 96846 16438 96898 16490
rect 127358 16438 127410 16490
rect 127462 16438 127514 16490
rect 127566 16438 127618 16490
rect 158078 16438 158130 16490
rect 158182 16438 158234 16490
rect 158286 16438 158338 16490
rect 188798 16438 188850 16490
rect 188902 16438 188954 16490
rect 189006 16438 189058 16490
rect 219518 16438 219570 16490
rect 219622 16438 219674 16490
rect 219726 16438 219778 16490
rect 250238 16438 250290 16490
rect 250342 16438 250394 16490
rect 250446 16438 250498 16490
rect 280958 16438 281010 16490
rect 281062 16438 281114 16490
rect 281166 16438 281218 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 81278 15654 81330 15706
rect 81382 15654 81434 15706
rect 81486 15654 81538 15706
rect 111998 15654 112050 15706
rect 112102 15654 112154 15706
rect 112206 15654 112258 15706
rect 142718 15654 142770 15706
rect 142822 15654 142874 15706
rect 142926 15654 142978 15706
rect 173438 15654 173490 15706
rect 173542 15654 173594 15706
rect 173646 15654 173698 15706
rect 204158 15654 204210 15706
rect 204262 15654 204314 15706
rect 204366 15654 204418 15706
rect 234878 15654 234930 15706
rect 234982 15654 235034 15706
rect 235086 15654 235138 15706
rect 265598 15654 265650 15706
rect 265702 15654 265754 15706
rect 265806 15654 265858 15706
rect 296318 15654 296370 15706
rect 296422 15654 296474 15706
rect 296526 15654 296578 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 96638 14870 96690 14922
rect 96742 14870 96794 14922
rect 96846 14870 96898 14922
rect 127358 14870 127410 14922
rect 127462 14870 127514 14922
rect 127566 14870 127618 14922
rect 158078 14870 158130 14922
rect 158182 14870 158234 14922
rect 158286 14870 158338 14922
rect 188798 14870 188850 14922
rect 188902 14870 188954 14922
rect 189006 14870 189058 14922
rect 219518 14870 219570 14922
rect 219622 14870 219674 14922
rect 219726 14870 219778 14922
rect 250238 14870 250290 14922
rect 250342 14870 250394 14922
rect 250446 14870 250498 14922
rect 280958 14870 281010 14922
rect 281062 14870 281114 14922
rect 281166 14870 281218 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 81278 14086 81330 14138
rect 81382 14086 81434 14138
rect 81486 14086 81538 14138
rect 111998 14086 112050 14138
rect 112102 14086 112154 14138
rect 112206 14086 112258 14138
rect 142718 14086 142770 14138
rect 142822 14086 142874 14138
rect 142926 14086 142978 14138
rect 173438 14086 173490 14138
rect 173542 14086 173594 14138
rect 173646 14086 173698 14138
rect 204158 14086 204210 14138
rect 204262 14086 204314 14138
rect 204366 14086 204418 14138
rect 234878 14086 234930 14138
rect 234982 14086 235034 14138
rect 235086 14086 235138 14138
rect 265598 14086 265650 14138
rect 265702 14086 265754 14138
rect 265806 14086 265858 14138
rect 296318 14086 296370 14138
rect 296422 14086 296474 14138
rect 296526 14086 296578 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 96638 13302 96690 13354
rect 96742 13302 96794 13354
rect 96846 13302 96898 13354
rect 127358 13302 127410 13354
rect 127462 13302 127514 13354
rect 127566 13302 127618 13354
rect 158078 13302 158130 13354
rect 158182 13302 158234 13354
rect 158286 13302 158338 13354
rect 188798 13302 188850 13354
rect 188902 13302 188954 13354
rect 189006 13302 189058 13354
rect 219518 13302 219570 13354
rect 219622 13302 219674 13354
rect 219726 13302 219778 13354
rect 250238 13302 250290 13354
rect 250342 13302 250394 13354
rect 250446 13302 250498 13354
rect 280958 13302 281010 13354
rect 281062 13302 281114 13354
rect 281166 13302 281218 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 81278 12518 81330 12570
rect 81382 12518 81434 12570
rect 81486 12518 81538 12570
rect 111998 12518 112050 12570
rect 112102 12518 112154 12570
rect 112206 12518 112258 12570
rect 142718 12518 142770 12570
rect 142822 12518 142874 12570
rect 142926 12518 142978 12570
rect 173438 12518 173490 12570
rect 173542 12518 173594 12570
rect 173646 12518 173698 12570
rect 204158 12518 204210 12570
rect 204262 12518 204314 12570
rect 204366 12518 204418 12570
rect 234878 12518 234930 12570
rect 234982 12518 235034 12570
rect 235086 12518 235138 12570
rect 265598 12518 265650 12570
rect 265702 12518 265754 12570
rect 265806 12518 265858 12570
rect 296318 12518 296370 12570
rect 296422 12518 296474 12570
rect 296526 12518 296578 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 96638 11734 96690 11786
rect 96742 11734 96794 11786
rect 96846 11734 96898 11786
rect 127358 11734 127410 11786
rect 127462 11734 127514 11786
rect 127566 11734 127618 11786
rect 158078 11734 158130 11786
rect 158182 11734 158234 11786
rect 158286 11734 158338 11786
rect 188798 11734 188850 11786
rect 188902 11734 188954 11786
rect 189006 11734 189058 11786
rect 219518 11734 219570 11786
rect 219622 11734 219674 11786
rect 219726 11734 219778 11786
rect 250238 11734 250290 11786
rect 250342 11734 250394 11786
rect 250446 11734 250498 11786
rect 280958 11734 281010 11786
rect 281062 11734 281114 11786
rect 281166 11734 281218 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 81278 10950 81330 11002
rect 81382 10950 81434 11002
rect 81486 10950 81538 11002
rect 111998 10950 112050 11002
rect 112102 10950 112154 11002
rect 112206 10950 112258 11002
rect 142718 10950 142770 11002
rect 142822 10950 142874 11002
rect 142926 10950 142978 11002
rect 173438 10950 173490 11002
rect 173542 10950 173594 11002
rect 173646 10950 173698 11002
rect 204158 10950 204210 11002
rect 204262 10950 204314 11002
rect 204366 10950 204418 11002
rect 234878 10950 234930 11002
rect 234982 10950 235034 11002
rect 235086 10950 235138 11002
rect 265598 10950 265650 11002
rect 265702 10950 265754 11002
rect 265806 10950 265858 11002
rect 296318 10950 296370 11002
rect 296422 10950 296474 11002
rect 296526 10950 296578 11002
rect 211934 10782 211986 10834
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 96638 10166 96690 10218
rect 96742 10166 96794 10218
rect 96846 10166 96898 10218
rect 127358 10166 127410 10218
rect 127462 10166 127514 10218
rect 127566 10166 127618 10218
rect 158078 10166 158130 10218
rect 158182 10166 158234 10218
rect 158286 10166 158338 10218
rect 188798 10166 188850 10218
rect 188902 10166 188954 10218
rect 189006 10166 189058 10218
rect 219518 10166 219570 10218
rect 219622 10166 219674 10218
rect 219726 10166 219778 10218
rect 250238 10166 250290 10218
rect 250342 10166 250394 10218
rect 250446 10166 250498 10218
rect 280958 10166 281010 10218
rect 281062 10166 281114 10218
rect 281166 10166 281218 10218
rect 199166 9886 199218 9938
rect 200062 9886 200114 9938
rect 217422 9886 217474 9938
rect 220894 9886 220946 9938
rect 211486 9774 211538 9826
rect 211710 9774 211762 9826
rect 212046 9774 212098 9826
rect 212494 9774 212546 9826
rect 211038 9662 211090 9714
rect 200958 9550 201010 9602
rect 210926 9550 210978 9602
rect 211262 9550 211314 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 81278 9382 81330 9434
rect 81382 9382 81434 9434
rect 81486 9382 81538 9434
rect 111998 9382 112050 9434
rect 112102 9382 112154 9434
rect 112206 9382 112258 9434
rect 142718 9382 142770 9434
rect 142822 9382 142874 9434
rect 142926 9382 142978 9434
rect 173438 9382 173490 9434
rect 173542 9382 173594 9434
rect 173646 9382 173698 9434
rect 204158 9382 204210 9434
rect 204262 9382 204314 9434
rect 204366 9382 204418 9434
rect 234878 9382 234930 9434
rect 234982 9382 235034 9434
rect 235086 9382 235138 9434
rect 265598 9382 265650 9434
rect 265702 9382 265754 9434
rect 265806 9382 265858 9434
rect 296318 9382 296370 9434
rect 296422 9382 296474 9434
rect 296526 9382 296578 9434
rect 188862 9214 188914 9266
rect 196030 9214 196082 9266
rect 198494 9214 198546 9266
rect 198830 9214 198882 9266
rect 201294 9214 201346 9266
rect 202302 9214 202354 9266
rect 203086 9214 203138 9266
rect 203646 9214 203698 9266
rect 216750 9214 216802 9266
rect 219102 9214 219154 9266
rect 219550 9214 219602 9266
rect 220446 9214 220498 9266
rect 222350 9214 222402 9266
rect 195582 9102 195634 9154
rect 199166 9102 199218 9154
rect 200398 9102 200450 9154
rect 208126 9102 208178 9154
rect 210142 9102 210194 9154
rect 211262 9102 211314 9154
rect 217198 9102 217250 9154
rect 217758 9102 217810 9154
rect 218430 9102 218482 9154
rect 219998 9102 220050 9154
rect 220670 9102 220722 9154
rect 221230 9102 221282 9154
rect 221902 9102 221954 9154
rect 192670 8990 192722 9042
rect 193006 8990 193058 9042
rect 193678 8990 193730 9042
rect 195358 8990 195410 9042
rect 199726 8990 199778 9042
rect 205774 8990 205826 9042
rect 207790 8990 207842 9042
rect 210814 8990 210866 9042
rect 212718 8990 212770 9042
rect 213390 8990 213442 9042
rect 213838 8990 213890 9042
rect 216526 8990 216578 9042
rect 216974 8990 217026 9042
rect 217982 8990 218034 9042
rect 218206 8990 218258 9042
rect 218766 8990 218818 9042
rect 220222 8990 220274 9042
rect 221454 8990 221506 9042
rect 221678 8990 221730 9042
rect 189422 8878 189474 8930
rect 199502 8878 199554 8930
rect 200958 8878 201010 8930
rect 201854 8878 201906 8930
rect 203198 8878 203250 8930
rect 206334 8878 206386 8930
rect 209246 8878 209298 8930
rect 210030 8878 210082 8930
rect 216414 8878 216466 8930
rect 200062 8766 200114 8818
rect 217870 8766 217922 8818
rect 220558 8766 220610 8818
rect 221790 8766 221842 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 96638 8598 96690 8650
rect 96742 8598 96794 8650
rect 96846 8598 96898 8650
rect 127358 8598 127410 8650
rect 127462 8598 127514 8650
rect 127566 8598 127618 8650
rect 158078 8598 158130 8650
rect 158182 8598 158234 8650
rect 158286 8598 158338 8650
rect 188798 8598 188850 8650
rect 188902 8598 188954 8650
rect 189006 8598 189058 8650
rect 219518 8598 219570 8650
rect 219622 8598 219674 8650
rect 219726 8598 219778 8650
rect 250238 8598 250290 8650
rect 250342 8598 250394 8650
rect 250446 8598 250498 8650
rect 280958 8598 281010 8650
rect 281062 8598 281114 8650
rect 281166 8598 281218 8650
rect 212270 8430 212322 8482
rect 221342 8430 221394 8482
rect 187630 8318 187682 8370
rect 189758 8318 189810 8370
rect 199054 8318 199106 8370
rect 199614 8318 199666 8370
rect 207678 8318 207730 8370
rect 222014 8318 222066 8370
rect 188638 8206 188690 8258
rect 189086 8206 189138 8258
rect 190766 8206 190818 8258
rect 199950 8206 200002 8258
rect 200846 8206 200898 8258
rect 203198 8206 203250 8258
rect 203422 8206 203474 8258
rect 204654 8206 204706 8258
rect 205102 8206 205154 8258
rect 205886 8206 205938 8258
rect 210702 8206 210754 8258
rect 211150 8206 211202 8258
rect 211710 8206 211762 8258
rect 212382 8206 212434 8258
rect 213390 8206 213442 8258
rect 217534 8206 217586 8258
rect 220782 8206 220834 8258
rect 221454 8206 221506 8258
rect 200062 8094 200114 8146
rect 202190 8094 202242 8146
rect 206894 8094 206946 8146
rect 210366 8094 210418 8146
rect 211374 8094 211426 8146
rect 212830 8094 212882 8146
rect 217758 8094 217810 8146
rect 221006 8094 221058 8146
rect 190430 7982 190482 8034
rect 201070 7982 201122 8034
rect 203086 7982 203138 8034
rect 205662 7982 205714 8034
rect 205998 7982 206050 8034
rect 209806 7982 209858 8034
rect 210590 7982 210642 8034
rect 210926 7982 210978 8034
rect 211934 7982 211986 8034
rect 212158 7982 212210 8034
rect 221230 7982 221282 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 81278 7814 81330 7866
rect 81382 7814 81434 7866
rect 81486 7814 81538 7866
rect 111998 7814 112050 7866
rect 112102 7814 112154 7866
rect 112206 7814 112258 7866
rect 142718 7814 142770 7866
rect 142822 7814 142874 7866
rect 142926 7814 142978 7866
rect 173438 7814 173490 7866
rect 173542 7814 173594 7866
rect 173646 7814 173698 7866
rect 204158 7814 204210 7866
rect 204262 7814 204314 7866
rect 204366 7814 204418 7866
rect 234878 7814 234930 7866
rect 234982 7814 235034 7866
rect 235086 7814 235138 7866
rect 265598 7814 265650 7866
rect 265702 7814 265754 7866
rect 265806 7814 265858 7866
rect 296318 7814 296370 7866
rect 296422 7814 296474 7866
rect 296526 7814 296578 7866
rect 196030 7646 196082 7698
rect 202862 7646 202914 7698
rect 204878 7646 204930 7698
rect 207342 7646 207394 7698
rect 215742 7646 215794 7698
rect 185390 7534 185442 7586
rect 186286 7534 186338 7586
rect 188078 7534 188130 7586
rect 188750 7534 188802 7586
rect 189310 7534 189362 7586
rect 191102 7534 191154 7586
rect 192670 7534 192722 7586
rect 195582 7534 195634 7586
rect 201070 7534 201122 7586
rect 202414 7534 202466 7586
rect 204654 7534 204706 7586
rect 209918 7534 209970 7586
rect 211598 7534 211650 7586
rect 185614 7422 185666 7474
rect 187854 7422 187906 7474
rect 189198 7422 189250 7474
rect 190654 7422 190706 7474
rect 192894 7422 192946 7474
rect 193790 7422 193842 7474
rect 195134 7422 195186 7474
rect 198494 7422 198546 7474
rect 200398 7422 200450 7474
rect 200846 7422 200898 7474
rect 202974 7422 203026 7474
rect 205774 7422 205826 7474
rect 210366 7422 210418 7474
rect 210926 7422 210978 7474
rect 214062 7422 214114 7474
rect 214510 7422 214562 7474
rect 216190 7422 216242 7474
rect 216414 7422 216466 7474
rect 216526 7422 216578 7474
rect 191662 7310 191714 7362
rect 199166 7310 199218 7362
rect 199614 7310 199666 7362
rect 203198 7310 203250 7362
rect 204878 7310 204930 7362
rect 205550 7310 205602 7362
rect 206334 7310 206386 7362
rect 206894 7310 206946 7362
rect 209470 7310 209522 7362
rect 216750 7310 216802 7362
rect 189870 7198 189922 7250
rect 197710 7198 197762 7250
rect 199838 7198 199890 7250
rect 200174 7198 200226 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 96638 7030 96690 7082
rect 96742 7030 96794 7082
rect 96846 7030 96898 7082
rect 127358 7030 127410 7082
rect 127462 7030 127514 7082
rect 127566 7030 127618 7082
rect 158078 7030 158130 7082
rect 158182 7030 158234 7082
rect 158286 7030 158338 7082
rect 188798 7030 188850 7082
rect 188902 7030 188954 7082
rect 189006 7030 189058 7082
rect 219518 7030 219570 7082
rect 219622 7030 219674 7082
rect 219726 7030 219778 7082
rect 250238 7030 250290 7082
rect 250342 7030 250394 7082
rect 250446 7030 250498 7082
rect 280958 7030 281010 7082
rect 281062 7030 281114 7082
rect 281166 7030 281218 7082
rect 199390 6750 199442 6802
rect 217758 6750 217810 6802
rect 184494 6638 184546 6690
rect 186734 6638 186786 6690
rect 187742 6638 187794 6690
rect 190318 6638 190370 6690
rect 190654 6638 190706 6690
rect 190990 6638 191042 6690
rect 192334 6638 192386 6690
rect 193230 6638 193282 6690
rect 193902 6638 193954 6690
rect 195918 6638 195970 6690
rect 196814 6638 196866 6690
rect 197598 6638 197650 6690
rect 197934 6638 197986 6690
rect 198606 6638 198658 6690
rect 201070 6638 201122 6690
rect 201630 6638 201682 6690
rect 203086 6638 203138 6690
rect 204654 6638 204706 6690
rect 206334 6638 206386 6690
rect 207454 6638 207506 6690
rect 213838 6638 213890 6690
rect 217198 6638 217250 6690
rect 218206 6638 218258 6690
rect 184382 6526 184434 6578
rect 188302 6526 188354 6578
rect 199614 6526 199666 6578
rect 204766 6526 204818 6578
rect 205102 6526 205154 6578
rect 184046 6414 184098 6466
rect 187406 6414 187458 6466
rect 192782 6414 192834 6466
rect 194350 6414 194402 6466
rect 204654 6414 204706 6466
rect 207006 6414 207058 6466
rect 207902 6414 207954 6466
rect 213614 6414 213666 6466
rect 217646 6414 217698 6466
rect 217870 6414 217922 6466
rect 218542 6414 218594 6466
rect 219102 6414 219154 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 81278 6246 81330 6298
rect 81382 6246 81434 6298
rect 81486 6246 81538 6298
rect 111998 6246 112050 6298
rect 112102 6246 112154 6298
rect 112206 6246 112258 6298
rect 142718 6246 142770 6298
rect 142822 6246 142874 6298
rect 142926 6246 142978 6298
rect 173438 6246 173490 6298
rect 173542 6246 173594 6298
rect 173646 6246 173698 6298
rect 204158 6246 204210 6298
rect 204262 6246 204314 6298
rect 204366 6246 204418 6298
rect 234878 6246 234930 6298
rect 234982 6246 235034 6298
rect 235086 6246 235138 6298
rect 265598 6246 265650 6298
rect 265702 6246 265754 6298
rect 265806 6246 265858 6298
rect 296318 6246 296370 6298
rect 296422 6246 296474 6298
rect 296526 6246 296578 6298
rect 185278 6078 185330 6130
rect 187518 6078 187570 6130
rect 193566 6078 193618 6130
rect 197710 6078 197762 6130
rect 203534 6078 203586 6130
rect 209470 6078 209522 6130
rect 214622 6078 214674 6130
rect 186398 5966 186450 6018
rect 187966 5966 188018 6018
rect 191662 5966 191714 6018
rect 191774 5966 191826 6018
rect 195582 5966 195634 6018
rect 199166 5966 199218 6018
rect 199502 5966 199554 6018
rect 205550 5966 205602 6018
rect 214958 5966 215010 6018
rect 216638 5966 216690 6018
rect 183710 5854 183762 5906
rect 184606 5854 184658 5906
rect 186174 5854 186226 5906
rect 186734 5854 186786 5906
rect 189310 5854 189362 5906
rect 191102 5854 191154 5906
rect 192894 5854 192946 5906
rect 193790 5854 193842 5906
rect 195358 5854 195410 5906
rect 196030 5854 196082 5906
rect 198046 5854 198098 5906
rect 200622 5854 200674 5906
rect 201294 5854 201346 5906
rect 201854 5854 201906 5906
rect 204542 5854 204594 5906
rect 205774 5854 205826 5906
rect 205998 5854 206050 5906
rect 206222 5854 206274 5906
rect 206558 5854 206610 5906
rect 210366 5854 210418 5906
rect 210814 5854 210866 5906
rect 211262 5854 211314 5906
rect 211374 5854 211426 5906
rect 216190 5854 216242 5906
rect 216414 5854 216466 5906
rect 188862 5742 188914 5794
rect 190430 5742 190482 5794
rect 203086 5742 203138 5794
rect 203982 5742 204034 5794
rect 204990 5742 205042 5794
rect 207006 5742 207058 5794
rect 207566 5742 207618 5794
rect 208014 5742 208066 5794
rect 208462 5742 208514 5794
rect 208910 5742 208962 5794
rect 209806 5742 209858 5794
rect 211598 5742 211650 5794
rect 215854 5742 215906 5794
rect 216526 5742 216578 5794
rect 217086 5742 217138 5794
rect 219550 5742 219602 5794
rect 223582 5742 223634 5794
rect 196814 5630 196866 5682
rect 206110 5630 206162 5682
rect 207454 5630 207506 5682
rect 208014 5630 208066 5682
rect 210590 5630 210642 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 96638 5462 96690 5514
rect 96742 5462 96794 5514
rect 96846 5462 96898 5514
rect 127358 5462 127410 5514
rect 127462 5462 127514 5514
rect 127566 5462 127618 5514
rect 158078 5462 158130 5514
rect 158182 5462 158234 5514
rect 158286 5462 158338 5514
rect 188798 5462 188850 5514
rect 188902 5462 188954 5514
rect 189006 5462 189058 5514
rect 219518 5462 219570 5514
rect 219622 5462 219674 5514
rect 219726 5462 219778 5514
rect 250238 5462 250290 5514
rect 250342 5462 250394 5514
rect 250446 5462 250498 5514
rect 280958 5462 281010 5514
rect 281062 5462 281114 5514
rect 281166 5462 281218 5514
rect 192782 5294 192834 5346
rect 204094 5294 204146 5346
rect 207342 5294 207394 5346
rect 210478 5294 210530 5346
rect 218318 5294 218370 5346
rect 220782 5294 220834 5346
rect 220894 5294 220946 5346
rect 93550 5182 93602 5234
rect 185950 5182 186002 5234
rect 192670 5182 192722 5234
rect 193230 5182 193282 5234
rect 195022 5182 195074 5234
rect 195470 5182 195522 5234
rect 206558 5182 206610 5234
rect 215294 5182 215346 5234
rect 217310 5182 217362 5234
rect 182702 5070 182754 5122
rect 183598 5070 183650 5122
rect 184718 5070 184770 5122
rect 185390 5070 185442 5122
rect 186398 5070 186450 5122
rect 187070 5070 187122 5122
rect 187518 5070 187570 5122
rect 190318 5070 190370 5122
rect 190654 5070 190706 5122
rect 190990 5070 191042 5122
rect 192334 5070 192386 5122
rect 194574 5070 194626 5122
rect 196254 5070 196306 5122
rect 199054 5070 199106 5122
rect 199726 5070 199778 5122
rect 201070 5070 201122 5122
rect 201742 5070 201794 5122
rect 202526 5070 202578 5122
rect 202974 5070 203026 5122
rect 204094 5070 204146 5122
rect 204542 5070 204594 5122
rect 205102 5070 205154 5122
rect 205774 5070 205826 5122
rect 206446 5070 206498 5122
rect 206782 5070 206834 5122
rect 207454 5070 207506 5122
rect 208014 5070 208066 5122
rect 208798 5070 208850 5122
rect 209470 5070 209522 5122
rect 210254 5070 210306 5122
rect 210702 5070 210754 5122
rect 212270 5070 212322 5122
rect 214286 5070 214338 5122
rect 214734 5070 214786 5122
rect 215182 5070 215234 5122
rect 215630 5070 215682 5122
rect 216190 5070 216242 5122
rect 216862 5070 216914 5122
rect 217982 5070 218034 5122
rect 218542 5070 218594 5122
rect 218990 5070 219042 5122
rect 219774 5070 219826 5122
rect 220558 5070 220610 5122
rect 221118 5070 221170 5122
rect 221566 5070 221618 5122
rect 221790 5070 221842 5122
rect 222574 5070 222626 5122
rect 223470 5070 223522 5122
rect 224030 5070 224082 5122
rect 186622 4958 186674 5010
rect 188862 4958 188914 5010
rect 197598 4958 197650 5010
rect 197934 4958 197986 5010
rect 201966 4958 202018 5010
rect 203534 4958 203586 5010
rect 203982 4958 204034 5010
rect 205998 4958 206050 5010
rect 207230 4958 207282 5010
rect 208350 4958 208402 5010
rect 209582 4958 209634 5010
rect 209918 4958 209970 5010
rect 212382 4958 212434 5010
rect 212606 4958 212658 5010
rect 212830 4958 212882 5010
rect 216078 4958 216130 5010
rect 217422 4958 217474 5010
rect 217758 4958 217810 5010
rect 218878 4958 218930 5010
rect 219998 4958 220050 5010
rect 220222 4958 220274 5010
rect 221678 4958 221730 5010
rect 183374 4846 183426 4898
rect 187406 4846 187458 4898
rect 193118 4846 193170 4898
rect 193790 4846 193842 4898
rect 196142 4846 196194 4898
rect 203086 4846 203138 4898
rect 203758 4846 203810 4898
rect 206222 4846 206274 4898
rect 207006 4846 207058 4898
rect 211038 4846 211090 4898
rect 211822 4846 211874 4898
rect 214510 4846 214562 4898
rect 215406 4846 215458 4898
rect 216302 4846 216354 4898
rect 219102 4846 219154 4898
rect 223022 4846 223074 4898
rect 223134 4846 223186 4898
rect 223246 4846 223298 4898
rect 223918 4846 223970 4898
rect 224142 4846 224194 4898
rect 224702 4846 224754 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 81278 4678 81330 4730
rect 81382 4678 81434 4730
rect 81486 4678 81538 4730
rect 111998 4678 112050 4730
rect 112102 4678 112154 4730
rect 112206 4678 112258 4730
rect 142718 4678 142770 4730
rect 142822 4678 142874 4730
rect 142926 4678 142978 4730
rect 173438 4678 173490 4730
rect 173542 4678 173594 4730
rect 173646 4678 173698 4730
rect 204158 4678 204210 4730
rect 204262 4678 204314 4730
rect 204366 4678 204418 4730
rect 234878 4678 234930 4730
rect 234982 4678 235034 4730
rect 235086 4678 235138 4730
rect 265598 4678 265650 4730
rect 265702 4678 265754 4730
rect 265806 4678 265858 4730
rect 296318 4678 296370 4730
rect 296422 4678 296474 4730
rect 296526 4678 296578 4730
rect 12462 4510 12514 4562
rect 54350 4510 54402 4562
rect 71150 4510 71202 4562
rect 74846 4510 74898 4562
rect 96238 4510 96290 4562
rect 122558 4510 122610 4562
rect 182366 4510 182418 4562
rect 184718 4510 184770 4562
rect 189310 4510 189362 4562
rect 189870 4510 189922 4562
rect 195358 4510 195410 4562
rect 196366 4510 196418 4562
rect 197150 4510 197202 4562
rect 197710 4510 197762 4562
rect 204878 4510 204930 4562
rect 212494 4510 212546 4562
rect 212606 4510 212658 4562
rect 215294 4510 215346 4562
rect 215406 4510 215458 4562
rect 215966 4510 216018 4562
rect 217086 4510 217138 4562
rect 217310 4510 217362 4562
rect 220110 4510 220162 4562
rect 11566 4398 11618 4450
rect 11902 4398 11954 4450
rect 71374 4398 71426 4450
rect 71710 4398 71762 4450
rect 75070 4398 75122 4450
rect 75406 4398 75458 4450
rect 83134 4398 83186 4450
rect 83470 4398 83522 4450
rect 86718 4398 86770 4450
rect 87054 4398 87106 4450
rect 93886 4398 93938 4450
rect 94222 4398 94274 4450
rect 96462 4398 96514 4450
rect 96798 4398 96850 4450
rect 187966 4398 188018 4450
rect 190542 4398 190594 4450
rect 191662 4398 191714 4450
rect 199166 4398 199218 4450
rect 199502 4398 199554 4450
rect 202974 4398 203026 4450
rect 207006 4398 207058 4450
rect 208238 4398 208290 4450
rect 210814 4398 210866 4450
rect 216750 4398 216802 4450
rect 217534 4398 217586 4450
rect 220670 4398 220722 4450
rect 221790 4398 221842 4450
rect 76638 4286 76690 4338
rect 80222 4286 80274 4338
rect 83806 4286 83858 4338
rect 87950 4286 88002 4338
rect 90974 4286 91026 4338
rect 182814 4286 182866 4338
rect 183710 4286 183762 4338
rect 184606 4286 184658 4338
rect 186174 4286 186226 4338
rect 186398 4286 186450 4338
rect 186734 4286 186786 4338
rect 189870 4286 189922 4338
rect 192782 4286 192834 4338
rect 193454 4286 193506 4338
rect 193678 4286 193730 4338
rect 197710 4286 197762 4338
rect 200622 4286 200674 4338
rect 201294 4286 201346 4338
rect 201854 4286 201906 4338
rect 203198 4286 203250 4338
rect 203758 4286 203810 4338
rect 204206 4286 204258 4338
rect 205550 4286 205602 4338
rect 208798 4286 208850 4338
rect 210030 4286 210082 4338
rect 210254 4286 210306 4338
rect 211934 4286 211986 4338
rect 212270 4286 212322 4338
rect 214846 4286 214898 4338
rect 215518 4286 215570 4338
rect 216526 4286 216578 4338
rect 217982 4286 218034 4338
rect 219550 4286 219602 4338
rect 219886 4286 219938 4338
rect 221342 4286 221394 4338
rect 221902 4286 221954 4338
rect 222014 4286 222066 4338
rect 222574 4286 222626 4338
rect 223022 4286 223074 4338
rect 223246 4286 223298 4338
rect 223694 4286 223746 4338
rect 50766 4174 50818 4226
rect 89070 4174 89122 4226
rect 111806 4174 111858 4226
rect 115390 4174 115442 4226
rect 181582 4174 181634 4226
rect 182254 4174 182306 4226
rect 182702 4174 182754 4226
rect 195806 4174 195858 4226
rect 206894 4174 206946 4226
rect 210366 4174 210418 4226
rect 217422 4174 217474 4226
rect 219326 4174 219378 4226
rect 219998 4174 220050 4226
rect 223134 4174 223186 4226
rect 77646 4062 77698 4114
rect 81230 4062 81282 4114
rect 84814 4062 84866 4114
rect 91982 4062 92034 4114
rect 186846 4062 186898 4114
rect 204542 4062 204594 4114
rect 221118 4062 221170 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 96638 3894 96690 3946
rect 96742 3894 96794 3946
rect 96846 3894 96898 3946
rect 127358 3894 127410 3946
rect 127462 3894 127514 3946
rect 127566 3894 127618 3946
rect 158078 3894 158130 3946
rect 158182 3894 158234 3946
rect 158286 3894 158338 3946
rect 188798 3894 188850 3946
rect 188902 3894 188954 3946
rect 189006 3894 189058 3946
rect 219518 3894 219570 3946
rect 219622 3894 219674 3946
rect 219726 3894 219778 3946
rect 250238 3894 250290 3946
rect 250342 3894 250394 3946
rect 250446 3894 250498 3946
rect 280958 3894 281010 3946
rect 281062 3894 281114 3946
rect 281166 3894 281218 3946
rect 182366 3726 182418 3778
rect 208238 3726 208290 3778
rect 208686 3726 208738 3778
rect 215406 3726 215458 3778
rect 216190 3726 216242 3778
rect 220782 3726 220834 3778
rect 221566 3726 221618 3778
rect 40686 3614 40738 3666
rect 43822 3614 43874 3666
rect 44494 3614 44546 3666
rect 47630 3614 47682 3666
rect 48190 3614 48242 3666
rect 51774 3614 51826 3666
rect 55358 3614 55410 3666
rect 58270 3614 58322 3666
rect 59054 3614 59106 3666
rect 61966 3614 62018 3666
rect 62862 3614 62914 3666
rect 65774 3614 65826 3666
rect 66670 3614 66722 3666
rect 69582 3614 69634 3666
rect 70478 3614 70530 3666
rect 73390 3614 73442 3666
rect 78318 3614 78370 3666
rect 82910 3614 82962 3666
rect 86494 3614 86546 3666
rect 88734 3614 88786 3666
rect 101614 3614 101666 3666
rect 105422 3614 105474 3666
rect 109118 3614 109170 3666
rect 112702 3614 112754 3666
rect 116286 3614 116338 3666
rect 119198 3614 119250 3666
rect 119982 3614 120034 3666
rect 182030 3614 182082 3666
rect 182254 3614 182306 3666
rect 196814 3614 196866 3666
rect 198158 3614 198210 3666
rect 204542 3614 204594 3666
rect 205662 3614 205714 3666
rect 206670 3614 206722 3666
rect 208686 3614 208738 3666
rect 209134 3614 209186 3666
rect 211374 3614 211426 3666
rect 215406 3614 215458 3666
rect 222014 3614 222066 3666
rect 267038 3614 267090 3666
rect 270622 3614 270674 3666
rect 281374 3614 281426 3666
rect 288542 3614 288594 3666
rect 292126 3614 292178 3666
rect 11566 3502 11618 3554
rect 43038 3502 43090 3554
rect 46846 3502 46898 3554
rect 50542 3502 50594 3554
rect 54126 3502 54178 3554
rect 57262 3502 57314 3554
rect 60958 3502 61010 3554
rect 65214 3502 65266 3554
rect 68910 3502 68962 3554
rect 72830 3502 72882 3554
rect 74062 3502 74114 3554
rect 78654 3502 78706 3554
rect 89406 3502 89458 3554
rect 94222 3502 94274 3554
rect 97582 3502 97634 3554
rect 103966 3502 104018 3554
rect 107774 3502 107826 3554
rect 111470 3502 111522 3554
rect 115054 3502 115106 3554
rect 118638 3502 118690 3554
rect 122334 3502 122386 3554
rect 182814 3502 182866 3554
rect 183710 3502 183762 3554
rect 185950 3502 186002 3554
rect 188526 3502 188578 3554
rect 193118 3502 193170 3554
rect 193566 3502 193618 3554
rect 194798 3502 194850 3554
rect 195358 3502 195410 3554
rect 201630 3502 201682 3554
rect 202414 3502 202466 3554
rect 202750 3502 202802 3554
rect 203534 3502 203586 3554
rect 203982 3502 204034 3554
rect 205102 3502 205154 3554
rect 205326 3502 205378 3554
rect 205550 3502 205602 3554
rect 206110 3502 206162 3554
rect 207566 3502 207618 3554
rect 208238 3502 208290 3554
rect 209470 3502 209522 3554
rect 210030 3502 210082 3554
rect 210590 3502 210642 3554
rect 211598 3502 211650 3554
rect 212046 3502 212098 3554
rect 213054 3502 213106 3554
rect 216638 3502 216690 3554
rect 220222 3502 220274 3554
rect 220894 3502 220946 3554
rect 223806 3502 223858 3554
rect 227390 3502 227442 3554
rect 230974 3502 231026 3554
rect 234558 3502 234610 3554
rect 238142 3502 238194 3554
rect 241838 3502 241890 3554
rect 245646 3502 245698 3554
rect 249454 3502 249506 3554
rect 253262 3502 253314 3554
rect 256062 3502 256114 3554
rect 259646 3502 259698 3554
rect 263230 3502 263282 3554
rect 285070 3502 285122 3554
rect 10110 3390 10162 3442
rect 75630 3390 75682 3442
rect 78990 3390 79042 3442
rect 89630 3390 89682 3442
rect 104750 3390 104802 3442
rect 108558 3390 108610 3442
rect 123118 3390 123170 3442
rect 123566 3390 123618 3442
rect 123902 3390 123954 3442
rect 126926 3390 126978 3442
rect 127374 3390 127426 3442
rect 127710 3390 127762 3442
rect 130734 3390 130786 3442
rect 131182 3390 131234 3442
rect 131518 3390 131570 3442
rect 133758 3390 133810 3442
rect 133982 3390 134034 3442
rect 134318 3390 134370 3442
rect 137342 3390 137394 3442
rect 137566 3390 137618 3442
rect 137902 3390 137954 3442
rect 140926 3390 140978 3442
rect 141150 3390 141202 3442
rect 141486 3390 141538 3442
rect 144510 3390 144562 3442
rect 144734 3390 144786 3442
rect 145070 3390 145122 3442
rect 148094 3390 148146 3442
rect 148318 3390 148370 3442
rect 148654 3390 148706 3442
rect 151678 3390 151730 3442
rect 151902 3390 151954 3442
rect 152238 3390 152290 3442
rect 155262 3390 155314 3442
rect 155486 3390 155538 3442
rect 155822 3390 155874 3442
rect 158846 3390 158898 3442
rect 159070 3390 159122 3442
rect 159406 3390 159458 3442
rect 162430 3390 162482 3442
rect 162654 3390 162706 3442
rect 166014 3390 166066 3442
rect 166238 3390 166290 3442
rect 166574 3390 166626 3442
rect 169598 3390 169650 3442
rect 169822 3390 169874 3442
rect 170158 3390 170210 3442
rect 172622 3390 172674 3442
rect 173406 3390 173458 3442
rect 173742 3390 173794 3442
rect 176430 3390 176482 3442
rect 176990 3390 177042 3442
rect 180238 3390 180290 3442
rect 180686 3390 180738 3442
rect 181022 3390 181074 3442
rect 183374 3390 183426 3442
rect 183934 3390 183986 3442
rect 184718 3390 184770 3442
rect 187854 3390 187906 3442
rect 188302 3390 188354 3442
rect 190094 3390 190146 3442
rect 190542 3390 190594 3442
rect 190766 3390 190818 3442
rect 190878 3390 190930 3442
rect 191214 3390 191266 3442
rect 191550 3390 191602 3442
rect 195918 3390 195970 3442
rect 196254 3390 196306 3442
rect 197150 3390 197202 3442
rect 197598 3390 197650 3442
rect 198494 3390 198546 3442
rect 198830 3390 198882 3442
rect 199838 3390 199890 3442
rect 200398 3390 200450 3442
rect 200846 3390 200898 3442
rect 201294 3390 201346 3442
rect 201742 3390 201794 3442
rect 203086 3390 203138 3442
rect 204878 3390 204930 3442
rect 205886 3390 205938 3442
rect 207342 3390 207394 3442
rect 209022 3390 209074 3442
rect 209246 3390 209298 3442
rect 209806 3390 209858 3442
rect 211150 3390 211202 3442
rect 211374 3390 211426 3442
rect 212606 3390 212658 3442
rect 212830 3390 212882 3442
rect 219326 3390 219378 3442
rect 219550 3390 219602 3442
rect 219886 3390 219938 3442
rect 220446 3390 220498 3442
rect 220670 3390 220722 3442
rect 221230 3390 221282 3442
rect 221454 3390 221506 3442
rect 223358 3390 223410 3442
rect 226942 3390 226994 3442
rect 230526 3390 230578 3442
rect 233550 3390 233602 3442
rect 237358 3390 237410 3442
rect 241166 3390 241218 3442
rect 244974 3390 245026 3442
rect 245422 3390 245474 3442
rect 248782 3390 248834 3442
rect 249230 3390 249282 3442
rect 252590 3390 252642 3442
rect 255614 3390 255666 3442
rect 259198 3390 259250 3442
rect 262782 3390 262834 3442
rect 266366 3390 266418 3442
rect 266590 3390 266642 3442
rect 269950 3390 270002 3442
rect 270174 3390 270226 3442
rect 273534 3390 273586 3442
rect 273758 3390 273810 3442
rect 274318 3390 274370 3442
rect 277118 3390 277170 3442
rect 277342 3390 277394 3442
rect 277902 3390 277954 3442
rect 280702 3390 280754 3442
rect 280926 3390 280978 3442
rect 284286 3390 284338 3442
rect 284510 3390 284562 3442
rect 287870 3390 287922 3442
rect 288094 3390 288146 3442
rect 291454 3390 291506 3442
rect 291678 3390 291730 3442
rect 12238 3278 12290 3330
rect 15710 3278 15762 3330
rect 19294 3278 19346 3330
rect 22878 3278 22930 3330
rect 26462 3278 26514 3330
rect 30046 3278 30098 3330
rect 33630 3278 33682 3330
rect 37214 3278 37266 3330
rect 94782 3278 94834 3330
rect 98590 3278 98642 3330
rect 162990 3278 163042 3330
rect 177326 3278 177378 3330
rect 184830 3278 184882 3330
rect 186734 3278 186786 3330
rect 193342 3278 193394 3330
rect 215854 3278 215906 3330
rect 216414 3278 216466 3330
rect 223582 3278 223634 3330
rect 227166 3278 227218 3330
rect 230750 3278 230802 3330
rect 234334 3278 234386 3330
rect 237918 3278 237970 3330
rect 241614 3278 241666 3330
rect 253038 3278 253090 3330
rect 255838 3278 255890 3330
rect 259422 3278 259474 3330
rect 263006 3278 263058 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 81278 3110 81330 3162
rect 81382 3110 81434 3162
rect 81486 3110 81538 3162
rect 111998 3110 112050 3162
rect 112102 3110 112154 3162
rect 112206 3110 112258 3162
rect 142718 3110 142770 3162
rect 142822 3110 142874 3162
rect 142926 3110 142978 3162
rect 173438 3110 173490 3162
rect 173542 3110 173594 3162
rect 173646 3110 173698 3162
rect 204158 3110 204210 3162
rect 204262 3110 204314 3162
rect 204366 3110 204418 3162
rect 234878 3110 234930 3162
rect 234982 3110 235034 3162
rect 235086 3110 235138 3162
rect 265598 3110 265650 3162
rect 265702 3110 265754 3162
rect 265806 3110 265858 3162
rect 296318 3110 296370 3162
rect 296422 3110 296474 3162
rect 296526 3110 296578 3162
<< metal2 >>
rect 7392 59200 7504 60000
rect 12768 59200 12880 60000
rect 18144 59200 18256 60000
rect 23520 59200 23632 60000
rect 28896 59200 29008 60000
rect 34272 59200 34384 60000
rect 39648 59200 39760 60000
rect 45024 59200 45136 60000
rect 50400 59200 50512 60000
rect 55776 59200 55888 60000
rect 61152 59200 61264 60000
rect 66528 59200 66640 60000
rect 71904 59200 72016 60000
rect 77280 59200 77392 60000
rect 82656 59200 82768 60000
rect 88032 59200 88144 60000
rect 93408 59200 93520 60000
rect 98784 59200 98896 60000
rect 104160 59200 104272 60000
rect 109536 59200 109648 60000
rect 114912 59200 115024 60000
rect 120288 59200 120400 60000
rect 125664 59200 125776 60000
rect 131040 59200 131152 60000
rect 136416 59200 136528 60000
rect 141792 59200 141904 60000
rect 147168 59200 147280 60000
rect 152544 59200 152656 60000
rect 157920 59200 158032 60000
rect 163296 59200 163408 60000
rect 168672 59200 168784 60000
rect 174048 59200 174160 60000
rect 179424 59200 179536 60000
rect 184800 59200 184912 60000
rect 190176 59200 190288 60000
rect 195552 59200 195664 60000
rect 200928 59200 201040 60000
rect 206304 59200 206416 60000
rect 211680 59200 211792 60000
rect 217056 59200 217168 60000
rect 222432 59200 222544 60000
rect 227808 59200 227920 60000
rect 233184 59200 233296 60000
rect 238560 59200 238672 60000
rect 243936 59200 244048 60000
rect 249312 59200 249424 60000
rect 254688 59200 254800 60000
rect 260064 59200 260176 60000
rect 265440 59200 265552 60000
rect 270816 59200 270928 60000
rect 276192 59200 276304 60000
rect 281568 59200 281680 60000
rect 286944 59200 287056 60000
rect 292320 59200 292432 60000
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 7420 52052 7476 59200
rect 7420 51986 7476 51996
rect 11900 56642 11956 56654
rect 11900 56590 11902 56642
rect 11954 56590 11956 56642
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 11900 4564 11956 56590
rect 12684 56308 12740 56318
rect 12796 56308 12852 59200
rect 13132 56642 13188 56654
rect 13132 56590 13134 56642
rect 13186 56590 13188 56642
rect 12684 56306 13076 56308
rect 12684 56254 12686 56306
rect 12738 56254 13076 56306
rect 12684 56252 13076 56254
rect 12684 56242 12740 56252
rect 13020 55972 13076 56252
rect 13132 56194 13188 56590
rect 18172 56308 18228 59200
rect 23548 56642 23604 59200
rect 23548 56590 23550 56642
rect 23602 56590 23604 56642
rect 23548 56578 23604 56590
rect 24108 56642 24164 56654
rect 24108 56590 24110 56642
rect 24162 56590 24164 56642
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 18396 56308 18452 56318
rect 18172 56306 18452 56308
rect 18172 56254 18174 56306
rect 18226 56254 18398 56306
rect 18450 56254 18452 56306
rect 18172 56252 18452 56254
rect 18172 56242 18228 56252
rect 18396 56242 18452 56252
rect 19180 56308 19236 56318
rect 19180 56214 19236 56252
rect 24108 56306 24164 56590
rect 24108 56254 24110 56306
rect 24162 56254 24164 56306
rect 24108 56242 24164 56254
rect 24556 56642 24612 56654
rect 24556 56590 24558 56642
rect 24610 56590 24612 56642
rect 24556 56306 24612 56590
rect 24556 56254 24558 56306
rect 24610 56254 24612 56306
rect 24556 56242 24612 56254
rect 28924 56308 28980 59200
rect 29148 56308 29204 56318
rect 28924 56306 29204 56308
rect 28924 56254 28926 56306
rect 28978 56254 29150 56306
rect 29202 56254 29204 56306
rect 28924 56252 29204 56254
rect 28924 56242 28980 56252
rect 29148 56242 29204 56252
rect 34300 56308 34356 59200
rect 34524 56308 34580 56318
rect 34300 56306 34580 56308
rect 34300 56254 34302 56306
rect 34354 56254 34526 56306
rect 34578 56254 34580 56306
rect 34300 56252 34580 56254
rect 34300 56242 34356 56252
rect 34524 56242 34580 56252
rect 39340 56308 39396 56318
rect 39676 56308 39732 59200
rect 39900 56308 39956 56318
rect 39340 56306 39956 56308
rect 39340 56254 39342 56306
rect 39394 56254 39902 56306
rect 39954 56254 39956 56306
rect 39340 56252 39956 56254
rect 39340 56242 39396 56252
rect 39900 56242 39956 56252
rect 45052 56308 45108 59200
rect 45276 56308 45332 56318
rect 45052 56306 45332 56308
rect 45052 56254 45054 56306
rect 45106 56254 45278 56306
rect 45330 56254 45332 56306
rect 45052 56252 45332 56254
rect 50428 56308 50484 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 50764 56308 50820 56318
rect 51212 56308 51268 56318
rect 50428 56306 51268 56308
rect 50428 56254 50766 56306
rect 50818 56254 51214 56306
rect 51266 56254 51268 56306
rect 50428 56252 51268 56254
rect 45052 56242 45108 56252
rect 45276 56242 45332 56252
rect 50764 56242 50820 56252
rect 51212 56242 51268 56252
rect 55804 56308 55860 59200
rect 56028 56308 56084 56318
rect 55804 56306 56084 56308
rect 55804 56254 55806 56306
rect 55858 56254 56030 56306
rect 56082 56254 56084 56306
rect 55804 56252 56084 56254
rect 55804 56242 55860 56252
rect 56028 56242 56084 56252
rect 61180 56308 61236 59200
rect 66556 57540 66612 59200
rect 66556 57484 67060 57540
rect 61404 56308 61460 56318
rect 61180 56306 61460 56308
rect 61180 56254 61182 56306
rect 61234 56254 61406 56306
rect 61458 56254 61460 56306
rect 61180 56252 61460 56254
rect 61180 56242 61236 56252
rect 61404 56242 61460 56252
rect 13132 56142 13134 56194
rect 13186 56142 13188 56194
rect 13132 56130 13188 56142
rect 13356 56082 13412 56094
rect 13356 56030 13358 56082
rect 13410 56030 13412 56082
rect 13356 55972 13412 56030
rect 13020 55916 13412 55972
rect 25116 55970 25172 55982
rect 25116 55918 25118 55970
rect 25170 55918 25172 55970
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 25116 7588 25172 55918
rect 29708 55970 29764 55982
rect 29708 55918 29710 55970
rect 29762 55918 29764 55970
rect 29708 9268 29764 55918
rect 35084 55970 35140 55982
rect 35084 55918 35086 55970
rect 35138 55918 35140 55970
rect 35084 19348 35140 55918
rect 40460 55970 40516 55982
rect 40460 55918 40462 55970
rect 40514 55918 40516 55970
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35084 19282 35140 19292
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 40460 15988 40516 55918
rect 45836 55970 45892 55982
rect 45836 55918 45838 55970
rect 45890 55918 45892 55970
rect 40460 15922 40516 15932
rect 43820 24500 43876 24510
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 29708 9202 29764 9212
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 25116 7522 25172 7532
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 12460 4564 12516 4574
rect 11900 4562 12516 4564
rect 11900 4510 12462 4562
rect 12514 4510 12516 4562
rect 11900 4508 12516 4510
rect 11564 4450 11620 4462
rect 11564 4398 11566 4450
rect 11618 4398 11620 4450
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 11564 3554 11620 4398
rect 11900 4450 11956 4508
rect 12460 4498 12516 4508
rect 11900 4398 11902 4450
rect 11954 4398 11956 4450
rect 11900 4386 11956 4398
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 40684 3668 40740 3678
rect 11564 3502 11566 3554
rect 11618 3502 11620 3554
rect 11564 3490 11620 3502
rect 40572 3666 40740 3668
rect 40572 3614 40686 3666
rect 40738 3614 40740 3666
rect 40572 3612 40740 3614
rect 8316 3444 8372 3454
rect 8316 800 8372 3388
rect 10108 3444 10164 3454
rect 10108 3350 10164 3388
rect 12236 3332 12292 3342
rect 15708 3332 15764 3342
rect 19292 3332 19348 3342
rect 22876 3332 22932 3342
rect 26460 3332 26516 3342
rect 30044 3332 30100 3342
rect 33628 3332 33684 3342
rect 37212 3332 37268 3342
rect 11900 3330 12292 3332
rect 11900 3278 12238 3330
rect 12290 3278 12292 3330
rect 11900 3276 12292 3278
rect 11900 800 11956 3276
rect 12236 3266 12292 3276
rect 15484 3330 15764 3332
rect 15484 3278 15710 3330
rect 15762 3278 15764 3330
rect 15484 3276 15764 3278
rect 15484 800 15540 3276
rect 15708 3266 15764 3276
rect 19068 3330 19348 3332
rect 19068 3278 19294 3330
rect 19346 3278 19348 3330
rect 19068 3276 19348 3278
rect 19068 800 19124 3276
rect 19292 3266 19348 3276
rect 22652 3330 22932 3332
rect 22652 3278 22878 3330
rect 22930 3278 22932 3330
rect 22652 3276 22932 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 22652 800 22708 3276
rect 22876 3266 22932 3276
rect 26236 3330 26516 3332
rect 26236 3278 26462 3330
rect 26514 3278 26516 3330
rect 26236 3276 26516 3278
rect 26236 800 26292 3276
rect 26460 3266 26516 3276
rect 29820 3330 30100 3332
rect 29820 3278 30046 3330
rect 30098 3278 30100 3330
rect 29820 3276 30100 3278
rect 29820 800 29876 3276
rect 30044 3266 30100 3276
rect 33404 3330 33684 3332
rect 33404 3278 33630 3330
rect 33682 3278 33684 3330
rect 33404 3276 33684 3278
rect 33404 800 33460 3276
rect 33628 3266 33684 3276
rect 36988 3330 37268 3332
rect 36988 3278 37214 3330
rect 37266 3278 37268 3330
rect 36988 3276 37268 3278
rect 36988 800 37044 3276
rect 37212 3266 37268 3276
rect 40572 800 40628 3612
rect 40684 3602 40740 3612
rect 43036 3668 43092 3678
rect 43036 3554 43092 3612
rect 43820 3668 43876 24444
rect 45836 21028 45892 55918
rect 51772 55972 51828 55982
rect 51772 55878 51828 55916
rect 52892 55972 52948 55982
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 45836 20962 45892 20972
rect 47628 26068 47684 26078
rect 44492 3668 44548 3678
rect 43820 3574 43876 3612
rect 44156 3666 44548 3668
rect 44156 3614 44494 3666
rect 44546 3614 44548 3666
rect 44156 3612 44548 3614
rect 43036 3502 43038 3554
rect 43090 3502 43092 3554
rect 43036 3490 43092 3502
rect 44156 800 44212 3612
rect 44492 3602 44548 3612
rect 46844 3668 46900 3678
rect 46844 3554 46900 3612
rect 47628 3668 47684 26012
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 52892 22932 52948 55916
rect 56588 55970 56644 55982
rect 56588 55918 56590 55970
rect 56642 55918 56644 55970
rect 52892 22866 52948 22876
rect 54348 41188 54404 41198
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 54348 4564 54404 41132
rect 56588 5908 56644 55918
rect 61964 55970 62020 55982
rect 61964 55918 61966 55970
rect 62018 55918 62020 55970
rect 61964 55524 62020 55918
rect 67004 55970 67060 57484
rect 67004 55918 67006 55970
rect 67058 55918 67060 55970
rect 67004 55906 67060 55918
rect 69356 56082 69412 56094
rect 69356 56030 69358 56082
rect 69410 56030 69412 56082
rect 69356 55972 69412 56030
rect 69356 55906 69412 55916
rect 70476 55972 70532 55982
rect 70476 55878 70532 55916
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 61964 55458 62020 55468
rect 71932 55468 71988 59200
rect 77308 57090 77364 59200
rect 77308 57038 77310 57090
rect 77362 57038 77364 57090
rect 77308 57026 77364 57038
rect 78092 57090 78148 57102
rect 78092 57038 78094 57090
rect 78146 57038 78148 57090
rect 73052 55972 73108 55982
rect 71932 55412 72436 55468
rect 72380 55410 72436 55412
rect 72380 55358 72382 55410
rect 72434 55358 72436 55410
rect 72380 55346 72436 55358
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 68236 36260 68292 36270
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 60956 32788 61012 32798
rect 56588 5842 56644 5852
rect 57260 31108 57316 31118
rect 54124 4562 54404 4564
rect 54124 4510 54350 4562
rect 54402 4510 54404 4562
rect 54124 4508 54404 4510
rect 50764 4226 50820 4238
rect 50764 4174 50766 4226
rect 50818 4174 50820 4226
rect 48188 3668 48244 3678
rect 47628 3574 47684 3612
rect 47740 3666 48244 3668
rect 47740 3614 48190 3666
rect 48242 3614 48244 3666
rect 47740 3612 48244 3614
rect 46844 3502 46846 3554
rect 46898 3502 46900 3554
rect 46844 3490 46900 3502
rect 47740 800 47796 3612
rect 48188 3602 48244 3612
rect 50540 3556 50596 3566
rect 50764 3556 50820 4174
rect 51772 3668 51828 3678
rect 50596 3500 50820 3556
rect 51324 3666 51828 3668
rect 51324 3614 51774 3666
rect 51826 3614 51828 3666
rect 51324 3612 51828 3614
rect 50540 3462 50596 3500
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 51324 800 51380 3612
rect 51772 3602 51828 3612
rect 54124 3554 54180 4508
rect 54348 4498 54404 4508
rect 55356 3668 55412 3678
rect 54124 3502 54126 3554
rect 54178 3502 54180 3554
rect 54124 3490 54180 3502
rect 54908 3666 55412 3668
rect 54908 3614 55358 3666
rect 55410 3614 55412 3666
rect 54908 3612 55412 3614
rect 54908 800 54964 3612
rect 55356 3602 55412 3612
rect 57260 3668 57316 31052
rect 59612 29428 59668 29438
rect 58268 3668 58324 3678
rect 59052 3668 59108 3678
rect 57260 3666 58324 3668
rect 57260 3614 58270 3666
rect 58322 3614 58324 3666
rect 57260 3612 58324 3614
rect 57260 3554 57316 3612
rect 58268 3602 58324 3612
rect 58492 3666 59108 3668
rect 58492 3614 59054 3666
rect 59106 3614 59108 3666
rect 58492 3612 59108 3614
rect 57260 3502 57262 3554
rect 57314 3502 57316 3554
rect 57260 3490 57316 3502
rect 58492 800 58548 3612
rect 59052 3602 59108 3612
rect 59612 3556 59668 29372
rect 59612 3490 59668 3500
rect 60956 3668 61012 32732
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 61964 3668 62020 3678
rect 60956 3666 62020 3668
rect 60956 3614 61966 3666
rect 62018 3614 62020 3666
rect 60956 3612 62020 3614
rect 60956 3554 61012 3612
rect 61964 3602 62020 3612
rect 62076 3668 62132 3678
rect 60956 3502 60958 3554
rect 61010 3502 61012 3554
rect 60956 3490 61012 3502
rect 62076 800 62132 3612
rect 62860 3668 62916 3678
rect 62860 3574 62916 3612
rect 65212 3668 65268 3678
rect 65212 3554 65268 3612
rect 65772 3668 65828 3678
rect 65772 3574 65828 3612
rect 66668 3666 66724 3678
rect 66668 3614 66670 3666
rect 66722 3614 66724 3666
rect 65212 3502 65214 3554
rect 65266 3502 65268 3554
rect 65212 3490 65268 3502
rect 65660 3444 65716 3454
rect 65660 800 65716 3388
rect 66668 3444 66724 3614
rect 68236 3668 68292 36204
rect 69580 34692 69636 34702
rect 68236 3602 68292 3612
rect 69244 3668 69300 3678
rect 68908 3556 68964 3566
rect 68908 3462 68964 3500
rect 66668 3378 66724 3388
rect 69244 800 69300 3612
rect 69580 3666 69636 34636
rect 73052 12740 73108 55916
rect 78092 55970 78148 57038
rect 81276 56476 81540 56486
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81276 56410 81540 56420
rect 78092 55918 78094 55970
rect 78146 55918 78148 55970
rect 78092 55906 78148 55918
rect 80444 56082 80500 56094
rect 80444 56030 80446 56082
rect 80498 56030 80500 56082
rect 80444 55972 80500 56030
rect 80444 55906 80500 55916
rect 81004 55972 81060 55982
rect 81004 55878 81060 55916
rect 82684 55970 82740 59200
rect 84924 56084 84980 56094
rect 84924 55990 84980 56028
rect 85708 56084 85764 56094
rect 82684 55918 82686 55970
rect 82738 55918 82740 55970
rect 82684 55906 82740 55918
rect 83132 55972 83188 55982
rect 74732 55298 74788 55310
rect 74732 55246 74734 55298
rect 74786 55246 74788 55298
rect 74732 55076 74788 55246
rect 75180 55076 75236 55086
rect 74732 55074 75236 55076
rect 74732 55022 75182 55074
rect 75234 55022 75236 55074
rect 74732 55020 75236 55022
rect 75180 14308 75236 55020
rect 81276 54908 81540 54918
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81276 54842 81540 54852
rect 81276 53340 81540 53350
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81276 53274 81540 53284
rect 81276 51772 81540 51782
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81276 51706 81540 51716
rect 81276 50204 81540 50214
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81276 50138 81540 50148
rect 81276 48636 81540 48646
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81276 48570 81540 48580
rect 81276 47068 81540 47078
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81276 47002 81540 47012
rect 81276 45500 81540 45510
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81276 45434 81540 45444
rect 81276 43932 81540 43942
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81276 43866 81540 43876
rect 81276 42364 81540 42374
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81276 42298 81540 42308
rect 81276 40796 81540 40806
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81276 40730 81540 40740
rect 81276 39228 81540 39238
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81276 39162 81540 39172
rect 81276 37660 81540 37670
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81276 37594 81540 37604
rect 81276 36092 81540 36102
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81276 36026 81540 36036
rect 81276 34524 81540 34534
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81276 34458 81540 34468
rect 81276 32956 81540 32966
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81276 32890 81540 32900
rect 81276 31388 81540 31398
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81276 31322 81540 31332
rect 81276 29820 81540 29830
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81276 29754 81540 29764
rect 81276 28252 81540 28262
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81276 28186 81540 28196
rect 81276 26684 81540 26694
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81276 26618 81540 26628
rect 81276 25116 81540 25126
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81276 25050 81540 25060
rect 81276 23548 81540 23558
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81276 23482 81540 23492
rect 81276 21980 81540 21990
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81276 21914 81540 21924
rect 81276 20412 81540 20422
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81276 20346 81540 20356
rect 75180 14242 75236 14252
rect 78652 19348 78708 19358
rect 73052 12674 73108 12684
rect 73388 11284 73444 11294
rect 71148 7588 71204 7598
rect 71148 4564 71204 7532
rect 71148 4562 71428 4564
rect 71148 4510 71150 4562
rect 71202 4510 71428 4562
rect 71148 4508 71428 4510
rect 71148 4498 71204 4508
rect 71372 4450 71428 4508
rect 71372 4398 71374 4450
rect 71426 4398 71428 4450
rect 71372 4386 71428 4398
rect 71708 4450 71764 4462
rect 71708 4398 71710 4450
rect 71762 4398 71764 4450
rect 69580 3614 69582 3666
rect 69634 3614 69636 3666
rect 69580 3556 69636 3614
rect 70476 3668 70532 3678
rect 70476 3574 70532 3612
rect 69580 3490 69636 3500
rect 71708 3556 71764 4398
rect 73388 3668 73444 11228
rect 74844 9268 74900 9278
rect 74844 4564 74900 9212
rect 74844 4562 75124 4564
rect 74844 4510 74846 4562
rect 74898 4510 75124 4562
rect 74844 4508 75124 4510
rect 74844 4498 74900 4508
rect 75068 4450 75124 4508
rect 75068 4398 75070 4450
rect 75122 4398 75124 4450
rect 75068 4386 75124 4398
rect 75404 4450 75460 4462
rect 75404 4398 75406 4450
rect 75458 4398 75460 4450
rect 75404 4340 75460 4398
rect 75404 4274 75460 4284
rect 76636 4340 76692 4350
rect 76636 4246 76692 4284
rect 71708 3490 71764 3500
rect 72828 3666 73444 3668
rect 72828 3614 73390 3666
rect 73442 3614 73444 3666
rect 72828 3612 73444 3614
rect 72828 3554 72884 3612
rect 73388 3602 73444 3612
rect 76412 4116 76468 4126
rect 72828 3502 72830 3554
rect 72882 3502 72884 3554
rect 72828 3490 72884 3502
rect 74060 3556 74116 3566
rect 74060 3462 74116 3500
rect 72940 3444 72996 3454
rect 72940 1652 72996 3388
rect 75628 3444 75684 3454
rect 75628 3350 75684 3388
rect 72828 1596 72996 1652
rect 72828 800 72884 1596
rect 76412 800 76468 4060
rect 77644 4116 77700 4126
rect 77644 4022 77700 4060
rect 78316 3668 78372 3678
rect 78652 3668 78708 19292
rect 81276 18844 81540 18854
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81276 18778 81540 18788
rect 83132 17668 83188 55916
rect 83132 17602 83188 17612
rect 85036 21028 85092 21038
rect 81276 17276 81540 17286
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81276 17210 81540 17220
rect 83132 15988 83188 15998
rect 81276 15708 81540 15718
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81276 15642 81540 15652
rect 81276 14140 81540 14150
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81276 14074 81540 14084
rect 81276 12572 81540 12582
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81276 12506 81540 12516
rect 81276 11004 81540 11014
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81276 10938 81540 10948
rect 81276 9436 81540 9446
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81276 9370 81540 9380
rect 81276 7868 81540 7878
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81276 7802 81540 7812
rect 81276 6300 81540 6310
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81276 6234 81540 6244
rect 81276 4732 81540 4742
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81276 4666 81540 4676
rect 83132 4452 83188 15932
rect 82908 4450 83188 4452
rect 82908 4398 83134 4450
rect 83186 4398 83188 4450
rect 82908 4396 83188 4398
rect 80220 4340 80276 4350
rect 78316 3666 78708 3668
rect 78316 3614 78318 3666
rect 78370 3614 78708 3666
rect 78316 3612 78708 3614
rect 78316 3602 78372 3612
rect 78652 3554 78708 3612
rect 78652 3502 78654 3554
rect 78706 3502 78708 3554
rect 78652 3490 78708 3502
rect 78988 4338 80276 4340
rect 78988 4286 80222 4338
rect 80274 4286 80276 4338
rect 78988 4284 80276 4286
rect 78988 3442 79044 4284
rect 80220 4274 80276 4284
rect 78988 3390 78990 3442
rect 79042 3390 79044 3442
rect 78988 3378 79044 3390
rect 79996 4116 80052 4126
rect 79996 800 80052 4060
rect 81228 4116 81284 4126
rect 81228 4022 81284 4060
rect 82908 3666 82964 4396
rect 83132 4386 83188 4396
rect 83468 4450 83524 4462
rect 83468 4398 83470 4450
rect 83522 4398 83524 4450
rect 83468 4340 83524 4398
rect 85036 4452 85092 20972
rect 85708 11172 85764 56028
rect 88060 55972 88116 59200
rect 91868 56084 91924 56094
rect 92428 56084 92484 56094
rect 91868 56082 92484 56084
rect 91868 56030 91870 56082
rect 91922 56030 92430 56082
rect 92482 56030 92484 56082
rect 91868 56028 92484 56030
rect 91868 56018 91924 56028
rect 88060 55906 88116 55916
rect 89516 55972 89572 55982
rect 89516 55878 89572 55916
rect 91644 55524 91700 55534
rect 85708 11106 85764 11116
rect 88732 22932 88788 22942
rect 86716 4452 86772 4462
rect 85036 4386 85092 4396
rect 86492 4396 86716 4452
rect 83804 4340 83860 4350
rect 83468 4338 83860 4340
rect 83468 4286 83806 4338
rect 83858 4286 83860 4338
rect 83468 4284 83860 4286
rect 83804 4274 83860 4284
rect 82908 3614 82910 3666
rect 82962 3614 82964 3666
rect 82908 3602 82964 3614
rect 83580 4116 83636 4126
rect 81276 3164 81540 3174
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81276 3098 81540 3108
rect 83580 800 83636 4060
rect 84812 4116 84868 4126
rect 84812 4022 84868 4060
rect 86492 3666 86548 4396
rect 86716 4358 86772 4396
rect 87052 4450 87108 4462
rect 87052 4398 87054 4450
rect 87106 4398 87108 4450
rect 87052 4340 87108 4398
rect 87052 4274 87108 4284
rect 87948 4340 88004 4350
rect 87948 4246 88004 4284
rect 86492 3614 86494 3666
rect 86546 3614 86548 3666
rect 86492 3602 86548 3614
rect 87164 4228 87220 4238
rect 87164 800 87220 4172
rect 88732 3666 88788 22876
rect 91644 4564 91700 55468
rect 92428 21028 92484 56028
rect 93436 55972 93492 59200
rect 96236 56082 96292 56094
rect 96236 56030 96238 56082
rect 96290 56030 96292 56082
rect 93884 55972 93940 55982
rect 93436 55970 93940 55972
rect 93436 55918 93886 55970
rect 93938 55918 93940 55970
rect 93436 55916 93940 55918
rect 93884 55906 93940 55916
rect 96236 55972 96292 56030
rect 96236 55906 96292 55916
rect 97132 55972 97188 55982
rect 97132 55878 97188 55916
rect 96636 55692 96900 55702
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96636 55626 96900 55636
rect 98812 55412 98868 59200
rect 98812 55346 98868 55356
rect 99932 55972 99988 55982
rect 104188 55972 104244 59200
rect 109564 56308 109620 59200
rect 114940 56642 114996 59200
rect 114940 56590 114942 56642
rect 114994 56590 114996 56642
rect 114940 56578 114996 56590
rect 115500 56642 115556 56654
rect 115500 56590 115502 56642
rect 115554 56590 115556 56642
rect 111996 56476 112260 56486
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 111996 56410 112260 56420
rect 109788 56308 109844 56318
rect 109564 56306 109844 56308
rect 109564 56254 109566 56306
rect 109618 56254 109790 56306
rect 109842 56254 109844 56306
rect 109564 56252 109844 56254
rect 109564 56242 109620 56252
rect 109788 56242 109844 56252
rect 115500 56306 115556 56590
rect 115500 56254 115502 56306
rect 115554 56254 115556 56306
rect 115500 56242 115556 56254
rect 115948 56642 116004 56654
rect 115948 56590 115950 56642
rect 116002 56590 116004 56642
rect 115948 56306 116004 56590
rect 115948 56254 115950 56306
rect 116002 56254 116004 56306
rect 115948 56242 116004 56254
rect 120316 56308 120372 59200
rect 120540 56308 120596 56318
rect 120316 56306 120596 56308
rect 120316 56254 120318 56306
rect 120370 56254 120542 56306
rect 120594 56254 120596 56306
rect 120316 56252 120596 56254
rect 120316 56242 120372 56252
rect 120540 56242 120596 56252
rect 125692 56308 125748 59200
rect 131068 57092 131124 59200
rect 130732 57036 131348 57092
rect 125916 56308 125972 56318
rect 125692 56306 125972 56308
rect 125692 56254 125694 56306
rect 125746 56254 125918 56306
rect 125970 56254 125972 56306
rect 125692 56252 125972 56254
rect 125692 56242 125748 56252
rect 125916 56242 125972 56252
rect 130732 56306 130788 57036
rect 130732 56254 130734 56306
rect 130786 56254 130788 56306
rect 130732 56242 130788 56254
rect 126252 56196 126308 56206
rect 126252 56102 126308 56140
rect 127820 56196 127876 56206
rect 107100 56084 107156 56094
rect 107660 56084 107716 56094
rect 107100 56082 107716 56084
rect 107100 56030 107102 56082
rect 107154 56030 107662 56082
rect 107714 56030 107716 56082
rect 107100 56028 107716 56030
rect 107100 56018 107156 56028
rect 104748 55972 104804 55982
rect 104188 55970 104804 55972
rect 104188 55918 104750 55970
rect 104802 55918 104804 55970
rect 104188 55916 104804 55918
rect 96636 54124 96900 54134
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96636 54058 96900 54068
rect 96636 52556 96900 52566
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96636 52490 96900 52500
rect 96636 50988 96900 50998
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96636 50922 96900 50932
rect 96636 49420 96900 49430
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96636 49354 96900 49364
rect 96636 47852 96900 47862
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96636 47786 96900 47796
rect 96636 46284 96900 46294
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96636 46218 96900 46228
rect 96636 44716 96900 44726
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96636 44650 96900 44660
rect 96636 43148 96900 43158
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96636 43082 96900 43092
rect 96636 41580 96900 41590
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96636 41514 96900 41524
rect 96636 40012 96900 40022
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96636 39946 96900 39956
rect 96636 38444 96900 38454
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96636 38378 96900 38388
rect 96636 36876 96900 36886
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96636 36810 96900 36820
rect 96636 35308 96900 35318
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96636 35242 96900 35252
rect 96636 33740 96900 33750
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96636 33674 96900 33684
rect 96636 32172 96900 32182
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96636 32106 96900 32116
rect 96636 30604 96900 30614
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96636 30538 96900 30548
rect 96636 29036 96900 29046
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96636 28970 96900 28980
rect 96636 27468 96900 27478
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96636 27402 96900 27412
rect 96636 25900 96900 25910
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96636 25834 96900 25844
rect 96636 24332 96900 24342
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96636 24266 96900 24276
rect 96636 22764 96900 22774
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96636 22698 96900 22708
rect 96636 21196 96900 21206
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96636 21130 96900 21140
rect 92428 20962 92484 20972
rect 96636 19628 96900 19638
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96636 19562 96900 19572
rect 96636 18060 96900 18070
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96636 17994 96900 18004
rect 96636 16492 96900 16502
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96636 16426 96900 16436
rect 96636 14924 96900 14934
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96636 14858 96900 14868
rect 96636 13356 96900 13366
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96636 13290 96900 13300
rect 96636 11788 96900 11798
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96636 11722 96900 11732
rect 96636 10220 96900 10230
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96636 10154 96900 10164
rect 99932 9268 99988 55916
rect 104748 55906 104804 55916
rect 100044 55412 100100 55422
rect 100044 55318 100100 55356
rect 102284 55298 102340 55310
rect 102284 55246 102286 55298
rect 102338 55246 102340 55298
rect 102284 55076 102340 55246
rect 102732 55076 102788 55086
rect 102284 55074 102788 55076
rect 102284 55022 102734 55074
rect 102786 55022 102788 55074
rect 102284 55020 102788 55022
rect 102508 49588 102564 55020
rect 102732 55010 102788 55020
rect 102508 49522 102564 49532
rect 107660 15988 107716 56028
rect 110348 55970 110404 55982
rect 110348 55918 110350 55970
rect 110402 55918 110404 55970
rect 110348 55188 110404 55918
rect 110348 55122 110404 55132
rect 116508 55970 116564 55982
rect 116508 55918 116510 55970
rect 116562 55918 116564 55970
rect 111996 54908 112260 54918
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 111996 54842 112260 54852
rect 111996 53340 112260 53350
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 111996 53274 112260 53284
rect 116508 52164 116564 55918
rect 121100 55972 121156 55982
rect 121100 55878 121156 55916
rect 127356 55692 127620 55702
rect 127412 55636 127460 55692
rect 127516 55636 127564 55692
rect 127356 55626 127620 55636
rect 127356 54124 127620 54134
rect 127412 54068 127460 54124
rect 127516 54068 127564 54124
rect 127356 54058 127620 54068
rect 127820 52836 127876 56140
rect 131292 56194 131348 57036
rect 136444 56420 136500 59200
rect 141820 57204 141876 59200
rect 141820 57148 142212 57204
rect 136444 56364 136948 56420
rect 136444 56306 136500 56364
rect 136444 56254 136446 56306
rect 136498 56254 136500 56306
rect 136444 56242 136500 56254
rect 131292 56142 131294 56194
rect 131346 56142 131348 56194
rect 131292 56130 131348 56142
rect 131628 56194 131684 56206
rect 131628 56142 131630 56194
rect 131682 56142 131684 56194
rect 131628 55468 131684 56142
rect 135772 56196 135828 56206
rect 131628 55412 131796 55468
rect 130284 54404 130340 54414
rect 130284 53730 130340 54348
rect 131740 54404 131796 55412
rect 132972 55300 133028 55310
rect 132972 54740 133028 55244
rect 135100 55300 135156 55310
rect 135100 55206 135156 55244
rect 132524 54738 133028 54740
rect 132524 54686 132974 54738
rect 133026 54686 133028 54738
rect 132524 54684 133028 54686
rect 132524 54514 132580 54684
rect 132972 54674 133028 54684
rect 135772 55186 135828 56140
rect 136668 56196 136724 56206
rect 136668 56102 136724 56140
rect 136892 56082 136948 56364
rect 142156 56306 142212 57148
rect 142716 56476 142980 56486
rect 142772 56420 142820 56476
rect 142876 56420 142924 56476
rect 142716 56410 142980 56420
rect 147196 56420 147252 59200
rect 142156 56254 142158 56306
rect 142210 56254 142212 56306
rect 142156 56196 142212 56254
rect 147196 56364 147700 56420
rect 147196 56306 147252 56364
rect 147196 56254 147198 56306
rect 147250 56254 147252 56306
rect 147196 56242 147252 56254
rect 142156 56130 142212 56140
rect 142604 56194 142660 56206
rect 142604 56142 142606 56194
rect 142658 56142 142660 56194
rect 136892 56030 136894 56082
rect 136946 56030 136948 56082
rect 136892 56018 136948 56030
rect 141260 55412 141316 55422
rect 141036 55356 141260 55412
rect 138348 55300 138404 55310
rect 138348 55206 138404 55244
rect 140476 55300 140532 55310
rect 140476 55206 140532 55244
rect 135772 55134 135774 55186
rect 135826 55134 135828 55186
rect 135772 54738 135828 55134
rect 135772 54686 135774 54738
rect 135826 54686 135828 54738
rect 135772 54674 135828 54686
rect 141036 54738 141092 55356
rect 141260 55318 141316 55356
rect 142604 55412 142660 56142
rect 142828 56196 142884 56206
rect 142828 56082 142884 56140
rect 142828 56030 142830 56082
rect 142882 56030 142884 56082
rect 142828 56018 142884 56030
rect 147420 56194 147476 56206
rect 147420 56142 147422 56194
rect 147474 56142 147476 56194
rect 142604 55346 142660 55356
rect 143836 55300 143892 55310
rect 143836 55206 143892 55244
rect 142716 54908 142980 54918
rect 142772 54852 142820 54908
rect 142876 54852 142924 54908
rect 142716 54842 142980 54852
rect 141036 54686 141038 54738
rect 141090 54686 141092 54738
rect 141036 54674 141092 54686
rect 132524 54462 132526 54514
rect 132578 54462 132580 54514
rect 132524 54450 132580 54462
rect 131740 54310 131796 54348
rect 145964 54404 146020 54414
rect 130284 53678 130286 53730
rect 130338 53678 130340 53730
rect 130284 53666 130340 53678
rect 134988 54290 135044 54302
rect 134988 54238 134990 54290
rect 135042 54238 135044 54290
rect 127820 52770 127876 52780
rect 129388 53618 129444 53630
rect 129388 53566 129390 53618
rect 129442 53566 129444 53618
rect 127356 52556 127620 52566
rect 127412 52500 127460 52556
rect 127516 52500 127564 52556
rect 127356 52490 127620 52500
rect 116508 52098 116564 52108
rect 111996 51772 112260 51782
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 111996 51706 112260 51716
rect 127356 50988 127620 50998
rect 127412 50932 127460 50988
rect 127516 50932 127564 50988
rect 127356 50922 127620 50932
rect 111996 50204 112260 50214
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 111996 50138 112260 50148
rect 127356 49420 127620 49430
rect 127412 49364 127460 49420
rect 127516 49364 127564 49420
rect 127356 49354 127620 49364
rect 111996 48636 112260 48646
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 111996 48570 112260 48580
rect 127356 47852 127620 47862
rect 127412 47796 127460 47852
rect 127516 47796 127564 47852
rect 127356 47786 127620 47796
rect 111996 47068 112260 47078
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 111996 47002 112260 47012
rect 127356 46284 127620 46294
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127356 46218 127620 46228
rect 111996 45500 112260 45510
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 111996 45434 112260 45444
rect 127356 44716 127620 44726
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127356 44650 127620 44660
rect 111996 43932 112260 43942
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 111996 43866 112260 43876
rect 127356 43148 127620 43158
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127356 43082 127620 43092
rect 111996 42364 112260 42374
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 111996 42298 112260 42308
rect 127356 41580 127620 41590
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127356 41514 127620 41524
rect 111996 40796 112260 40806
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 111996 40730 112260 40740
rect 127356 40012 127620 40022
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127356 39946 127620 39956
rect 111996 39228 112260 39238
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 111996 39162 112260 39172
rect 127356 38444 127620 38454
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127356 38378 127620 38388
rect 111996 37660 112260 37670
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 111996 37594 112260 37604
rect 127356 36876 127620 36886
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127356 36810 127620 36820
rect 111996 36092 112260 36102
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 111996 36026 112260 36036
rect 127356 35308 127620 35318
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127356 35242 127620 35252
rect 111996 34524 112260 34534
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 111996 34458 112260 34468
rect 127356 33740 127620 33750
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127356 33674 127620 33684
rect 111996 32956 112260 32966
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 111996 32890 112260 32900
rect 127356 32172 127620 32182
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127356 32106 127620 32116
rect 111996 31388 112260 31398
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 111996 31322 112260 31332
rect 127356 30604 127620 30614
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127356 30538 127620 30548
rect 111996 29820 112260 29830
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 111996 29754 112260 29764
rect 127356 29036 127620 29046
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127356 28970 127620 28980
rect 111996 28252 112260 28262
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 111996 28186 112260 28196
rect 127356 27468 127620 27478
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127356 27402 127620 27412
rect 111996 26684 112260 26694
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 111996 26618 112260 26628
rect 127356 25900 127620 25910
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127356 25834 127620 25844
rect 111996 25116 112260 25126
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 111996 25050 112260 25060
rect 129388 24500 129444 53566
rect 134988 31948 135044 54238
rect 134876 31892 135044 31948
rect 140252 54290 140308 54302
rect 140252 54238 140254 54290
rect 140306 54238 140308 54290
rect 134876 26068 134932 31892
rect 140252 29428 140308 54238
rect 145964 53730 146020 54348
rect 147420 54404 147476 56142
rect 147644 56082 147700 56364
rect 152572 56308 152628 59200
rect 157388 57090 157444 57102
rect 157388 57038 157390 57090
rect 157442 57038 157444 57090
rect 152572 56306 152852 56308
rect 152572 56254 152574 56306
rect 152626 56254 152852 56306
rect 152572 56252 152852 56254
rect 152572 56242 152628 56252
rect 152796 56194 152852 56252
rect 157388 56306 157444 57038
rect 157948 57090 158004 59200
rect 157948 57038 157950 57090
rect 158002 57038 158004 57090
rect 157948 57026 158004 57038
rect 158508 57090 158564 57102
rect 158508 57038 158510 57090
rect 158562 57038 158564 57090
rect 157388 56254 157390 56306
rect 157442 56254 157444 56306
rect 157388 56242 157444 56254
rect 152796 56142 152798 56194
rect 152850 56142 152852 56194
rect 152796 56130 152852 56142
rect 153132 56194 153188 56206
rect 158172 56196 158228 56206
rect 153132 56142 153134 56194
rect 153186 56142 153188 56194
rect 147644 56030 147646 56082
rect 147698 56030 147700 56082
rect 147644 56018 147700 56030
rect 147868 55300 147924 55310
rect 147868 55188 147924 55244
rect 152684 55298 152740 55310
rect 152684 55246 152686 55298
rect 152738 55246 152740 55298
rect 147868 55186 148148 55188
rect 147868 55134 147870 55186
rect 147922 55134 148148 55186
rect 147868 55132 148148 55134
rect 147868 55122 147924 55132
rect 148092 54740 148148 55132
rect 152684 55076 152740 55246
rect 152684 55010 152740 55020
rect 148092 54514 148148 54684
rect 148652 54740 148708 54750
rect 148652 54646 148708 54684
rect 150108 54740 150164 54750
rect 150108 54646 150164 54684
rect 148092 54462 148094 54514
rect 148146 54462 148148 54514
rect 148092 54450 148148 54462
rect 147420 54310 147476 54348
rect 151564 54404 151620 54414
rect 145964 53678 145966 53730
rect 146018 53678 146020 53730
rect 145964 53666 146020 53678
rect 151564 53730 151620 54348
rect 153132 54404 153188 56142
rect 157500 56194 158228 56196
rect 157500 56142 158174 56194
rect 158226 56142 158228 56194
rect 157500 56140 158228 56142
rect 157500 55468 157556 56140
rect 158172 56130 158228 56140
rect 158508 56194 158564 57038
rect 163324 56420 163380 59200
rect 168700 56642 168756 59200
rect 168700 56590 168702 56642
rect 168754 56590 168756 56642
rect 163324 56364 163828 56420
rect 163324 56306 163380 56364
rect 163324 56254 163326 56306
rect 163378 56254 163380 56306
rect 163324 56242 163380 56254
rect 158508 56142 158510 56194
rect 158562 56142 158564 56194
rect 158508 56130 158564 56142
rect 163548 56194 163604 56206
rect 163548 56142 163550 56194
rect 163602 56142 163604 56194
rect 158076 55692 158340 55702
rect 158132 55636 158180 55692
rect 158236 55636 158284 55692
rect 158076 55626 158340 55636
rect 163548 55468 163604 56142
rect 163772 56082 163828 56364
rect 168700 56308 168756 56590
rect 169596 56642 169652 56654
rect 169596 56590 169598 56642
rect 169650 56590 169652 56642
rect 168812 56308 168868 56318
rect 168700 56306 168868 56308
rect 168700 56254 168814 56306
rect 168866 56254 168868 56306
rect 168700 56252 168868 56254
rect 168812 56242 168868 56252
rect 163772 56030 163774 56082
rect 163826 56030 163828 56082
rect 163772 56018 163828 56030
rect 169260 56194 169316 56206
rect 169260 56142 169262 56194
rect 169314 56142 169316 56194
rect 169260 55468 169316 56142
rect 169596 56194 169652 56590
rect 173436 56476 173700 56486
rect 173492 56420 173540 56476
rect 173596 56420 173644 56476
rect 173436 56410 173700 56420
rect 174076 56420 174132 59200
rect 174076 56364 174580 56420
rect 174076 56306 174132 56364
rect 174076 56254 174078 56306
rect 174130 56254 174132 56306
rect 174076 56242 174132 56254
rect 169596 56142 169598 56194
rect 169650 56142 169652 56194
rect 169596 56130 169652 56142
rect 174300 56194 174356 56206
rect 174300 56142 174302 56194
rect 174354 56142 174356 56194
rect 153916 55412 153972 55422
rect 153244 55076 153300 55086
rect 153244 54982 153300 55020
rect 153916 54740 153972 55356
rect 156268 55412 156324 55422
rect 156268 55318 156324 55356
rect 156716 55412 156772 55422
rect 156716 55298 156772 55356
rect 156716 55246 156718 55298
rect 156770 55246 156772 55298
rect 156716 55234 156772 55246
rect 157388 55412 157556 55468
rect 161868 55412 161924 55422
rect 157388 55186 157444 55412
rect 161868 55318 161924 55356
rect 162428 55412 162484 55422
rect 162428 55298 162484 55356
rect 162428 55246 162430 55298
rect 162482 55246 162484 55298
rect 162428 55234 162484 55246
rect 163212 55412 163604 55468
rect 168924 55412 169316 55468
rect 157388 55134 157390 55186
rect 157442 55134 157444 55186
rect 153916 54514 153972 54684
rect 157164 54740 157220 54750
rect 157388 54740 157444 55134
rect 163212 55186 163268 55412
rect 163212 55134 163214 55186
rect 163266 55134 163268 55186
rect 157164 54738 157444 54740
rect 157164 54686 157166 54738
rect 157218 54686 157444 54738
rect 157164 54684 157444 54686
rect 162316 54740 162372 54750
rect 157164 54674 157220 54684
rect 162316 54646 162372 54684
rect 163212 54740 163268 55134
rect 168924 55186 168980 55412
rect 169708 55300 169764 55310
rect 169708 55206 169764 55244
rect 170380 55300 170436 55310
rect 170380 55206 170436 55244
rect 168924 55134 168926 55186
rect 168978 55134 168980 55186
rect 163212 54674 163268 54684
rect 166236 55076 166292 55086
rect 153916 54462 153918 54514
rect 153970 54462 153972 54514
rect 153916 54450 153972 54462
rect 153132 54310 153188 54348
rect 151564 53678 151566 53730
rect 151618 53678 151620 53730
rect 151564 53666 151620 53678
rect 156380 54290 156436 54302
rect 156380 54238 156382 54290
rect 156434 54238 156436 54290
rect 145180 53506 145236 53518
rect 145180 53454 145182 53506
rect 145234 53454 145236 53506
rect 142716 53340 142980 53350
rect 142772 53284 142820 53340
rect 142876 53284 142924 53340
rect 142716 53274 142980 53284
rect 142716 51772 142980 51782
rect 142772 51716 142820 51772
rect 142876 51716 142924 51772
rect 142716 51706 142980 51716
rect 142716 50204 142980 50214
rect 142772 50148 142820 50204
rect 142876 50148 142924 50204
rect 142716 50138 142980 50148
rect 142716 48636 142980 48646
rect 142772 48580 142820 48636
rect 142876 48580 142924 48636
rect 142716 48570 142980 48580
rect 142716 47068 142980 47078
rect 142772 47012 142820 47068
rect 142876 47012 142924 47068
rect 142716 47002 142980 47012
rect 142716 45500 142980 45510
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142716 45434 142980 45444
rect 142716 43932 142980 43942
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142716 43866 142980 43876
rect 142716 42364 142980 42374
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142716 42298 142980 42308
rect 145180 41188 145236 53454
rect 145180 41122 145236 41132
rect 150780 53506 150836 53518
rect 150780 53454 150782 53506
rect 150834 53454 150836 53506
rect 142716 40796 142980 40806
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142716 40730 142980 40740
rect 142716 39228 142980 39238
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142716 39162 142980 39172
rect 142716 37660 142980 37670
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142716 37594 142980 37604
rect 142716 36092 142980 36102
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142716 36026 142980 36036
rect 142716 34524 142980 34534
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142716 34458 142980 34468
rect 142716 32956 142980 32966
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142716 32890 142980 32900
rect 142716 31388 142980 31398
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142716 31322 142980 31332
rect 150780 31108 150836 53454
rect 156380 32788 156436 54238
rect 161532 54290 161588 54302
rect 161532 54238 161534 54290
rect 161586 54238 161588 54290
rect 158076 54124 158340 54134
rect 158132 54068 158180 54124
rect 158236 54068 158284 54124
rect 158076 54058 158340 54068
rect 158076 52556 158340 52566
rect 158132 52500 158180 52556
rect 158236 52500 158284 52556
rect 158076 52490 158340 52500
rect 158076 50988 158340 50998
rect 158132 50932 158180 50988
rect 158236 50932 158284 50988
rect 158076 50922 158340 50932
rect 158076 49420 158340 49430
rect 158132 49364 158180 49420
rect 158236 49364 158284 49420
rect 158076 49354 158340 49364
rect 158076 47852 158340 47862
rect 158132 47796 158180 47852
rect 158236 47796 158284 47852
rect 158076 47786 158340 47796
rect 158076 46284 158340 46294
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158076 46218 158340 46228
rect 158076 44716 158340 44726
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158076 44650 158340 44660
rect 158076 43148 158340 43158
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158076 43082 158340 43092
rect 158076 41580 158340 41590
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158076 41514 158340 41524
rect 158076 40012 158340 40022
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158076 39946 158340 39956
rect 158076 38444 158340 38454
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158076 38378 158340 38388
rect 158076 36876 158340 36886
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158076 36810 158340 36820
rect 161532 36260 161588 54238
rect 161980 53732 162036 53742
rect 162428 53732 162484 53742
rect 161980 53730 162484 53732
rect 161980 53678 161982 53730
rect 162034 53678 162430 53730
rect 162482 53678 162484 53730
rect 161980 53676 162484 53678
rect 161980 52052 162036 53676
rect 162428 53666 162484 53676
rect 166236 53620 166292 55020
rect 167916 54740 167972 54750
rect 167916 54646 167972 54684
rect 168924 54740 168980 55134
rect 174300 55186 174356 56142
rect 174524 56082 174580 56364
rect 179452 56308 179508 59200
rect 184828 56420 184884 59200
rect 190204 56642 190260 59200
rect 190204 56590 190206 56642
rect 190258 56590 190260 56642
rect 190204 56578 190260 56590
rect 191436 56642 191492 56654
rect 191436 56590 191438 56642
rect 191490 56590 191492 56642
rect 184828 56364 185332 56420
rect 179452 56306 179732 56308
rect 179452 56254 179454 56306
rect 179506 56254 179732 56306
rect 179452 56252 179732 56254
rect 179452 56242 179508 56252
rect 179676 56194 179732 56252
rect 184828 56306 184884 56364
rect 184828 56254 184830 56306
rect 184882 56254 184884 56306
rect 184828 56242 184884 56254
rect 179676 56142 179678 56194
rect 179730 56142 179732 56194
rect 179676 56130 179732 56142
rect 180012 56194 180068 56206
rect 180012 56142 180014 56194
rect 180066 56142 180068 56194
rect 174524 56030 174526 56082
rect 174578 56030 174580 56082
rect 174524 56018 174580 56030
rect 180012 55468 180068 56142
rect 184044 56196 184100 56206
rect 183372 55860 183428 55870
rect 180012 55412 180292 55468
rect 180236 55410 180292 55412
rect 180236 55358 180238 55410
rect 180290 55358 180292 55410
rect 180236 55346 180292 55358
rect 182364 55412 182420 55422
rect 182364 55318 182420 55356
rect 174972 55300 175028 55310
rect 174972 55206 175028 55244
rect 175532 55300 175588 55310
rect 175532 55206 175588 55244
rect 179452 55300 179508 55310
rect 174300 55134 174302 55186
rect 174354 55134 174356 55186
rect 173436 54908 173700 54918
rect 173492 54852 173540 54908
rect 173596 54852 173644 54908
rect 173436 54842 173700 54852
rect 168924 54674 168980 54684
rect 172732 54740 172788 54750
rect 172732 54646 172788 54684
rect 174300 54740 174356 55134
rect 174300 54674 174356 54684
rect 166236 53554 166292 53564
rect 167132 54290 167188 54302
rect 167132 54238 167134 54290
rect 167186 54238 167188 54290
rect 161980 51986 162036 51996
rect 161532 36194 161588 36204
rect 158076 35308 158340 35318
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158076 35242 158340 35252
rect 167132 34692 167188 54238
rect 171948 54290 172004 54302
rect 171948 54238 171950 54290
rect 172002 54238 172004 54290
rect 167468 53620 167524 53630
rect 167468 53526 167524 53564
rect 167132 34626 167188 34636
rect 158076 33740 158340 33750
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158076 33674 158340 33684
rect 156380 32722 156436 32732
rect 158076 32172 158340 32182
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158076 32106 158340 32116
rect 150780 31042 150836 31052
rect 158076 30604 158340 30614
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158076 30538 158340 30548
rect 142716 29820 142980 29830
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142716 29754 142980 29764
rect 140252 29362 140308 29372
rect 158076 29036 158340 29046
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158076 28970 158340 28980
rect 142716 28252 142980 28262
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142716 28186 142980 28196
rect 158076 27468 158340 27478
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158076 27402 158340 27412
rect 142716 26684 142980 26694
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142716 26618 142980 26628
rect 134876 26002 134932 26012
rect 158076 25900 158340 25910
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158076 25834 158340 25844
rect 142716 25116 142980 25126
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142716 25050 142980 25060
rect 129388 24434 129444 24444
rect 127356 24332 127620 24342
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127356 24266 127620 24276
rect 158076 24332 158340 24342
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158076 24266 158340 24276
rect 111996 23548 112260 23558
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 111996 23482 112260 23492
rect 142716 23548 142980 23558
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142716 23482 142980 23492
rect 127356 22764 127620 22774
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127356 22698 127620 22708
rect 158076 22764 158340 22774
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158076 22698 158340 22708
rect 111996 21980 112260 21990
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 111996 21914 112260 21924
rect 142716 21980 142980 21990
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142716 21914 142980 21924
rect 127356 21196 127620 21206
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127356 21130 127620 21140
rect 158076 21196 158340 21206
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158076 21130 158340 21140
rect 111996 20412 112260 20422
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 111996 20346 112260 20356
rect 142716 20412 142980 20422
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142716 20346 142980 20356
rect 127356 19628 127620 19638
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127356 19562 127620 19572
rect 158076 19628 158340 19638
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158076 19562 158340 19572
rect 111996 18844 112260 18854
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 111996 18778 112260 18788
rect 142716 18844 142980 18854
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142716 18778 142980 18788
rect 127356 18060 127620 18070
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127356 17994 127620 18004
rect 158076 18060 158340 18070
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158076 17994 158340 18004
rect 111996 17276 112260 17286
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 111996 17210 112260 17220
rect 142716 17276 142980 17286
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142716 17210 142980 17220
rect 127356 16492 127620 16502
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127356 16426 127620 16436
rect 158076 16492 158340 16502
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158076 16426 158340 16436
rect 107660 15922 107716 15932
rect 111996 15708 112260 15718
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 111996 15642 112260 15652
rect 142716 15708 142980 15718
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142716 15642 142980 15652
rect 127356 14924 127620 14934
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127356 14858 127620 14868
rect 158076 14924 158340 14934
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158076 14858 158340 14868
rect 111996 14140 112260 14150
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 111996 14074 112260 14084
rect 142716 14140 142980 14150
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142716 14074 142980 14084
rect 127356 13356 127620 13366
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127356 13290 127620 13300
rect 158076 13356 158340 13366
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158076 13290 158340 13300
rect 111996 12572 112260 12582
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 111996 12506 112260 12516
rect 142716 12572 142980 12582
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142716 12506 142980 12516
rect 127356 11788 127620 11798
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127356 11722 127620 11732
rect 158076 11788 158340 11798
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158076 11722 158340 11732
rect 171948 11284 172004 54238
rect 179452 53844 179508 55244
rect 182812 55074 182868 55086
rect 182812 55022 182814 55074
rect 182866 55022 182868 55074
rect 182812 54404 182868 55022
rect 183260 54514 183316 54526
rect 183260 54462 183262 54514
rect 183314 54462 183316 54514
rect 182924 54404 182980 54414
rect 183260 54404 183316 54462
rect 182812 54402 183316 54404
rect 182812 54350 182926 54402
rect 182978 54350 183316 54402
rect 182812 54348 183316 54350
rect 179452 53778 179508 53788
rect 180124 53844 180180 53854
rect 180124 53750 180180 53788
rect 182140 53844 182196 53854
rect 178108 53730 178164 53742
rect 178108 53678 178110 53730
rect 178162 53678 178164 53730
rect 177660 53620 177716 53630
rect 177660 53526 177716 53564
rect 178108 53620 178164 53678
rect 178108 53554 178164 53564
rect 173436 53340 173700 53350
rect 173492 53284 173540 53340
rect 173596 53284 173644 53340
rect 173436 53274 173700 53284
rect 182140 53172 182196 53788
rect 182812 53844 182868 54348
rect 182924 54338 182980 54348
rect 182812 53778 182868 53788
rect 183372 53508 183428 55804
rect 184044 54626 184100 56140
rect 185052 56196 185108 56206
rect 185052 56102 185108 56140
rect 185276 56082 185332 56364
rect 185276 56030 185278 56082
rect 185330 56030 185332 56082
rect 185276 56018 185332 56030
rect 187180 56196 187236 56206
rect 186172 55412 186228 55422
rect 186172 55318 186228 55356
rect 186396 55412 186452 55422
rect 186396 55318 186452 55356
rect 184044 54574 184046 54626
rect 184098 54574 184100 54626
rect 184044 54562 184100 54574
rect 186060 55298 186116 55310
rect 186060 55246 186062 55298
rect 186114 55246 186116 55298
rect 186060 54404 186116 55246
rect 187180 55298 187236 56140
rect 189868 56196 189924 56206
rect 189868 56102 189924 56140
rect 191212 56194 191268 56206
rect 191212 56142 191214 56194
rect 191266 56142 191268 56194
rect 190876 56084 190932 56094
rect 190876 55990 190932 56028
rect 187852 55972 187908 55982
rect 187852 55878 187908 55916
rect 188524 55970 188580 55982
rect 188524 55918 188526 55970
rect 188578 55918 188580 55970
rect 188524 55468 188580 55918
rect 189084 55972 189140 55982
rect 189084 55878 189140 55916
rect 188796 55692 189060 55702
rect 188852 55636 188900 55692
rect 188956 55636 189004 55692
rect 188796 55626 189060 55636
rect 191212 55468 191268 56142
rect 191436 56082 191492 56590
rect 192220 56642 192276 56654
rect 192220 56590 192222 56642
rect 192274 56590 192276 56642
rect 192220 56306 192276 56590
rect 195580 56420 195636 59200
rect 195580 56364 196196 56420
rect 192220 56254 192222 56306
rect 192274 56254 192276 56306
rect 192220 56242 192276 56254
rect 195468 56308 195524 56318
rect 195580 56308 195636 56364
rect 195468 56306 195636 56308
rect 195468 56254 195470 56306
rect 195522 56254 195636 56306
rect 195468 56252 195636 56254
rect 195468 56242 195524 56252
rect 193900 56196 193956 56206
rect 191436 56030 191438 56082
rect 191490 56030 191492 56082
rect 191436 56018 191492 56030
rect 191772 56084 191828 56094
rect 188300 55412 188356 55422
rect 188524 55412 188692 55468
rect 188300 55318 188356 55356
rect 187180 55246 187182 55298
rect 187234 55246 187236 55298
rect 187180 55234 187236 55246
rect 186508 55188 186564 55198
rect 186844 55188 186900 55198
rect 186508 55186 186900 55188
rect 186508 55134 186510 55186
rect 186562 55134 186846 55186
rect 186898 55134 186900 55186
rect 186508 55132 186900 55134
rect 186508 55122 186564 55132
rect 186844 55122 186900 55132
rect 186956 55188 187012 55198
rect 186956 55094 187012 55132
rect 187516 55188 187572 55198
rect 187516 55094 187572 55132
rect 187964 55074 188020 55086
rect 187964 55022 187966 55074
rect 188018 55022 188020 55074
rect 186172 54404 186228 54414
rect 186060 54402 186228 54404
rect 186060 54350 186174 54402
rect 186226 54350 186228 54402
rect 186060 54348 186228 54350
rect 186172 54338 186228 54348
rect 183372 53442 183428 53452
rect 186508 53732 186564 53742
rect 182476 53172 182532 53182
rect 182140 53170 182476 53172
rect 182140 53118 182142 53170
rect 182194 53118 182476 53170
rect 182140 53116 182476 53118
rect 182140 53106 182196 53116
rect 182476 52946 182532 53116
rect 185836 53172 185892 53182
rect 185836 53078 185892 53116
rect 186508 53172 186564 53676
rect 187964 53732 188020 55022
rect 187964 53666 188020 53676
rect 182476 52894 182478 52946
rect 182530 52894 182532 52946
rect 182476 52882 182532 52894
rect 186508 52946 186564 53116
rect 186508 52894 186510 52946
rect 186562 52894 186564 52946
rect 186508 52882 186564 52894
rect 181468 52836 181524 52846
rect 181468 52742 181524 52780
rect 183260 52836 183316 52846
rect 183260 52742 183316 52780
rect 185388 52834 185444 52846
rect 185388 52782 185390 52834
rect 185442 52782 185444 52834
rect 173436 51772 173700 51782
rect 173492 51716 173540 51772
rect 173596 51716 173644 51772
rect 173436 51706 173700 51716
rect 173436 50204 173700 50214
rect 173492 50148 173540 50204
rect 173596 50148 173644 50204
rect 173436 50138 173700 50148
rect 173436 48636 173700 48646
rect 173492 48580 173540 48636
rect 173596 48580 173644 48636
rect 173436 48570 173700 48580
rect 173436 47068 173700 47078
rect 173492 47012 173540 47068
rect 173596 47012 173644 47068
rect 173436 47002 173700 47012
rect 173436 45500 173700 45510
rect 173492 45444 173540 45500
rect 173596 45444 173644 45500
rect 173436 45434 173700 45444
rect 173436 43932 173700 43942
rect 173492 43876 173540 43932
rect 173596 43876 173644 43932
rect 173436 43866 173700 43876
rect 173436 42364 173700 42374
rect 173492 42308 173540 42364
rect 173596 42308 173644 42364
rect 173436 42298 173700 42308
rect 173436 40796 173700 40806
rect 173492 40740 173540 40796
rect 173596 40740 173644 40796
rect 173436 40730 173700 40740
rect 173436 39228 173700 39238
rect 173492 39172 173540 39228
rect 173596 39172 173644 39228
rect 173436 39162 173700 39172
rect 173436 37660 173700 37670
rect 173492 37604 173540 37660
rect 173596 37604 173644 37660
rect 173436 37594 173700 37604
rect 173436 36092 173700 36102
rect 173492 36036 173540 36092
rect 173596 36036 173644 36092
rect 173436 36026 173700 36036
rect 173436 34524 173700 34534
rect 173492 34468 173540 34524
rect 173596 34468 173644 34524
rect 173436 34458 173700 34468
rect 173436 32956 173700 32966
rect 173492 32900 173540 32956
rect 173596 32900 173644 32956
rect 173436 32890 173700 32900
rect 173436 31388 173700 31398
rect 173492 31332 173540 31388
rect 173596 31332 173644 31388
rect 173436 31322 173700 31332
rect 173436 29820 173700 29830
rect 173492 29764 173540 29820
rect 173596 29764 173644 29820
rect 173436 29754 173700 29764
rect 173436 28252 173700 28262
rect 173492 28196 173540 28252
rect 173596 28196 173644 28252
rect 173436 28186 173700 28196
rect 173436 26684 173700 26694
rect 173492 26628 173540 26684
rect 173596 26628 173644 26684
rect 173436 26618 173700 26628
rect 173436 25116 173700 25126
rect 173492 25060 173540 25116
rect 173596 25060 173644 25116
rect 173436 25050 173700 25060
rect 173436 23548 173700 23558
rect 173492 23492 173540 23548
rect 173596 23492 173644 23548
rect 173436 23482 173700 23492
rect 173436 21980 173700 21990
rect 173492 21924 173540 21980
rect 173596 21924 173644 21980
rect 173436 21914 173700 21924
rect 178892 21028 178948 21038
rect 173436 20412 173700 20422
rect 173492 20356 173540 20412
rect 173596 20356 173644 20412
rect 173436 20346 173700 20356
rect 173436 18844 173700 18854
rect 173492 18788 173540 18844
rect 173596 18788 173644 18844
rect 173436 18778 173700 18788
rect 173436 17276 173700 17286
rect 173492 17220 173540 17276
rect 173596 17220 173644 17276
rect 173436 17210 173700 17220
rect 173436 15708 173700 15718
rect 173492 15652 173540 15708
rect 173596 15652 173644 15708
rect 173436 15642 173700 15652
rect 173436 14140 173700 14150
rect 173492 14084 173540 14140
rect 173596 14084 173644 14140
rect 173436 14074 173700 14084
rect 173436 12572 173700 12582
rect 173492 12516 173540 12572
rect 173596 12516 173644 12572
rect 173436 12506 173700 12516
rect 171948 11218 172004 11228
rect 111996 11004 112260 11014
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 111996 10938 112260 10948
rect 142716 11004 142980 11014
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142716 10938 142980 10948
rect 173436 11004 173700 11014
rect 173492 10948 173540 11004
rect 173596 10948 173644 11004
rect 173436 10938 173700 10948
rect 127356 10220 127620 10230
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127356 10154 127620 10164
rect 158076 10220 158340 10230
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158076 10154 158340 10164
rect 111996 9436 112260 9446
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 111996 9370 112260 9380
rect 142716 9436 142980 9446
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142716 9370 142980 9380
rect 173436 9436 173700 9446
rect 173492 9380 173540 9436
rect 173596 9380 173644 9436
rect 173436 9370 173700 9380
rect 99932 9202 99988 9212
rect 119196 9156 119252 9166
rect 96636 8652 96900 8662
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96636 8586 96900 8596
rect 111996 7868 112260 7878
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 111996 7802 112260 7812
rect 96636 7084 96900 7094
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96636 7018 96900 7028
rect 111996 6300 112260 6310
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 111996 6234 112260 6244
rect 93548 5908 93604 5918
rect 93548 5236 93604 5852
rect 96636 5516 96900 5526
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96636 5450 96900 5460
rect 93548 5234 93940 5236
rect 93548 5182 93550 5234
rect 93602 5182 93940 5234
rect 93548 5180 93940 5182
rect 93548 5170 93604 5180
rect 91644 4498 91700 4508
rect 93884 4450 93940 5180
rect 111996 4732 112260 4742
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 111996 4666 112260 4676
rect 96236 4564 96292 4574
rect 96292 4508 96516 4564
rect 96236 4470 96292 4508
rect 93884 4398 93886 4450
rect 93938 4398 93940 4450
rect 93884 4386 93940 4398
rect 94220 4450 94276 4462
rect 94220 4398 94222 4450
rect 94274 4398 94276 4450
rect 89628 4340 89684 4350
rect 89068 4228 89124 4238
rect 89068 4134 89124 4172
rect 88732 3614 88734 3666
rect 88786 3614 88788 3666
rect 88732 3556 88788 3614
rect 88732 3490 88788 3500
rect 89404 3556 89460 3566
rect 89404 3462 89460 3500
rect 89628 3442 89684 4284
rect 90972 4340 91028 4350
rect 90972 4246 91028 4284
rect 89628 3390 89630 3442
rect 89682 3390 89684 3442
rect 89628 3378 89684 3390
rect 90748 4116 90804 4126
rect 90748 800 90804 4060
rect 91980 4116 92036 4126
rect 91980 4022 92036 4060
rect 94220 3554 94276 4398
rect 96460 4450 96516 4508
rect 96460 4398 96462 4450
rect 96514 4398 96516 4450
rect 96460 4386 96516 4398
rect 96796 4452 96852 4462
rect 96796 4358 96852 4396
rect 97580 4452 97636 4462
rect 96636 3948 96900 3958
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96636 3882 96900 3892
rect 94220 3502 94222 3554
rect 94274 3502 94276 3554
rect 94220 3490 94276 3502
rect 97580 3554 97636 4396
rect 111804 4226 111860 4238
rect 111804 4174 111806 4226
rect 111858 4174 111860 4226
rect 101612 3668 101668 3678
rect 105420 3668 105476 3678
rect 109116 3668 109172 3678
rect 97580 3502 97582 3554
rect 97634 3502 97636 3554
rect 97580 3490 97636 3502
rect 101500 3666 101668 3668
rect 101500 3614 101614 3666
rect 101666 3614 101668 3666
rect 101500 3612 101668 3614
rect 94780 3332 94836 3342
rect 94332 3330 94836 3332
rect 94332 3278 94782 3330
rect 94834 3278 94836 3330
rect 94332 3276 94836 3278
rect 94332 800 94388 3276
rect 94780 3266 94836 3276
rect 98588 3330 98644 3342
rect 98588 3278 98590 3330
rect 98642 3278 98644 3330
rect 97916 924 98308 980
rect 97916 800 97972 924
rect 8288 0 8400 800
rect 11872 0 11984 800
rect 15456 0 15568 800
rect 19040 0 19152 800
rect 22624 0 22736 800
rect 26208 0 26320 800
rect 29792 0 29904 800
rect 33376 0 33488 800
rect 36960 0 37072 800
rect 40544 0 40656 800
rect 44128 0 44240 800
rect 47712 0 47824 800
rect 51296 0 51408 800
rect 54880 0 54992 800
rect 58464 0 58576 800
rect 62048 0 62160 800
rect 65632 0 65744 800
rect 69216 0 69328 800
rect 72800 0 72912 800
rect 76384 0 76496 800
rect 79968 0 80080 800
rect 83552 0 83664 800
rect 87136 0 87248 800
rect 90720 0 90832 800
rect 94304 0 94416 800
rect 97888 0 98000 800
rect 98252 756 98308 924
rect 98588 756 98644 3278
rect 101500 800 101556 3612
rect 101612 3602 101668 3612
rect 105084 3666 105476 3668
rect 105084 3614 105422 3666
rect 105474 3614 105476 3666
rect 105084 3612 105476 3614
rect 103964 3554 104020 3566
rect 103964 3502 103966 3554
rect 104018 3502 104020 3554
rect 103964 3444 104020 3502
rect 103964 3378 104020 3388
rect 104748 3444 104804 3454
rect 104748 3350 104804 3388
rect 105084 800 105140 3612
rect 105420 3602 105476 3612
rect 108892 3666 109172 3668
rect 108892 3614 109118 3666
rect 109170 3614 109172 3666
rect 108892 3612 109172 3614
rect 107772 3554 107828 3566
rect 107772 3502 107774 3554
rect 107826 3502 107828 3554
rect 107772 3444 107828 3502
rect 107772 3378 107828 3388
rect 108556 3444 108612 3454
rect 108556 3350 108612 3388
rect 108892 980 108948 3612
rect 109116 3602 109172 3612
rect 111468 3556 111524 3566
rect 111468 3462 111524 3500
rect 111804 3556 111860 4174
rect 115388 4226 115444 4238
rect 115388 4174 115390 4226
rect 115442 4174 115444 4226
rect 112700 3668 112756 3678
rect 111804 3490 111860 3500
rect 112364 3666 112756 3668
rect 112364 3614 112702 3666
rect 112754 3614 112756 3666
rect 112364 3612 112756 3614
rect 109340 3444 109396 3454
rect 109340 1092 109396 3388
rect 111996 3164 112260 3174
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 111996 3098 112260 3108
rect 112364 1652 112420 3612
rect 112700 3602 112756 3612
rect 112812 3556 112868 3566
rect 112812 2324 112868 3500
rect 115052 3556 115108 3566
rect 115052 3462 115108 3500
rect 115388 3556 115444 4174
rect 116284 3668 116340 3678
rect 119196 3668 119252 9100
rect 127356 8652 127620 8662
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127356 8586 127620 8596
rect 158076 8652 158340 8662
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158076 8586 158340 8596
rect 142716 7868 142980 7878
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142716 7802 142980 7812
rect 173436 7868 173700 7878
rect 173492 7812 173540 7868
rect 173596 7812 173644 7868
rect 173436 7802 173700 7812
rect 137900 7700 137956 7710
rect 127356 7084 127620 7094
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127356 7018 127620 7028
rect 127356 5516 127620 5526
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127356 5450 127620 5460
rect 122556 5124 122612 5134
rect 122556 4564 122612 5068
rect 122332 4562 122612 4564
rect 122332 4510 122558 4562
rect 122610 4510 122612 4562
rect 122332 4508 122612 4510
rect 119980 3668 120036 3678
rect 115388 3490 115444 3500
rect 115836 3666 116340 3668
rect 115836 3614 116286 3666
rect 116338 3614 116340 3666
rect 115836 3612 116340 3614
rect 112812 2258 112868 2268
rect 109340 1026 109396 1036
rect 112252 1596 112420 1652
rect 108668 924 108948 980
rect 108668 800 108724 924
rect 112252 800 112308 1596
rect 115836 800 115892 3612
rect 116284 3602 116340 3612
rect 118636 3666 119252 3668
rect 118636 3614 119198 3666
rect 119250 3614 119252 3666
rect 118636 3612 119252 3614
rect 118636 3554 118692 3612
rect 119196 3602 119252 3612
rect 119420 3666 120036 3668
rect 119420 3614 119982 3666
rect 120034 3614 120036 3666
rect 119420 3612 120036 3614
rect 118636 3502 118638 3554
rect 118690 3502 118692 3554
rect 118636 3490 118692 3502
rect 119420 800 119476 3612
rect 119980 3602 120036 3612
rect 122332 3554 122388 4508
rect 122556 4498 122612 4508
rect 134316 4900 134372 4910
rect 122332 3502 122334 3554
rect 122386 3502 122388 3554
rect 122332 3490 122388 3502
rect 123900 4116 123956 4126
rect 123116 3444 123172 3454
rect 123564 3444 123620 3454
rect 123004 3442 123620 3444
rect 123004 3390 123118 3442
rect 123170 3390 123566 3442
rect 123618 3390 123620 3442
rect 123004 3388 123620 3390
rect 123004 800 123060 3388
rect 123116 3378 123172 3388
rect 123564 3378 123620 3388
rect 123900 3442 123956 4060
rect 127356 3948 127620 3958
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127356 3882 127620 3892
rect 131516 3780 131572 3790
rect 123900 3390 123902 3442
rect 123954 3390 123956 3442
rect 123900 3378 123956 3390
rect 124348 3556 124404 3566
rect 124348 1540 124404 3500
rect 127708 3556 127764 3566
rect 126924 3444 126980 3454
rect 127372 3444 127428 3454
rect 126924 3442 127428 3444
rect 126924 3390 126926 3442
rect 126978 3390 127374 3442
rect 127426 3390 127428 3442
rect 126924 3388 127428 3390
rect 126924 2212 126980 3388
rect 127372 3378 127428 3388
rect 127708 3442 127764 3500
rect 127708 3390 127710 3442
rect 127762 3390 127764 3442
rect 127708 3378 127764 3390
rect 130732 3444 130788 3454
rect 131180 3444 131236 3454
rect 130732 3442 131236 3444
rect 130732 3390 130734 3442
rect 130786 3390 131182 3442
rect 131234 3390 131236 3442
rect 130732 3388 131236 3390
rect 130732 2212 130788 3388
rect 131180 3378 131236 3388
rect 131516 3442 131572 3724
rect 131516 3390 131518 3442
rect 131570 3390 131572 3442
rect 131516 3378 131572 3390
rect 133756 3444 133812 3454
rect 133980 3444 134036 3454
rect 133756 3442 134036 3444
rect 133756 3390 133758 3442
rect 133810 3390 133982 3442
rect 134034 3390 134036 3442
rect 133756 3388 134036 3390
rect 124348 1474 124404 1484
rect 126588 2156 126980 2212
rect 130172 2156 130788 2212
rect 126588 800 126644 2156
rect 130172 800 130228 2156
rect 133756 800 133812 3388
rect 133980 3378 134036 3388
rect 134316 3442 134372 4844
rect 134316 3390 134318 3442
rect 134370 3390 134372 3442
rect 134316 3378 134372 3390
rect 137340 3444 137396 3454
rect 137564 3444 137620 3454
rect 137340 3442 137620 3444
rect 137340 3390 137342 3442
rect 137394 3390 137566 3442
rect 137618 3390 137620 3442
rect 137340 3388 137620 3390
rect 137340 800 137396 3388
rect 137564 3378 137620 3388
rect 137900 3442 137956 7644
rect 158076 7084 158340 7094
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158076 7018 158340 7028
rect 145068 6916 145124 6926
rect 142716 6300 142980 6310
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142716 6234 142980 6244
rect 141484 6132 141540 6142
rect 137900 3390 137902 3442
rect 137954 3390 137956 3442
rect 137900 3378 137956 3390
rect 140924 3444 140980 3454
rect 141148 3444 141204 3454
rect 140924 3442 141204 3444
rect 140924 3390 140926 3442
rect 140978 3390 141150 3442
rect 141202 3390 141204 3442
rect 140924 3388 141204 3390
rect 140924 800 140980 3388
rect 141148 3378 141204 3388
rect 141484 3442 141540 6076
rect 142716 4732 142980 4742
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142716 4666 142980 4676
rect 141484 3390 141486 3442
rect 141538 3390 141540 3442
rect 141484 3378 141540 3390
rect 144508 3444 144564 3454
rect 144732 3444 144788 3454
rect 144508 3442 144788 3444
rect 144508 3390 144510 3442
rect 144562 3390 144734 3442
rect 144786 3390 144788 3442
rect 144508 3388 144788 3390
rect 142716 3164 142980 3174
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142716 3098 142980 3108
rect 144508 800 144564 3388
rect 144732 3378 144788 3388
rect 145068 3442 145124 6860
rect 148652 6468 148708 6478
rect 145068 3390 145070 3442
rect 145122 3390 145124 3442
rect 145068 3378 145124 3390
rect 148092 3444 148148 3454
rect 148316 3444 148372 3454
rect 148092 3442 148372 3444
rect 148092 3390 148094 3442
rect 148146 3390 148318 3442
rect 148370 3390 148372 3442
rect 148092 3388 148372 3390
rect 148092 800 148148 3388
rect 148316 3378 148372 3388
rect 148652 3442 148708 6412
rect 173436 6300 173700 6310
rect 173492 6244 173540 6300
rect 173596 6244 173644 6300
rect 173436 6234 173700 6244
rect 158076 5516 158340 5526
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158076 5450 158340 5460
rect 173436 4732 173700 4742
rect 173492 4676 173540 4732
rect 173596 4676 173644 4732
rect 173436 4666 173700 4676
rect 173740 4564 173796 4574
rect 152236 4228 152292 4238
rect 148652 3390 148654 3442
rect 148706 3390 148708 3442
rect 148652 3378 148708 3390
rect 151676 3444 151732 3454
rect 151900 3444 151956 3454
rect 151676 3442 151956 3444
rect 151676 3390 151678 3442
rect 151730 3390 151902 3442
rect 151954 3390 151956 3442
rect 151676 3388 151956 3390
rect 151676 800 151732 3388
rect 151900 3378 151956 3388
rect 152236 3442 152292 4172
rect 158076 3948 158340 3958
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158076 3882 158340 3892
rect 170156 3892 170212 3902
rect 152236 3390 152238 3442
rect 152290 3390 152292 3442
rect 152236 3378 152292 3390
rect 155260 3444 155316 3454
rect 155484 3444 155540 3454
rect 155260 3442 155540 3444
rect 155260 3390 155262 3442
rect 155314 3390 155486 3442
rect 155538 3390 155540 3442
rect 155260 3388 155540 3390
rect 155260 800 155316 3388
rect 155484 3378 155540 3388
rect 155820 3444 155876 3454
rect 158844 3444 158900 3454
rect 159068 3444 159124 3454
rect 155820 3442 156324 3444
rect 155820 3390 155822 3442
rect 155874 3390 156324 3442
rect 155820 3388 156324 3390
rect 155820 3378 155876 3388
rect 156268 2436 156324 3388
rect 156268 2370 156324 2380
rect 158844 3442 159124 3444
rect 158844 3390 158846 3442
rect 158898 3390 159070 3442
rect 159122 3390 159124 3442
rect 158844 3388 159124 3390
rect 158844 800 158900 3388
rect 159068 3378 159124 3388
rect 159404 3444 159460 3454
rect 162428 3444 162484 3454
rect 162652 3444 162708 3454
rect 159404 3442 159684 3444
rect 159404 3390 159406 3442
rect 159458 3390 159684 3442
rect 159404 3388 159684 3390
rect 159404 3378 159460 3388
rect 159628 1988 159684 3388
rect 159628 1922 159684 1932
rect 162428 3442 162708 3444
rect 162428 3390 162430 3442
rect 162482 3390 162654 3442
rect 162706 3390 162708 3442
rect 162428 3388 162708 3390
rect 162428 800 162484 3388
rect 162652 3378 162708 3388
rect 166012 3444 166068 3454
rect 166236 3444 166292 3454
rect 166012 3442 166292 3444
rect 166012 3390 166014 3442
rect 166066 3390 166238 3442
rect 166290 3390 166292 3442
rect 166012 3388 166292 3390
rect 162988 3330 163044 3342
rect 162988 3278 162990 3330
rect 163042 3278 163044 3330
rect 162988 2884 163044 3278
rect 162988 2818 163044 2828
rect 166012 800 166068 3388
rect 166236 3378 166292 3388
rect 166572 3444 166628 3454
rect 166572 3350 166628 3388
rect 169596 3444 169652 3454
rect 169820 3444 169876 3454
rect 169596 3442 169876 3444
rect 169596 3390 169598 3442
rect 169650 3390 169822 3442
rect 169874 3390 169876 3442
rect 169596 3388 169876 3390
rect 169596 800 169652 3388
rect 169820 3378 169876 3388
rect 169932 3444 169988 3454
rect 169932 2772 169988 3388
rect 170156 3442 170212 3836
rect 170156 3390 170158 3442
rect 170210 3390 170212 3442
rect 170156 3378 170212 3390
rect 172620 3444 172676 3454
rect 173404 3444 173460 3454
rect 172620 3442 173460 3444
rect 172620 3390 172622 3442
rect 172674 3390 173406 3442
rect 173458 3390 173460 3442
rect 172620 3388 173460 3390
rect 172620 3378 172676 3388
rect 169932 2706 169988 2716
rect 173180 800 173236 3388
rect 173404 3378 173460 3388
rect 173740 3442 173796 4508
rect 173740 3390 173742 3442
rect 173794 3390 173796 3442
rect 173740 3378 173796 3390
rect 176428 3444 176484 3454
rect 176988 3444 177044 3454
rect 176428 3442 177044 3444
rect 176428 3390 176430 3442
rect 176482 3390 176990 3442
rect 177042 3390 177044 3442
rect 176428 3388 177044 3390
rect 176428 3378 176484 3388
rect 173436 3164 173700 3174
rect 173492 3108 173540 3164
rect 173596 3108 173644 3164
rect 173436 3098 173700 3108
rect 176764 800 176820 3388
rect 176988 3378 177044 3388
rect 177324 3330 177380 3342
rect 177324 3278 177326 3330
rect 177378 3278 177380 3330
rect 177324 1204 177380 3278
rect 178892 2548 178948 20972
rect 185388 19348 185444 52782
rect 186172 52836 186228 52846
rect 186172 52276 186228 52780
rect 187180 52836 187236 52846
rect 187180 52742 187236 52780
rect 186172 52182 186228 52220
rect 185388 19282 185444 19292
rect 187292 49588 187348 49598
rect 183372 17668 183428 17678
rect 182252 15988 182308 15998
rect 182252 7588 182308 15932
rect 182252 7522 182308 7532
rect 182364 5908 182420 5918
rect 182364 4562 182420 5852
rect 182700 5124 182756 5134
rect 182364 4510 182366 4562
rect 182418 4510 182420 4562
rect 182364 4498 182420 4510
rect 182476 5122 182756 5124
rect 182476 5070 182702 5122
rect 182754 5070 182756 5122
rect 182476 5068 182756 5070
rect 181580 4226 181636 4238
rect 181580 4174 181582 4226
rect 181634 4174 181636 4226
rect 181580 4116 181636 4174
rect 181580 4050 181636 4060
rect 182252 4226 182308 4238
rect 182252 4174 182254 4226
rect 182306 4174 182308 4226
rect 182252 4116 182308 4174
rect 182252 4050 182308 4060
rect 182028 3780 182084 3790
rect 181020 3668 181076 3678
rect 180236 3444 180292 3454
rect 180684 3444 180740 3454
rect 180236 3442 180740 3444
rect 180236 3390 180238 3442
rect 180290 3390 180686 3442
rect 180738 3390 180740 3442
rect 180236 3388 180740 3390
rect 180236 3378 180292 3388
rect 178892 2482 178948 2492
rect 177324 1138 177380 1148
rect 180348 800 180404 3388
rect 180684 3378 180740 3388
rect 181020 3442 181076 3612
rect 182028 3668 182084 3724
rect 182364 3780 182420 3790
rect 182476 3780 182532 5068
rect 182700 5058 182756 5068
rect 183372 4898 183428 17612
rect 184828 14308 184884 14318
rect 184492 7476 184548 7486
rect 184492 6690 184548 7420
rect 184492 6638 184494 6690
rect 184546 6638 184548 6690
rect 184492 6626 184548 6638
rect 184380 6578 184436 6590
rect 184380 6526 184382 6578
rect 184434 6526 184436 6578
rect 184044 6468 184100 6478
rect 184380 6468 184436 6526
rect 184100 6412 184436 6468
rect 184044 6374 184100 6412
rect 183708 5908 183764 5918
rect 183708 5814 183764 5852
rect 184604 5908 184660 5918
rect 183596 5122 183652 5134
rect 183596 5070 183598 5122
rect 183650 5070 183652 5122
rect 183596 5012 183652 5070
rect 183596 4946 183652 4956
rect 184604 5012 184660 5852
rect 184716 5348 184772 5358
rect 184716 5122 184772 5292
rect 184716 5070 184718 5122
rect 184770 5070 184772 5122
rect 184716 5058 184772 5070
rect 183372 4846 183374 4898
rect 183426 4846 183428 4898
rect 183372 4834 183428 4846
rect 182812 4340 182868 4350
rect 182812 4246 182868 4284
rect 183708 4340 183764 4350
rect 183708 4246 183764 4284
rect 184604 4338 184660 4956
rect 184716 4564 184772 4574
rect 184828 4564 184884 14252
rect 185276 12740 185332 12750
rect 185276 6130 185332 12684
rect 187292 9044 187348 49532
rect 187292 8978 187348 8988
rect 188636 9268 188692 55412
rect 190428 55412 191268 55468
rect 190428 55410 190484 55412
rect 190428 55358 190430 55410
rect 190482 55358 190484 55410
rect 190428 55346 190484 55358
rect 191212 55298 191268 55310
rect 191212 55246 191214 55298
rect 191266 55246 191268 55298
rect 190428 54516 190484 54526
rect 191212 54516 191268 55246
rect 191436 54516 191492 54526
rect 191212 54460 191436 54516
rect 188796 54124 189060 54134
rect 188852 54068 188900 54124
rect 188956 54068 189004 54124
rect 188796 54058 189060 54068
rect 189756 53732 189812 53742
rect 189756 53638 189812 53676
rect 190428 53732 190484 54460
rect 191436 54422 191492 54460
rect 191772 54402 191828 56028
rect 193900 54626 193956 56140
rect 195916 56196 195972 56206
rect 195916 56102 195972 56140
rect 196140 56082 196196 56364
rect 196140 56030 196142 56082
rect 196194 56030 196196 56082
rect 196140 56018 196196 56030
rect 200956 55970 201012 59200
rect 204156 56476 204420 56486
rect 204212 56420 204260 56476
rect 204316 56420 204364 56476
rect 204156 56410 204420 56420
rect 206332 56308 206388 59200
rect 206332 56242 206388 56252
rect 208348 56308 208404 56318
rect 208348 56214 208404 56252
rect 211708 56308 211764 59200
rect 217084 56420 217140 59200
rect 222460 57204 222516 59200
rect 222124 57148 222516 57204
rect 222124 56642 222180 57148
rect 222124 56590 222126 56642
rect 222178 56590 222180 56642
rect 217084 56364 217588 56420
rect 211932 56308 211988 56318
rect 211708 56306 211988 56308
rect 211708 56254 211710 56306
rect 211762 56254 211934 56306
rect 211986 56254 211988 56306
rect 211708 56252 211988 56254
rect 211708 56242 211764 56252
rect 211932 56242 211988 56252
rect 217084 56306 217140 56364
rect 217084 56254 217086 56306
rect 217138 56254 217140 56306
rect 217084 56242 217140 56254
rect 212268 56194 212324 56206
rect 212268 56142 212270 56194
rect 212322 56142 212324 56194
rect 200956 55918 200958 55970
rect 201010 55918 201012 55970
rect 200956 55906 201012 55918
rect 202972 56082 203028 56094
rect 202972 56030 202974 56082
rect 203026 56030 203028 56082
rect 202972 55972 203028 56030
rect 206892 56084 206948 56094
rect 207340 56084 207396 56094
rect 206892 56082 207396 56084
rect 206892 56030 206894 56082
rect 206946 56030 207342 56082
rect 207394 56030 207396 56082
rect 206892 56028 207396 56030
rect 202972 55906 203028 55916
rect 203756 55972 203812 55982
rect 203756 55878 203812 55916
rect 205772 55972 205828 55982
rect 204156 54908 204420 54918
rect 204212 54852 204260 54908
rect 204316 54852 204364 54908
rect 204156 54842 204420 54852
rect 193900 54574 193902 54626
rect 193954 54574 193956 54626
rect 193900 54562 193956 54574
rect 194572 54516 194628 54526
rect 194572 54422 194628 54460
rect 191772 54350 191774 54402
rect 191826 54350 191828 54402
rect 191772 54338 191828 54350
rect 193228 53844 193284 53854
rect 193228 53750 193284 53788
rect 195804 53844 195860 53854
rect 190428 53638 190484 53676
rect 191100 53618 191156 53630
rect 191100 53566 191102 53618
rect 191154 53566 191156 53618
rect 189420 53508 189476 53518
rect 189420 53414 189476 53452
rect 191100 53508 191156 53566
rect 191100 53442 191156 53452
rect 189308 52834 189364 52846
rect 189308 52782 189310 52834
rect 189362 52782 189364 52834
rect 188796 52556 189060 52566
rect 188852 52500 188900 52556
rect 188956 52500 189004 52556
rect 188796 52490 189060 52500
rect 189308 52164 189364 52782
rect 189308 52098 189364 52108
rect 190652 52164 190708 52174
rect 188796 50988 189060 50998
rect 188852 50932 188900 50988
rect 188956 50932 189004 50988
rect 188796 50922 189060 50932
rect 188796 49420 189060 49430
rect 188852 49364 188900 49420
rect 188956 49364 189004 49420
rect 188796 49354 189060 49364
rect 188796 47852 189060 47862
rect 188852 47796 188900 47852
rect 188956 47796 189004 47852
rect 188796 47786 189060 47796
rect 188796 46284 189060 46294
rect 188852 46228 188900 46284
rect 188956 46228 189004 46284
rect 188796 46218 189060 46228
rect 188796 44716 189060 44726
rect 188852 44660 188900 44716
rect 188956 44660 189004 44716
rect 188796 44650 189060 44660
rect 188796 43148 189060 43158
rect 188852 43092 188900 43148
rect 188956 43092 189004 43148
rect 188796 43082 189060 43092
rect 188796 41580 189060 41590
rect 188852 41524 188900 41580
rect 188956 41524 189004 41580
rect 188796 41514 189060 41524
rect 188796 40012 189060 40022
rect 188852 39956 188900 40012
rect 188956 39956 189004 40012
rect 188796 39946 189060 39956
rect 188796 38444 189060 38454
rect 188852 38388 188900 38444
rect 188956 38388 189004 38444
rect 188796 38378 189060 38388
rect 188796 36876 189060 36886
rect 188852 36820 188900 36876
rect 188956 36820 189004 36876
rect 188796 36810 189060 36820
rect 188796 35308 189060 35318
rect 188852 35252 188900 35308
rect 188956 35252 189004 35308
rect 188796 35242 189060 35252
rect 188796 33740 189060 33750
rect 188852 33684 188900 33740
rect 188956 33684 189004 33740
rect 188796 33674 189060 33684
rect 188796 32172 189060 32182
rect 188852 32116 188900 32172
rect 188956 32116 189004 32172
rect 188796 32106 189060 32116
rect 188796 30604 189060 30614
rect 188852 30548 188900 30604
rect 188956 30548 189004 30604
rect 188796 30538 189060 30548
rect 188796 29036 189060 29046
rect 188852 28980 188900 29036
rect 188956 28980 189004 29036
rect 188796 28970 189060 28980
rect 188796 27468 189060 27478
rect 188852 27412 188900 27468
rect 188956 27412 189004 27468
rect 188796 27402 189060 27412
rect 188796 25900 189060 25910
rect 188852 25844 188900 25900
rect 188956 25844 189004 25900
rect 188796 25834 189060 25844
rect 188796 24332 189060 24342
rect 188852 24276 188900 24332
rect 188956 24276 189004 24332
rect 188796 24266 189060 24276
rect 188796 22764 189060 22774
rect 188852 22708 188900 22764
rect 188956 22708 189004 22764
rect 188796 22698 189060 22708
rect 188796 21196 189060 21206
rect 188852 21140 188900 21196
rect 188956 21140 189004 21196
rect 188796 21130 189060 21140
rect 188796 19628 189060 19638
rect 188852 19572 188900 19628
rect 188956 19572 189004 19628
rect 188796 19562 189060 19572
rect 188796 18060 189060 18070
rect 188852 18004 188900 18060
rect 188956 18004 189004 18060
rect 188796 17994 189060 18004
rect 188796 16492 189060 16502
rect 188852 16436 188900 16492
rect 188956 16436 189004 16492
rect 188796 16426 189060 16436
rect 188796 14924 189060 14934
rect 188852 14868 188900 14924
rect 188956 14868 189004 14924
rect 188796 14858 189060 14868
rect 188796 13356 189060 13366
rect 188852 13300 188900 13356
rect 188956 13300 189004 13356
rect 188796 13290 189060 13300
rect 188796 11788 189060 11798
rect 188852 11732 188900 11788
rect 188956 11732 189004 11788
rect 188796 11722 189060 11732
rect 190652 10276 190708 52108
rect 188796 10220 189060 10230
rect 188852 10164 188900 10220
rect 188956 10164 189004 10220
rect 190652 10210 190708 10220
rect 191324 17668 191380 17678
rect 188796 10154 189060 10164
rect 188860 9268 188916 9278
rect 188636 9266 188916 9268
rect 188636 9214 188862 9266
rect 188914 9214 188916 9266
rect 188636 9212 188916 9214
rect 187628 8370 187684 8382
rect 187628 8318 187630 8370
rect 187682 8318 187684 8370
rect 187628 7700 187684 8318
rect 188636 8260 188692 9212
rect 188860 9202 188916 9212
rect 189420 8930 189476 8942
rect 189420 8878 189422 8930
rect 189474 8878 189476 8930
rect 188796 8652 189060 8662
rect 188852 8596 188900 8652
rect 188956 8596 189004 8652
rect 188796 8586 189060 8596
rect 188636 8166 188692 8204
rect 189084 8260 189140 8270
rect 189084 8166 189140 8204
rect 185388 7588 185444 7598
rect 185388 7494 185444 7532
rect 186284 7586 186340 7598
rect 186284 7534 186286 7586
rect 186338 7534 186340 7586
rect 185612 7476 185668 7486
rect 185612 7382 185668 7420
rect 186284 7476 186340 7534
rect 186284 7410 186340 7420
rect 187516 7476 187572 7486
rect 186732 6916 186788 6926
rect 186732 6692 186788 6860
rect 185276 6078 185278 6130
rect 185330 6078 185332 6130
rect 185276 6066 185332 6078
rect 186396 6690 186788 6692
rect 186396 6638 186734 6690
rect 186786 6638 186788 6690
rect 186396 6636 186788 6638
rect 186396 6018 186452 6636
rect 186732 6626 186788 6636
rect 186396 5966 186398 6018
rect 186450 5966 186452 6018
rect 186396 5954 186452 5966
rect 187404 6466 187460 6478
rect 187404 6414 187406 6466
rect 187458 6414 187460 6466
rect 186172 5906 186228 5918
rect 186172 5854 186174 5906
rect 186226 5854 186228 5906
rect 185388 5460 185444 5470
rect 185388 5122 185444 5404
rect 185948 5236 186004 5246
rect 185948 5142 186004 5180
rect 185388 5070 185390 5122
rect 185442 5070 185444 5122
rect 185388 5058 185444 5070
rect 186172 5124 186228 5854
rect 186732 5908 186788 5918
rect 186732 5814 186788 5852
rect 186172 5058 186228 5068
rect 186396 5684 186452 5694
rect 186396 5122 186452 5628
rect 186396 5070 186398 5122
rect 186450 5070 186452 5122
rect 186396 5058 186452 5070
rect 187068 5460 187124 5470
rect 187068 5122 187124 5404
rect 187404 5348 187460 6414
rect 187516 6356 187572 7420
rect 187516 6130 187572 6300
rect 187516 6078 187518 6130
rect 187570 6078 187572 6130
rect 187516 6020 187572 6078
rect 187516 5954 187572 5964
rect 187404 5282 187460 5292
rect 187068 5070 187070 5122
rect 187122 5070 187124 5122
rect 186620 5012 186676 5022
rect 184716 4562 184884 4564
rect 184716 4510 184718 4562
rect 184770 4510 184884 4562
rect 184716 4508 184884 4510
rect 186172 4900 186228 4910
rect 184716 4498 184772 4508
rect 184604 4286 184606 4338
rect 184658 4286 184660 4338
rect 182364 3778 182532 3780
rect 182364 3726 182366 3778
rect 182418 3726 182532 3778
rect 182364 3724 182532 3726
rect 182700 4226 182756 4238
rect 182700 4174 182702 4226
rect 182754 4174 182756 4226
rect 182364 3714 182420 3724
rect 182252 3668 182308 3678
rect 182028 3666 182308 3668
rect 182028 3614 182030 3666
rect 182082 3614 182254 3666
rect 182306 3614 182308 3666
rect 182028 3612 182308 3614
rect 182028 3602 182084 3612
rect 182252 3602 182308 3612
rect 182700 3556 182756 4174
rect 183932 3780 183988 3790
rect 182812 3556 182868 3566
rect 182700 3500 182812 3556
rect 182812 3462 182868 3500
rect 183708 3554 183764 3566
rect 183708 3502 183710 3554
rect 183762 3502 183764 3554
rect 181020 3390 181022 3442
rect 181074 3390 181076 3442
rect 181020 3378 181076 3390
rect 183372 3444 183428 3454
rect 183708 3444 183764 3502
rect 183372 3442 183764 3444
rect 183372 3390 183374 3442
rect 183426 3390 183764 3442
rect 183372 3388 183764 3390
rect 183372 3378 183428 3388
rect 183708 2548 183764 3388
rect 183932 3442 183988 3724
rect 183932 3390 183934 3442
rect 183986 3390 183988 3442
rect 183932 3378 183988 3390
rect 184604 3444 184660 4286
rect 186172 4338 186228 4844
rect 186172 4286 186174 4338
rect 186226 4286 186228 4338
rect 186172 4274 186228 4286
rect 186396 4340 186452 4350
rect 186620 4340 186676 4956
rect 186732 4340 186788 4350
rect 186396 4338 186564 4340
rect 186396 4286 186398 4338
rect 186450 4286 186564 4338
rect 186396 4284 186564 4286
rect 186620 4338 186788 4340
rect 186620 4286 186734 4338
rect 186786 4286 186788 4338
rect 186620 4284 186788 4286
rect 186396 4274 186452 4284
rect 186284 4228 186340 4238
rect 185948 3556 186004 3566
rect 185948 3462 186004 3500
rect 184716 3444 184772 3454
rect 184604 3442 184772 3444
rect 184604 3390 184718 3442
rect 184770 3390 184772 3442
rect 184604 3388 184772 3390
rect 184716 3378 184772 3388
rect 184828 3332 184884 3342
rect 184828 3238 184884 3276
rect 186284 2660 186340 4172
rect 186508 3332 186564 4284
rect 186732 3556 186788 4284
rect 186732 3490 186788 3500
rect 186844 4114 186900 4126
rect 186844 4062 186846 4114
rect 186898 4062 186900 4114
rect 186732 3332 186788 3342
rect 186508 3330 186788 3332
rect 186508 3278 186734 3330
rect 186786 3278 186788 3330
rect 186508 3276 186788 3278
rect 186284 2594 186340 2604
rect 183708 2492 183988 2548
rect 183932 800 183988 2492
rect 186732 2212 186788 3276
rect 186844 2324 186900 4062
rect 186844 2258 186900 2268
rect 187068 2324 187124 5070
rect 187516 5122 187572 5134
rect 187516 5070 187518 5122
rect 187570 5070 187572 5122
rect 187404 4900 187460 4910
rect 187404 4806 187460 4844
rect 187516 3780 187572 5070
rect 187628 5012 187684 7644
rect 187852 8036 187908 8046
rect 187852 7474 187908 7980
rect 188636 7700 188692 7710
rect 189308 7700 189364 7710
rect 188692 7644 188804 7700
rect 188636 7634 188692 7644
rect 188076 7588 188132 7598
rect 188076 7494 188132 7532
rect 188748 7586 188804 7644
rect 188748 7534 188750 7586
rect 188802 7534 188804 7586
rect 188748 7522 188804 7534
rect 189308 7586 189364 7644
rect 189308 7534 189310 7586
rect 189362 7534 189364 7586
rect 189308 7522 189364 7534
rect 187852 7422 187854 7474
rect 187906 7422 187908 7474
rect 187852 7410 187908 7422
rect 189196 7474 189252 7486
rect 189196 7422 189198 7474
rect 189250 7422 189252 7474
rect 188300 7252 188356 7262
rect 187740 6690 187796 6702
rect 187740 6638 187742 6690
rect 187794 6638 187796 6690
rect 187740 6356 187796 6638
rect 188300 6578 188356 7196
rect 188796 7084 189060 7094
rect 188852 7028 188900 7084
rect 188956 7028 189004 7084
rect 188796 7018 189060 7028
rect 188300 6526 188302 6578
rect 188354 6526 188356 6578
rect 187740 6300 188244 6356
rect 187964 6020 188020 6030
rect 187964 5926 188020 5964
rect 187628 4946 187684 4956
rect 187964 4452 188020 4462
rect 187964 4358 188020 4396
rect 187516 3714 187572 3724
rect 187068 2258 187124 2268
rect 187852 3444 187908 3454
rect 188188 3444 188244 6300
rect 188300 4452 188356 6526
rect 188860 5794 188916 5806
rect 188860 5742 188862 5794
rect 188914 5742 188916 5794
rect 188860 5684 188916 5742
rect 189196 5796 189252 7422
rect 189420 6356 189476 8878
rect 191100 8596 191156 8606
rect 189756 8372 189812 8382
rect 189756 8278 189812 8316
rect 190764 8260 190820 8270
rect 190764 8166 190820 8204
rect 190428 8036 190484 8046
rect 190428 7942 190484 7980
rect 191100 7588 191156 8540
rect 191324 7700 191380 17612
rect 193228 15988 193284 15998
rect 192556 11172 192612 11182
rect 192556 8428 192612 11116
rect 192668 9044 192724 9054
rect 192668 8950 192724 8988
rect 193004 9042 193060 9054
rect 193004 8990 193006 9042
rect 193058 8990 193060 9042
rect 192556 8372 192724 8428
rect 191324 7634 191380 7644
rect 191100 7494 191156 7532
rect 192668 7586 192724 8372
rect 192668 7534 192670 7586
rect 192722 7534 192724 7586
rect 192668 7522 192724 7534
rect 190652 7476 190708 7486
rect 190652 7382 190708 7420
rect 192892 7474 192948 7486
rect 192892 7422 192894 7474
rect 192946 7422 192948 7474
rect 191660 7362 191716 7374
rect 191660 7310 191662 7362
rect 191714 7310 191716 7362
rect 189868 7252 189924 7262
rect 189868 7158 189924 7196
rect 190876 6804 190932 6814
rect 190316 6690 190372 6702
rect 190316 6638 190318 6690
rect 190370 6638 190372 6690
rect 190316 6468 190372 6638
rect 190316 6402 190372 6412
rect 190652 6690 190708 6702
rect 190652 6638 190654 6690
rect 190706 6638 190708 6690
rect 189420 6290 189476 6300
rect 189308 5908 189364 5918
rect 189308 5906 189476 5908
rect 189308 5854 189310 5906
rect 189362 5854 189476 5906
rect 189308 5852 189476 5854
rect 189308 5842 189364 5852
rect 189196 5730 189252 5740
rect 188860 5618 188916 5628
rect 188796 5516 189060 5526
rect 188852 5460 188900 5516
rect 188956 5460 189004 5516
rect 188796 5450 189060 5460
rect 188300 4386 188356 4396
rect 188860 5010 188916 5022
rect 188860 4958 188862 5010
rect 188914 4958 188916 5010
rect 188860 4452 188916 4958
rect 189420 4676 189476 5852
rect 190428 5796 190484 5806
rect 190428 5702 190484 5740
rect 190652 5684 190708 6638
rect 190316 5348 190372 5358
rect 189308 4564 189364 4574
rect 189420 4564 189476 4620
rect 189308 4562 189476 4564
rect 189308 4510 189310 4562
rect 189362 4510 189476 4562
rect 189308 4508 189476 4510
rect 189868 5124 189924 5134
rect 189868 4562 189924 5068
rect 190316 5122 190372 5292
rect 190316 5070 190318 5122
rect 190370 5070 190372 5122
rect 190316 5058 190372 5070
rect 190652 5236 190708 5628
rect 190652 5122 190708 5180
rect 190652 5070 190654 5122
rect 190706 5070 190708 5122
rect 190652 5058 190708 5070
rect 189868 4510 189870 4562
rect 189922 4510 189924 4562
rect 189308 4498 189364 4508
rect 189868 4498 189924 4510
rect 190316 4788 190372 4798
rect 188860 4386 188916 4396
rect 189868 4338 189924 4350
rect 189868 4286 189870 4338
rect 189922 4286 189924 4338
rect 188796 3948 189060 3958
rect 188852 3892 188900 3948
rect 188956 3892 189004 3948
rect 188796 3882 189060 3892
rect 189868 3668 189924 4286
rect 189868 3602 189924 3612
rect 188524 3554 188580 3566
rect 188524 3502 188526 3554
rect 188578 3502 188580 3554
rect 188300 3444 188356 3454
rect 188188 3442 188356 3444
rect 188188 3390 188302 3442
rect 188354 3390 188356 3442
rect 188188 3388 188356 3390
rect 187852 2212 187908 3388
rect 188300 3378 188356 3388
rect 188524 3444 188580 3502
rect 188524 3378 188580 3388
rect 190092 3442 190148 3454
rect 190092 3390 190094 3442
rect 190146 3390 190148 3442
rect 190092 3220 190148 3390
rect 190316 3444 190372 4732
rect 190540 4452 190596 4462
rect 190540 4358 190596 4396
rect 190540 3444 190596 3454
rect 190764 3444 190820 3454
rect 190316 3442 190820 3444
rect 190316 3390 190542 3442
rect 190594 3390 190766 3442
rect 190818 3390 190820 3442
rect 190316 3388 190820 3390
rect 190540 3378 190596 3388
rect 190764 3378 190820 3388
rect 190876 3442 190932 6748
rect 190988 6692 191044 6702
rect 190988 6598 191044 6636
rect 191660 6132 191716 7310
rect 192892 6804 192948 7422
rect 192892 6738 192948 6748
rect 191660 6018 191716 6076
rect 192332 6690 192388 6702
rect 192332 6638 192334 6690
rect 192386 6638 192388 6690
rect 191660 5966 191662 6018
rect 191714 5966 191716 6018
rect 191660 5954 191716 5966
rect 191772 6020 191828 6030
rect 191772 5926 191828 5964
rect 191100 5908 191156 5918
rect 191100 5814 191156 5852
rect 192332 5796 192388 6638
rect 191660 5236 191716 5246
rect 190988 5124 191044 5134
rect 190988 5030 191044 5068
rect 191660 4450 191716 5180
rect 192332 5236 192388 5740
rect 192332 5122 192388 5180
rect 192668 6580 192724 6590
rect 192668 5460 192724 6524
rect 192780 6468 192836 6478
rect 192780 6374 192836 6412
rect 192892 6020 192948 6030
rect 192892 5906 192948 5964
rect 192892 5854 192894 5906
rect 192946 5854 192948 5906
rect 192892 5842 192948 5854
rect 192668 5234 192724 5404
rect 192780 5348 192836 5358
rect 193004 5348 193060 8990
rect 193228 6692 193284 15932
rect 195020 11172 195076 11182
rect 193564 9268 193620 9278
rect 193228 6598 193284 6636
rect 193340 7812 193396 7822
rect 192780 5346 193060 5348
rect 192780 5294 192782 5346
rect 192834 5294 193060 5346
rect 192780 5292 193060 5294
rect 193116 6468 193172 6478
rect 192780 5282 192836 5292
rect 193116 5236 193172 6412
rect 192668 5182 192670 5234
rect 192722 5182 192724 5234
rect 192668 5170 192724 5182
rect 193004 5180 193172 5236
rect 193228 5236 193284 5246
rect 193340 5236 193396 7756
rect 193564 6130 193620 9212
rect 193676 9042 193732 9054
rect 193676 8990 193678 9042
rect 193730 8990 193732 9042
rect 193676 7476 193732 8990
rect 193900 7812 193956 7822
rect 193788 7476 193844 7486
rect 193676 7474 193844 7476
rect 193676 7422 193790 7474
rect 193842 7422 193844 7474
rect 193676 7420 193844 7422
rect 193564 6078 193566 6130
rect 193618 6078 193620 6130
rect 193564 6066 193620 6078
rect 193788 5906 193844 7420
rect 193900 6690 193956 7756
rect 193900 6638 193902 6690
rect 193954 6638 193956 6690
rect 193900 6626 193956 6638
rect 193788 5854 193790 5906
rect 193842 5854 193844 5906
rect 193228 5234 193396 5236
rect 193228 5182 193230 5234
rect 193282 5182 193396 5234
rect 193228 5180 193396 5182
rect 193676 5236 193732 5246
rect 192332 5070 192334 5122
rect 192386 5070 192388 5122
rect 192332 5058 192388 5070
rect 191660 4398 191662 4450
rect 191714 4398 191716 4450
rect 191660 4386 191716 4398
rect 192780 4338 192836 4350
rect 192780 4286 192782 4338
rect 192834 4286 192836 4338
rect 191660 4228 191716 4238
rect 191212 3444 191268 3454
rect 190876 3390 190878 3442
rect 190930 3390 190932 3442
rect 190876 3378 190932 3390
rect 191100 3442 191268 3444
rect 191100 3390 191214 3442
rect 191266 3390 191268 3442
rect 191100 3388 191268 3390
rect 191100 3220 191156 3388
rect 191212 3378 191268 3388
rect 191548 3444 191604 3454
rect 191660 3444 191716 4172
rect 192780 4116 192836 4286
rect 192780 4050 192836 4060
rect 191548 3442 191716 3444
rect 191548 3390 191550 3442
rect 191602 3390 191716 3442
rect 191548 3388 191716 3390
rect 191548 3378 191604 3388
rect 190092 3164 191156 3220
rect 186732 2146 186788 2156
rect 187516 2156 187908 2212
rect 187516 800 187572 2156
rect 191100 800 191156 3164
rect 193004 1428 193060 5180
rect 193228 5170 193284 5180
rect 193116 4898 193172 4910
rect 193116 4846 193118 4898
rect 193170 4846 193172 4898
rect 193116 3554 193172 4846
rect 193452 4340 193508 4350
rect 193452 4246 193508 4284
rect 193676 4338 193732 5180
rect 193676 4286 193678 4338
rect 193730 4286 193732 4338
rect 193676 4274 193732 4286
rect 193788 4898 193844 5854
rect 194348 6468 194404 6478
rect 195020 6468 195076 11116
rect 195804 10164 195860 53788
rect 204156 53340 204420 53350
rect 204212 53284 204260 53340
rect 204316 53284 204364 53340
rect 204156 53274 204420 53284
rect 204156 51772 204420 51782
rect 204212 51716 204260 51772
rect 204316 51716 204364 51772
rect 204156 51706 204420 51716
rect 204156 50204 204420 50214
rect 204212 50148 204260 50204
rect 204316 50148 204364 50204
rect 204156 50138 204420 50148
rect 204156 48636 204420 48646
rect 204212 48580 204260 48636
rect 204316 48580 204364 48636
rect 204156 48570 204420 48580
rect 204156 47068 204420 47078
rect 204212 47012 204260 47068
rect 204316 47012 204364 47068
rect 204156 47002 204420 47012
rect 204156 45500 204420 45510
rect 204212 45444 204260 45500
rect 204316 45444 204364 45500
rect 204156 45434 204420 45444
rect 204156 43932 204420 43942
rect 204212 43876 204260 43932
rect 204316 43876 204364 43932
rect 204156 43866 204420 43876
rect 204156 42364 204420 42374
rect 204212 42308 204260 42364
rect 204316 42308 204364 42364
rect 204156 42298 204420 42308
rect 204156 40796 204420 40806
rect 204212 40740 204260 40796
rect 204316 40740 204364 40796
rect 204156 40730 204420 40740
rect 204156 39228 204420 39238
rect 204212 39172 204260 39228
rect 204316 39172 204364 39228
rect 204156 39162 204420 39172
rect 204156 37660 204420 37670
rect 204212 37604 204260 37660
rect 204316 37604 204364 37660
rect 204156 37594 204420 37604
rect 204156 36092 204420 36102
rect 204212 36036 204260 36092
rect 204316 36036 204364 36092
rect 204156 36026 204420 36036
rect 204156 34524 204420 34534
rect 204212 34468 204260 34524
rect 204316 34468 204364 34524
rect 204156 34458 204420 34468
rect 204156 32956 204420 32966
rect 204212 32900 204260 32956
rect 204316 32900 204364 32956
rect 204156 32890 204420 32900
rect 204156 31388 204420 31398
rect 204212 31332 204260 31388
rect 204316 31332 204364 31388
rect 204156 31322 204420 31332
rect 205772 30324 205828 55916
rect 205772 30258 205828 30268
rect 204156 29820 204420 29830
rect 204212 29764 204260 29820
rect 204316 29764 204364 29820
rect 204156 29754 204420 29764
rect 204156 28252 204420 28262
rect 204212 28196 204260 28252
rect 204316 28196 204364 28252
rect 204156 28186 204420 28196
rect 202300 27748 202356 27758
rect 198492 19348 198548 19358
rect 196700 14308 196756 14318
rect 195804 10098 195860 10108
rect 196140 10388 196196 10398
rect 195468 9940 195524 9950
rect 195356 9042 195412 9054
rect 195356 8990 195358 9042
rect 195410 8990 195412 9042
rect 195356 7700 195412 8990
rect 195356 7634 195412 7644
rect 195244 7588 195300 7598
rect 194348 6466 195076 6468
rect 194348 6414 194350 6466
rect 194402 6414 195076 6466
rect 194348 6412 195076 6414
rect 195132 7474 195188 7486
rect 195132 7422 195134 7474
rect 195186 7422 195188 7474
rect 194348 5124 194404 6412
rect 195020 5460 195076 5470
rect 194348 5058 194404 5068
rect 194572 5236 194628 5246
rect 194572 5122 194628 5180
rect 195020 5234 195076 5404
rect 195020 5182 195022 5234
rect 195074 5182 195076 5234
rect 195020 5170 195076 5182
rect 194572 5070 194574 5122
rect 194626 5070 194628 5122
rect 194572 5058 194628 5070
rect 195132 5124 195188 7422
rect 195132 5058 195188 5068
rect 195244 6356 195300 7532
rect 195244 5236 195300 6300
rect 195356 6132 195412 6142
rect 195356 5906 195412 6076
rect 195356 5854 195358 5906
rect 195410 5854 195412 5906
rect 195356 5842 195412 5854
rect 193788 4846 193790 4898
rect 193842 4846 193844 4898
rect 193116 3502 193118 3554
rect 193170 3502 193172 3554
rect 193116 3490 193172 3502
rect 193564 3556 193620 3566
rect 193788 3556 193844 4846
rect 193564 3554 193844 3556
rect 193564 3502 193566 3554
rect 193618 3502 193844 3554
rect 193564 3500 193844 3502
rect 194796 4900 194852 4910
rect 194796 3554 194852 4844
rect 195244 4564 195300 5180
rect 195468 5348 195524 9884
rect 196028 9828 196084 9838
rect 196028 9268 196084 9772
rect 195580 9266 196084 9268
rect 195580 9214 196030 9266
rect 196082 9214 196084 9266
rect 195580 9212 196084 9214
rect 195580 9154 195636 9212
rect 196028 9202 196084 9212
rect 195580 9102 195582 9154
rect 195634 9102 195636 9154
rect 195580 9090 195636 9102
rect 196028 7700 196084 7710
rect 196140 7700 196196 10332
rect 195580 7698 196196 7700
rect 195580 7646 196030 7698
rect 196082 7646 196196 7698
rect 195580 7644 196196 7646
rect 196252 10052 196308 10062
rect 195580 7586 195636 7644
rect 196028 7634 196084 7644
rect 195580 7534 195582 7586
rect 195634 7534 195636 7586
rect 195580 7522 195636 7534
rect 195916 6692 195972 6702
rect 196252 6692 196308 9996
rect 195580 6690 196308 6692
rect 195580 6638 195918 6690
rect 195970 6638 196308 6690
rect 195580 6636 196308 6638
rect 195580 6018 195636 6636
rect 195916 6626 195972 6636
rect 195580 5966 195582 6018
rect 195634 5966 195636 6018
rect 195580 5954 195636 5966
rect 196028 6468 196084 6478
rect 196028 5908 196084 6412
rect 196028 5814 196084 5852
rect 195468 5234 195524 5292
rect 195468 5182 195470 5234
rect 195522 5182 195524 5234
rect 195468 5170 195524 5182
rect 196252 5122 196308 5134
rect 196252 5070 196254 5122
rect 196306 5070 196308 5122
rect 196140 4900 196196 4910
rect 196140 4806 196196 4844
rect 195356 4564 195412 4574
rect 195244 4562 195412 4564
rect 195244 4510 195358 4562
rect 195410 4510 195412 4562
rect 195244 4508 195412 4510
rect 195356 4498 195412 4508
rect 195804 4226 195860 4238
rect 195804 4174 195806 4226
rect 195858 4174 195860 4226
rect 195804 4116 195860 4174
rect 194796 3502 194798 3554
rect 194850 3502 194852 3554
rect 193564 3490 193620 3500
rect 194796 3490 194852 3502
rect 195356 3556 195412 3566
rect 195356 3462 195412 3500
rect 194684 3444 194740 3454
rect 193340 3330 193396 3342
rect 193340 3278 193342 3330
rect 193394 3278 193396 3330
rect 193340 2548 193396 3278
rect 193340 2482 193396 2492
rect 193004 1362 193060 1372
rect 194684 800 194740 3388
rect 195804 1652 195860 4060
rect 195916 3444 195972 3454
rect 195916 3350 195972 3388
rect 196252 3442 196308 5070
rect 196364 4676 196420 4686
rect 196364 4562 196420 4620
rect 196364 4510 196366 4562
rect 196418 4510 196420 4562
rect 196364 4498 196420 4510
rect 196700 4452 196756 14252
rect 197596 9268 197652 9278
rect 196812 6690 196868 6702
rect 196812 6638 196814 6690
rect 196866 6638 196868 6690
rect 196812 5682 196868 6638
rect 197596 6690 197652 9212
rect 198492 9268 198548 19292
rect 199164 10276 199220 10286
rect 199164 9940 199220 10220
rect 199724 10164 199780 10174
rect 199780 10108 199892 10164
rect 199724 10098 199780 10108
rect 199836 10052 199892 10108
rect 199836 9996 200116 10052
rect 199164 9938 199780 9940
rect 199164 9886 199166 9938
rect 199218 9886 199780 9938
rect 199164 9884 199780 9886
rect 199164 9874 199220 9884
rect 199724 9604 199780 9884
rect 198828 9268 198884 9278
rect 198492 9266 198884 9268
rect 198492 9214 198494 9266
rect 198546 9214 198830 9266
rect 198882 9214 198884 9266
rect 198492 9212 198884 9214
rect 198492 9202 198548 9212
rect 198828 8372 198884 9212
rect 199164 9154 199220 9166
rect 199164 9102 199166 9154
rect 199218 9102 199220 9154
rect 198828 8306 198884 8316
rect 199052 8820 199108 8830
rect 199052 8370 199108 8764
rect 199164 8428 199220 9102
rect 199724 9042 199780 9548
rect 199724 8990 199726 9042
rect 199778 8990 199780 9042
rect 199724 8978 199780 8990
rect 199836 9156 199892 9996
rect 200060 9938 200116 9996
rect 200060 9886 200062 9938
rect 200114 9886 200116 9938
rect 200060 9874 200116 9886
rect 200956 9604 201012 9614
rect 201012 9548 201348 9604
rect 200956 9510 201012 9548
rect 201292 9266 201348 9548
rect 201292 9214 201294 9266
rect 201346 9214 201348 9266
rect 201292 9202 201348 9214
rect 202300 9268 202356 27692
rect 204156 26684 204420 26694
rect 204212 26628 204260 26684
rect 204316 26628 204364 26684
rect 204156 26618 204420 26628
rect 204156 25116 204420 25126
rect 204212 25060 204260 25116
rect 204316 25060 204364 25116
rect 204156 25050 204420 25060
rect 204156 23548 204420 23558
rect 204212 23492 204260 23548
rect 204316 23492 204364 23548
rect 204156 23482 204420 23492
rect 204156 21980 204420 21990
rect 204212 21924 204260 21980
rect 204316 21924 204364 21980
rect 204156 21914 204420 21924
rect 204156 20412 204420 20422
rect 204212 20356 204260 20412
rect 204316 20356 204364 20412
rect 204156 20346 204420 20356
rect 204156 18844 204420 18854
rect 204212 18788 204260 18844
rect 204316 18788 204364 18844
rect 204156 18778 204420 18788
rect 206892 17668 206948 56028
rect 207340 56018 207396 56028
rect 209132 55860 209188 55870
rect 206892 17602 206948 17612
rect 207900 21028 207956 21038
rect 204156 17276 204420 17286
rect 204212 17220 204260 17276
rect 204316 17220 204364 17276
rect 204156 17210 204420 17220
rect 204156 15708 204420 15718
rect 204212 15652 204260 15708
rect 204316 15652 204364 15708
rect 204156 15642 204420 15652
rect 204156 14140 204420 14150
rect 204212 14084 204260 14140
rect 204316 14084 204364 14140
rect 204156 14074 204420 14084
rect 203644 12740 203700 12750
rect 202300 9174 202356 9212
rect 203084 9604 203140 9614
rect 203084 9268 203140 9548
rect 203084 9266 203252 9268
rect 203084 9214 203086 9266
rect 203138 9214 203252 9266
rect 203084 9212 203252 9214
rect 203084 9202 203140 9212
rect 200396 9156 200452 9166
rect 199836 9154 200452 9156
rect 199836 9102 200398 9154
rect 200450 9102 200452 9154
rect 199836 9100 200452 9102
rect 203196 9156 203252 9212
rect 203644 9266 203700 12684
rect 204156 12572 204420 12582
rect 204212 12516 204260 12572
rect 204316 12516 204364 12572
rect 204156 12506 204420 12516
rect 204156 11004 204420 11014
rect 204212 10948 204260 11004
rect 204316 10948 204364 11004
rect 204156 10938 204420 10948
rect 204156 9436 204420 9446
rect 204212 9380 204260 9436
rect 204316 9380 204364 9436
rect 204156 9370 204420 9380
rect 203644 9214 203646 9266
rect 203698 9214 203700 9266
rect 203196 9100 203364 9156
rect 199500 8930 199556 8942
rect 199500 8878 199502 8930
rect 199554 8878 199556 8930
rect 199500 8820 199556 8878
rect 199836 8820 199892 9100
rect 200396 9090 200452 9100
rect 201292 9044 201348 9054
rect 200956 8930 201012 8942
rect 200956 8878 200958 8930
rect 201010 8878 201012 8930
rect 199556 8764 199892 8820
rect 200060 8818 200116 8830
rect 200060 8766 200062 8818
rect 200114 8766 200116 8818
rect 199500 8726 199556 8764
rect 200060 8428 200116 8766
rect 199164 8372 199332 8428
rect 199052 8318 199054 8370
rect 199106 8318 199108 8370
rect 199052 8306 199108 8318
rect 198492 7474 198548 7486
rect 198492 7422 198494 7474
rect 198546 7422 198548 7474
rect 198492 7364 198548 7422
rect 199276 7476 199332 8372
rect 199612 8372 199668 8382
rect 200060 8372 200228 8428
rect 199668 8316 200004 8372
rect 199612 8278 199668 8316
rect 199948 8258 200004 8316
rect 199948 8206 199950 8258
rect 200002 8206 200004 8258
rect 199948 8194 200004 8206
rect 200060 8148 200116 8158
rect 200060 8054 200116 8092
rect 199724 8036 199780 8046
rect 199276 7410 199332 7420
rect 199388 7700 199444 7710
rect 198492 7298 198548 7308
rect 199164 7362 199220 7374
rect 199164 7310 199166 7362
rect 199218 7310 199220 7362
rect 197596 6638 197598 6690
rect 197650 6638 197652 6690
rect 197596 6626 197652 6638
rect 197708 7250 197764 7262
rect 197708 7198 197710 7250
rect 197762 7198 197764 7250
rect 197708 6356 197764 7198
rect 196812 5630 196814 5682
rect 196866 5630 196868 5682
rect 196812 5236 196868 5630
rect 196812 5170 196868 5180
rect 197596 6300 197764 6356
rect 197932 6690 197988 6702
rect 197932 6638 197934 6690
rect 197986 6638 197988 6690
rect 197596 5012 197652 6300
rect 197708 6132 197764 6142
rect 197708 6038 197764 6076
rect 197596 4918 197652 4956
rect 197708 5124 197764 5134
rect 197148 4564 197204 4574
rect 197148 4470 197204 4508
rect 197708 4562 197764 5068
rect 197708 4510 197710 4562
rect 197762 4510 197764 4562
rect 197708 4498 197764 4510
rect 197932 5010 197988 6638
rect 198604 6692 198660 6702
rect 199164 6692 199220 7310
rect 199388 6802 199444 7644
rect 199612 7362 199668 7374
rect 199612 7310 199614 7362
rect 199666 7310 199668 7362
rect 199612 7252 199668 7310
rect 199612 7186 199668 7196
rect 199388 6750 199390 6802
rect 199442 6750 199444 6802
rect 199388 6738 199444 6750
rect 198604 6690 199220 6692
rect 198604 6638 198606 6690
rect 198658 6638 199220 6690
rect 198604 6636 199220 6638
rect 198044 5908 198100 5918
rect 198044 5906 198324 5908
rect 198044 5854 198046 5906
rect 198098 5854 198324 5906
rect 198044 5852 198324 5854
rect 198044 5842 198100 5852
rect 197932 4958 197934 5010
rect 197986 4958 197988 5010
rect 197932 4564 197988 4958
rect 197932 4498 197988 4508
rect 198156 5684 198212 5694
rect 198156 4676 198212 5628
rect 196756 4396 196868 4452
rect 196700 4386 196756 4396
rect 196812 3666 196868 4396
rect 197708 4340 197764 4350
rect 197708 4246 197764 4284
rect 196812 3614 196814 3666
rect 196866 3614 196868 3666
rect 196812 3602 196868 3614
rect 198156 3666 198212 4620
rect 198156 3614 198158 3666
rect 198210 3614 198212 3666
rect 198156 3602 198212 3614
rect 196252 3390 196254 3442
rect 196306 3390 196308 3442
rect 196252 3378 196308 3390
rect 197148 3444 197204 3454
rect 197148 3350 197204 3388
rect 197596 3444 197652 3454
rect 198268 3444 198324 5852
rect 198492 3444 198548 3454
rect 198268 3442 198548 3444
rect 198268 3390 198494 3442
rect 198546 3390 198548 3442
rect 198268 3388 198548 3390
rect 197596 2100 197652 3388
rect 198492 3378 198548 3388
rect 198604 2548 198660 6636
rect 199612 6580 199668 6590
rect 199164 6578 199668 6580
rect 199164 6526 199614 6578
rect 199666 6526 199668 6578
rect 199164 6524 199668 6526
rect 199164 6018 199220 6524
rect 199612 6514 199668 6524
rect 199164 5966 199166 6018
rect 199218 5966 199220 6018
rect 199052 5122 199108 5134
rect 199052 5070 199054 5122
rect 199106 5070 199108 5122
rect 199052 3668 199108 5070
rect 199164 5012 199220 5966
rect 199164 4450 199220 4956
rect 199164 4398 199166 4450
rect 199218 4398 199220 4450
rect 199164 4386 199220 4398
rect 199500 6018 199556 6030
rect 199500 5966 199502 6018
rect 199554 5966 199556 6018
rect 199500 4564 199556 5966
rect 199724 6020 199780 7980
rect 199836 7250 199892 7262
rect 199836 7198 199838 7250
rect 199890 7198 199892 7250
rect 199836 6692 199892 7198
rect 200172 7252 200228 8372
rect 200844 8258 200900 8270
rect 200844 8206 200846 8258
rect 200898 8206 200900 8258
rect 200844 8148 200900 8206
rect 200396 7476 200452 7486
rect 200396 7382 200452 7420
rect 200844 7474 200900 8092
rect 200956 8036 201012 8878
rect 200956 7970 201012 7980
rect 201068 8036 201124 8046
rect 201068 8034 201236 8036
rect 201068 7982 201070 8034
rect 201122 7982 201236 8034
rect 201068 7980 201236 7982
rect 201068 7970 201124 7980
rect 201068 7588 201124 7598
rect 200844 7422 200846 7474
rect 200898 7422 200900 7474
rect 200844 7410 200900 7422
rect 200956 7586 201124 7588
rect 200956 7534 201070 7586
rect 201122 7534 201124 7586
rect 200956 7532 201124 7534
rect 200172 7158 200228 7196
rect 199836 6626 199892 6636
rect 199724 5954 199780 5964
rect 200620 5908 200676 5918
rect 200620 5814 200676 5852
rect 199724 5796 199780 5806
rect 199724 5122 199780 5740
rect 200956 5460 201012 7532
rect 201068 7522 201124 7532
rect 201180 6916 201236 7980
rect 201180 6850 201236 6860
rect 201068 6692 201124 6702
rect 201068 6690 201236 6692
rect 201068 6638 201070 6690
rect 201122 6638 201236 6690
rect 201068 6636 201236 6638
rect 201068 6626 201124 6636
rect 200956 5394 201012 5404
rect 199724 5070 199726 5122
rect 199778 5070 199780 5122
rect 199724 5058 199780 5070
rect 200844 5348 200900 5358
rect 199500 4450 199556 4508
rect 199500 4398 199502 4450
rect 199554 4398 199556 4450
rect 199500 4386 199556 4398
rect 200620 4564 200676 4574
rect 200620 4338 200676 4508
rect 200620 4286 200622 4338
rect 200674 4286 200676 4338
rect 200620 4274 200676 4286
rect 199052 3602 199108 3612
rect 198716 3444 198772 3454
rect 198716 2884 198772 3388
rect 198716 2818 198772 2828
rect 198828 3444 198884 3454
rect 199836 3444 199892 3454
rect 198828 3442 199892 3444
rect 198828 3390 198830 3442
rect 198882 3390 199838 3442
rect 199890 3390 199892 3442
rect 198828 3388 199892 3390
rect 198716 2548 198772 2558
rect 198604 2492 198716 2548
rect 198716 2482 198772 2492
rect 198828 2212 198884 3388
rect 199836 3378 199892 3388
rect 200396 3444 200452 3454
rect 200396 3350 200452 3388
rect 200844 3442 200900 5292
rect 201068 5236 201124 5246
rect 201068 5122 201124 5180
rect 201068 5070 201070 5122
rect 201122 5070 201124 5122
rect 201068 5058 201124 5070
rect 201180 4228 201236 6636
rect 201292 5906 201348 8988
rect 201852 8930 201908 8942
rect 203196 8932 203252 8942
rect 201852 8878 201854 8930
rect 201906 8878 201908 8930
rect 201852 8372 201908 8878
rect 203084 8930 203252 8932
rect 203084 8878 203198 8930
rect 203250 8878 203252 8930
rect 203084 8876 203252 8878
rect 203084 8428 203140 8876
rect 203196 8866 203252 8876
rect 203308 8708 203364 9100
rect 203644 9044 203700 9214
rect 203644 8978 203700 8988
rect 205772 9042 205828 9054
rect 205772 8990 205774 9042
rect 205826 8990 205828 9042
rect 201852 8306 201908 8316
rect 202972 8372 203140 8428
rect 203196 8652 203364 8708
rect 203868 8820 203924 8830
rect 202188 8148 202244 8158
rect 202188 8054 202244 8092
rect 202412 8148 202468 8158
rect 202412 7586 202468 8092
rect 202412 7534 202414 7586
rect 202466 7534 202468 7586
rect 202412 7476 202468 7534
rect 202412 7410 202468 7420
rect 202860 7698 202916 7710
rect 202860 7646 202862 7698
rect 202914 7646 202916 7698
rect 202860 7364 202916 7646
rect 202972 7476 203028 8316
rect 203196 8258 203252 8652
rect 203196 8206 203198 8258
rect 203250 8206 203252 8258
rect 203196 8194 203252 8206
rect 203420 8258 203476 8270
rect 203420 8206 203422 8258
rect 203474 8206 203476 8258
rect 202972 7382 203028 7420
rect 203084 8034 203140 8046
rect 203084 7982 203086 8034
rect 203138 7982 203140 8034
rect 201628 6692 201684 6702
rect 201628 6598 201684 6636
rect 202860 6580 202916 7308
rect 203084 6916 203140 7982
rect 203420 8036 203476 8206
rect 203420 7970 203476 7980
rect 202860 6514 202916 6524
rect 202972 6860 203140 6916
rect 203196 7362 203252 7374
rect 203196 7310 203198 7362
rect 203250 7310 203252 7362
rect 202972 6692 203028 6860
rect 201292 5854 201294 5906
rect 201346 5854 201348 5906
rect 201292 5842 201348 5854
rect 201852 5906 201908 5918
rect 201852 5854 201854 5906
rect 201906 5854 201908 5906
rect 201852 5236 201908 5854
rect 202972 5684 203028 6636
rect 203084 6690 203140 6702
rect 203084 6638 203086 6690
rect 203138 6638 203140 6690
rect 203084 6468 203140 6638
rect 203196 6468 203252 7310
rect 203196 6412 203364 6468
rect 203084 6402 203140 6412
rect 203308 6132 203364 6412
rect 203532 6132 203588 6142
rect 203308 6076 203532 6132
rect 203532 6038 203588 6076
rect 202972 5618 203028 5628
rect 203084 5794 203140 5806
rect 203084 5742 203086 5794
rect 203138 5742 203140 5794
rect 201740 5124 201796 5134
rect 201628 5068 201740 5124
rect 201180 4162 201236 4172
rect 201292 4338 201348 4350
rect 201292 4286 201294 4338
rect 201346 4286 201348 4338
rect 201292 4004 201348 4286
rect 201292 3938 201348 3948
rect 200844 3390 200846 3442
rect 200898 3390 200900 3442
rect 200844 2772 200900 3390
rect 200844 2706 200900 2716
rect 201292 3668 201348 3678
rect 201292 3442 201348 3612
rect 201628 3554 201684 5068
rect 201740 5030 201796 5068
rect 201628 3502 201630 3554
rect 201682 3502 201684 3554
rect 201628 3490 201684 3502
rect 201740 4452 201796 4462
rect 201292 3390 201294 3442
rect 201346 3390 201348 3442
rect 197596 2034 197652 2044
rect 198268 2156 198884 2212
rect 195804 1586 195860 1596
rect 198268 800 198324 2156
rect 201292 1316 201348 3390
rect 201740 3442 201796 4396
rect 201852 4338 201908 5180
rect 202972 5348 203028 5358
rect 202524 5124 202580 5134
rect 202412 5122 202580 5124
rect 202412 5070 202526 5122
rect 202578 5070 202580 5122
rect 202412 5068 202580 5070
rect 201964 5010 202020 5022
rect 201964 4958 201966 5010
rect 202018 4958 202020 5010
rect 201964 4452 202020 4958
rect 202076 4452 202132 4462
rect 201964 4396 202076 4452
rect 202076 4386 202132 4396
rect 201852 4286 201854 4338
rect 201906 4286 201908 4338
rect 201852 4274 201908 4286
rect 201740 3390 201742 3442
rect 201794 3390 201796 3442
rect 201740 3378 201796 3390
rect 201852 3892 201908 3902
rect 201292 1250 201348 1260
rect 201852 800 201908 3836
rect 202412 3556 202468 5068
rect 202524 5058 202580 5068
rect 202972 5122 203028 5292
rect 202972 5070 202974 5122
rect 203026 5070 203028 5122
rect 202972 5058 203028 5070
rect 203084 5124 203140 5742
rect 203868 5796 203924 8764
rect 203980 8484 204036 8494
rect 203980 6132 204036 8428
rect 205212 8372 205268 8382
rect 204652 8258 204708 8270
rect 204652 8206 204654 8258
rect 204706 8206 204708 8258
rect 204156 7868 204420 7878
rect 204212 7812 204260 7868
rect 204316 7812 204364 7868
rect 204156 7802 204420 7812
rect 204652 7586 204708 8206
rect 205100 8260 205156 8270
rect 205212 8260 205268 8316
rect 205100 8258 205268 8260
rect 205100 8206 205102 8258
rect 205154 8206 205268 8258
rect 205100 8204 205268 8206
rect 205100 8194 205156 8204
rect 204876 8036 204932 8046
rect 204876 7698 204932 7980
rect 204876 7646 204878 7698
rect 204930 7646 204932 7698
rect 204876 7634 204932 7646
rect 204652 7534 204654 7586
rect 204706 7534 204708 7586
rect 204652 7476 204708 7534
rect 204652 7410 204708 7420
rect 204876 7364 204932 7374
rect 204876 7270 204932 7308
rect 204988 6916 205044 6926
rect 204428 6692 204484 6702
rect 204652 6692 204708 6702
rect 204484 6636 204596 6692
rect 204428 6626 204484 6636
rect 204540 6356 204596 6636
rect 204652 6598 204708 6636
rect 204764 6578 204820 6590
rect 204764 6526 204766 6578
rect 204818 6526 204820 6578
rect 204156 6300 204420 6310
rect 204212 6244 204260 6300
rect 204316 6244 204364 6300
rect 204540 6290 204596 6300
rect 204652 6466 204708 6478
rect 204652 6414 204654 6466
rect 204706 6414 204708 6466
rect 204156 6234 204420 6244
rect 204540 6132 204596 6142
rect 203980 6076 204148 6132
rect 203980 5796 204036 5806
rect 203868 5740 203980 5796
rect 203980 5702 204036 5740
rect 203868 5572 203924 5582
rect 203140 5068 203252 5124
rect 203084 5058 203140 5068
rect 203196 5012 203252 5068
rect 203532 5012 203588 5022
rect 203196 5010 203588 5012
rect 203196 4958 203534 5010
rect 203586 4958 203588 5010
rect 203196 4956 203588 4958
rect 203084 4898 203140 4910
rect 203084 4846 203086 4898
rect 203138 4846 203140 4898
rect 202972 4452 203028 4462
rect 202972 4358 203028 4396
rect 203084 3668 203140 4846
rect 203196 4338 203252 4956
rect 203532 4946 203588 4956
rect 203196 4286 203198 4338
rect 203250 4286 203252 4338
rect 203196 4274 203252 4286
rect 203756 4898 203812 4910
rect 203756 4846 203758 4898
rect 203810 4846 203812 4898
rect 203756 4338 203812 4846
rect 203756 4286 203758 4338
rect 203810 4286 203812 4338
rect 203084 3612 203252 3668
rect 202412 3462 202468 3500
rect 202748 3554 202804 3566
rect 202748 3502 202750 3554
rect 202802 3502 202804 3554
rect 202748 3444 202804 3502
rect 202748 3378 202804 3388
rect 203084 3442 203140 3454
rect 203084 3390 203086 3442
rect 203138 3390 203140 3442
rect 203084 2772 203140 3390
rect 203196 2884 203252 3612
rect 203532 3556 203588 3566
rect 203756 3556 203812 4286
rect 203588 3500 203812 3556
rect 203868 3556 203924 5516
rect 203980 5460 204036 5470
rect 203980 5010 204036 5404
rect 204092 5346 204148 6076
rect 204540 5906 204596 6076
rect 204652 6020 204708 6414
rect 204764 6356 204820 6526
rect 204988 6356 205044 6860
rect 205100 6580 205156 6590
rect 205100 6486 205156 6524
rect 204988 6300 205156 6356
rect 204764 6290 204820 6300
rect 204652 5954 204708 5964
rect 204540 5854 204542 5906
rect 204594 5854 204596 5906
rect 204540 5842 204596 5854
rect 204876 5908 204932 5918
rect 204092 5294 204094 5346
rect 204146 5294 204148 5346
rect 204092 5282 204148 5294
rect 203980 4958 203982 5010
rect 204034 4958 204036 5010
rect 203980 4946 204036 4958
rect 204092 5122 204148 5134
rect 204092 5070 204094 5122
rect 204146 5070 204148 5122
rect 204092 4900 204148 5070
rect 204092 4834 204148 4844
rect 204540 5122 204596 5134
rect 204540 5070 204542 5122
rect 204594 5070 204596 5122
rect 204156 4732 204420 4742
rect 204212 4676 204260 4732
rect 204316 4676 204364 4732
rect 204156 4666 204420 4676
rect 204540 4452 204596 5070
rect 204540 4386 204596 4396
rect 204652 4900 204708 4910
rect 204204 4338 204260 4350
rect 204204 4286 204206 4338
rect 204258 4286 204260 4338
rect 204204 3780 204260 4286
rect 204540 4116 204596 4126
rect 204540 4022 204596 4060
rect 204204 3714 204260 3724
rect 204540 3668 204596 3678
rect 204652 3668 204708 4844
rect 204876 4564 204932 5852
rect 204988 5796 205044 5806
rect 204988 5702 205044 5740
rect 205100 5122 205156 6300
rect 205212 5572 205268 8204
rect 205660 8034 205716 8046
rect 205660 7982 205662 8034
rect 205714 7982 205716 8034
rect 205548 7362 205604 7374
rect 205548 7310 205550 7362
rect 205602 7310 205604 7362
rect 205548 6132 205604 7310
rect 205548 6018 205604 6076
rect 205548 5966 205550 6018
rect 205602 5966 205604 6018
rect 205548 5954 205604 5966
rect 205548 5796 205604 5806
rect 205212 5506 205268 5516
rect 205436 5740 205548 5796
rect 205100 5070 205102 5122
rect 205154 5070 205156 5122
rect 205100 5058 205156 5070
rect 204540 3666 204708 3668
rect 204540 3614 204542 3666
rect 204594 3614 204708 3666
rect 204540 3612 204708 3614
rect 204764 4562 204932 4564
rect 204764 4510 204878 4562
rect 204930 4510 204932 4562
rect 204764 4508 204932 4510
rect 204540 3602 204596 3612
rect 203980 3556 204036 3566
rect 203868 3554 204036 3556
rect 203868 3502 203982 3554
rect 204034 3502 204036 3554
rect 203868 3500 204036 3502
rect 203532 3462 203588 3500
rect 203980 3490 204036 3500
rect 204156 3164 204420 3174
rect 204212 3108 204260 3164
rect 204316 3108 204364 3164
rect 204156 3098 204420 3108
rect 204764 2996 204820 4508
rect 204876 4498 204932 4508
rect 205100 4452 205156 4462
rect 205100 3554 205156 4396
rect 205100 3502 205102 3554
rect 205154 3502 205156 3554
rect 205100 3490 205156 3502
rect 205324 4340 205380 4350
rect 205324 3554 205380 4284
rect 205324 3502 205326 3554
rect 205378 3502 205380 3554
rect 205324 3490 205380 3502
rect 205436 3556 205492 5740
rect 205548 5730 205604 5740
rect 205548 4340 205604 4350
rect 205548 4246 205604 4284
rect 205660 3892 205716 7982
rect 205772 8036 205828 8990
rect 207788 9042 207844 9054
rect 207788 8990 207790 9042
rect 207842 8990 207844 9042
rect 206332 8932 206388 8942
rect 206332 8838 206388 8876
rect 207676 8932 207732 8942
rect 205884 8372 205940 8382
rect 205884 8258 205940 8316
rect 207676 8370 207732 8876
rect 207676 8318 207678 8370
rect 207730 8318 207732 8370
rect 207676 8306 207732 8318
rect 205884 8206 205886 8258
rect 205938 8206 205940 8258
rect 205884 8194 205940 8206
rect 206892 8146 206948 8158
rect 206892 8094 206894 8146
rect 206946 8094 206948 8146
rect 205772 7474 205828 7980
rect 205996 8036 206052 8046
rect 205996 7942 206052 7980
rect 205772 7422 205774 7474
rect 205826 7422 205828 7474
rect 205772 7410 205828 7422
rect 206892 7812 206948 8094
rect 206332 7362 206388 7374
rect 206332 7310 206334 7362
rect 206386 7310 206388 7362
rect 206332 7252 206388 7310
rect 206892 7362 206948 7756
rect 207340 8148 207396 8158
rect 207340 7924 207396 8092
rect 207788 7924 207844 8990
rect 207340 7868 207844 7924
rect 207340 7698 207396 7868
rect 207340 7646 207342 7698
rect 207394 7646 207396 7698
rect 207340 7634 207396 7646
rect 206892 7310 206894 7362
rect 206946 7310 206948 7362
rect 206892 7298 206948 7310
rect 205996 7196 206388 7252
rect 205996 6132 206052 7196
rect 205884 6076 206052 6132
rect 206108 7028 206164 7038
rect 205772 5908 205828 5918
rect 205772 5572 205828 5852
rect 205772 5506 205828 5516
rect 205660 3826 205716 3836
rect 205772 5124 205828 5134
rect 205884 5124 205940 6076
rect 205996 5906 206052 5918
rect 205996 5854 205998 5906
rect 206050 5854 206052 5906
rect 205996 5460 206052 5854
rect 206108 5682 206164 6972
rect 206332 6690 206388 6702
rect 206332 6638 206334 6690
rect 206386 6638 206388 6690
rect 206108 5630 206110 5682
rect 206162 5630 206164 5682
rect 206108 5618 206164 5630
rect 206220 5906 206276 5918
rect 206220 5854 206222 5906
rect 206274 5854 206276 5906
rect 206220 5684 206276 5854
rect 205996 5394 206052 5404
rect 206220 5124 206276 5628
rect 205772 5122 205940 5124
rect 205772 5070 205774 5122
rect 205826 5070 205940 5122
rect 205772 5068 205940 5070
rect 206108 5068 206276 5124
rect 206332 5124 206388 6638
rect 207452 6692 207508 6702
rect 207004 6466 207060 6478
rect 207004 6414 207006 6466
rect 207058 6414 207060 6466
rect 207004 6356 207060 6414
rect 207004 6290 207060 6300
rect 207452 6020 207508 6636
rect 207900 6468 207956 20972
rect 208236 12852 208292 12862
rect 208124 9154 208180 9166
rect 208124 9102 208126 9154
rect 208178 9102 208180 9154
rect 208124 8372 208180 9102
rect 208124 8306 208180 8316
rect 207900 6374 207956 6412
rect 207452 5954 207508 5964
rect 206556 5908 206612 5918
rect 206556 5814 206612 5852
rect 205660 3668 205716 3678
rect 205660 3574 205716 3612
rect 205548 3556 205604 3566
rect 205436 3554 205604 3556
rect 205436 3502 205550 3554
rect 205602 3502 205604 3554
rect 205436 3500 205604 3502
rect 205548 3490 205604 3500
rect 204764 2930 204820 2940
rect 204876 3444 204932 3454
rect 203196 2818 203252 2828
rect 203084 2706 203140 2716
rect 204876 1988 204932 3388
rect 205660 3444 205716 3454
rect 205660 2436 205716 3388
rect 204876 1922 204932 1932
rect 205436 2380 205716 2436
rect 205772 2436 205828 5068
rect 205996 5012 206052 5022
rect 205996 4918 206052 4956
rect 206108 4340 206164 5068
rect 206332 5058 206388 5068
rect 206444 5796 206500 5806
rect 206444 5460 206500 5740
rect 207004 5794 207060 5806
rect 207004 5742 207006 5794
rect 207058 5742 207060 5794
rect 206444 5404 206836 5460
rect 206444 5122 206500 5404
rect 206556 5236 206612 5246
rect 206556 5142 206612 5180
rect 206444 5070 206446 5122
rect 206498 5070 206500 5122
rect 206444 5058 206500 5070
rect 206780 5124 206836 5404
rect 206780 5122 206948 5124
rect 206780 5070 206782 5122
rect 206834 5070 206948 5122
rect 206780 5068 206948 5070
rect 206780 5058 206836 5068
rect 205996 4284 206164 4340
rect 206220 4900 206276 4910
rect 206220 4340 206276 4844
rect 206892 4452 206948 5068
rect 207004 4900 207060 5742
rect 207564 5794 207620 5806
rect 207564 5742 207566 5794
rect 207618 5742 207620 5794
rect 207452 5682 207508 5694
rect 207452 5630 207454 5682
rect 207506 5630 207508 5682
rect 207340 5348 207396 5358
rect 207340 5254 207396 5292
rect 207340 5124 207396 5134
rect 207228 5012 207284 5022
rect 207228 4918 207284 4956
rect 207004 4806 207060 4844
rect 207004 4452 207060 4462
rect 206892 4450 207060 4452
rect 206892 4398 207006 4450
rect 207058 4398 207060 4450
rect 206892 4396 207060 4398
rect 207004 4386 207060 4396
rect 205884 4228 205940 4238
rect 205884 3442 205940 4172
rect 205884 3390 205886 3442
rect 205938 3390 205940 3442
rect 205884 3378 205940 3390
rect 205436 800 205492 2380
rect 205772 2370 205828 2380
rect 205996 1204 206052 4284
rect 206220 4274 206276 4284
rect 206892 4226 206948 4238
rect 206892 4174 206894 4226
rect 206946 4174 206948 4226
rect 206108 3892 206164 3902
rect 206108 3554 206164 3836
rect 206668 3780 206724 3790
rect 206668 3666 206724 3724
rect 206668 3614 206670 3666
rect 206722 3614 206724 3666
rect 206668 3602 206724 3614
rect 206108 3502 206110 3554
rect 206162 3502 206164 3554
rect 206108 3490 206164 3502
rect 205996 1138 206052 1148
rect 206892 1092 206948 4174
rect 207340 3442 207396 5068
rect 207340 3390 207342 3442
rect 207394 3390 207396 3442
rect 207340 3378 207396 3390
rect 207452 5122 207508 5630
rect 207564 5684 207620 5742
rect 207564 5618 207620 5628
rect 208012 5794 208068 5806
rect 208012 5742 208014 5794
rect 208066 5742 208068 5794
rect 208012 5682 208068 5742
rect 208012 5630 208014 5682
rect 208066 5630 208068 5682
rect 208012 5618 208068 5630
rect 208236 5348 208292 12796
rect 209132 8932 209188 55804
rect 212268 55468 212324 56142
rect 217308 56194 217364 56206
rect 217308 56142 217310 56194
rect 217362 56142 217364 56194
rect 212268 55412 212884 55468
rect 210028 30324 210084 30334
rect 209916 9156 209972 9166
rect 209132 8866 209188 8876
rect 209244 8930 209300 8942
rect 209244 8878 209246 8930
rect 209298 8878 209300 8930
rect 209244 8428 209300 8878
rect 209244 8372 209524 8428
rect 209468 8260 209524 8372
rect 209468 7476 209524 8204
rect 209804 8034 209860 8046
rect 209804 7982 209806 8034
rect 209858 7982 209860 8034
rect 209804 7812 209860 7982
rect 209804 7746 209860 7756
rect 209916 7586 209972 9100
rect 210028 8930 210084 30268
rect 211932 11732 211988 11742
rect 211932 10836 211988 11676
rect 211708 10834 211988 10836
rect 211708 10782 211934 10834
rect 211986 10782 211988 10834
rect 211708 10780 211988 10782
rect 210812 9884 211204 9940
rect 210700 9716 210756 9726
rect 210028 8878 210030 8930
rect 210082 8878 210084 8930
rect 210028 8866 210084 8878
rect 210140 9154 210196 9166
rect 210140 9102 210142 9154
rect 210194 9102 210196 9154
rect 210140 8260 210196 9102
rect 210700 9156 210756 9660
rect 210140 8194 210196 8204
rect 210364 8260 210420 8270
rect 209916 7534 209918 7586
rect 209970 7534 209972 7586
rect 209916 7522 209972 7534
rect 210364 8146 210420 8204
rect 210700 8258 210756 9100
rect 210812 9042 210868 9884
rect 211148 9828 211204 9884
rect 211484 9828 211540 9838
rect 211148 9826 211540 9828
rect 211148 9774 211486 9826
rect 211538 9774 211540 9826
rect 211148 9772 211540 9774
rect 211036 9716 211092 9726
rect 211036 9622 211092 9660
rect 210812 8990 210814 9042
rect 210866 8990 210868 9042
rect 210812 8978 210868 8990
rect 210924 9602 210980 9614
rect 210924 9550 210926 9602
rect 210978 9550 210980 9602
rect 210924 8428 210980 9550
rect 211148 9380 211204 9772
rect 211484 9762 211540 9772
rect 211708 9826 211764 10780
rect 211932 10770 211988 10780
rect 211708 9774 211710 9826
rect 211762 9774 211764 9826
rect 211708 9762 211764 9774
rect 212044 9826 212100 9838
rect 212044 9774 212046 9826
rect 212098 9774 212100 9826
rect 211260 9604 211316 9614
rect 211260 9602 211428 9604
rect 211260 9550 211262 9602
rect 211314 9550 211428 9602
rect 211260 9548 211428 9550
rect 211260 9538 211316 9548
rect 210700 8206 210702 8258
rect 210754 8206 210756 8258
rect 210700 8194 210756 8206
rect 210812 8372 210980 8428
rect 211036 9324 211204 9380
rect 211036 8428 211092 9324
rect 211260 9156 211316 9166
rect 211260 9062 211316 9100
rect 211372 8428 211428 9548
rect 211036 8372 211204 8428
rect 210364 8094 210366 8146
rect 210418 8094 210420 8146
rect 209468 7364 209524 7420
rect 210364 7474 210420 8094
rect 210588 8036 210644 8046
rect 210364 7422 210366 7474
rect 210418 7422 210420 7474
rect 210364 7410 210420 7422
rect 210476 8034 210644 8036
rect 210476 7982 210590 8034
rect 210642 7982 210644 8034
rect 210476 7980 210644 7982
rect 209356 7362 209524 7364
rect 209356 7310 209470 7362
rect 209522 7310 209524 7362
rect 209356 7308 209524 7310
rect 208124 5292 208292 5348
rect 208460 5794 208516 5806
rect 208460 5742 208462 5794
rect 208514 5742 208516 5794
rect 207452 5070 207454 5122
rect 207506 5070 207508 5122
rect 207340 2660 207396 2670
rect 207452 2660 207508 5070
rect 208012 5122 208068 5134
rect 208012 5070 208014 5122
rect 208066 5070 208068 5122
rect 208012 4564 208068 5070
rect 207564 3554 207620 3566
rect 207564 3502 207566 3554
rect 207618 3502 207620 3554
rect 207564 3444 207620 3502
rect 207564 3378 207620 3388
rect 208012 3220 208068 4508
rect 208124 4004 208180 5292
rect 208348 5010 208404 5022
rect 208348 4958 208350 5010
rect 208402 4958 208404 5010
rect 208124 3556 208180 3948
rect 208236 4788 208292 4798
rect 208236 4450 208292 4732
rect 208236 4398 208238 4450
rect 208290 4398 208292 4450
rect 208236 3778 208292 4398
rect 208348 4340 208404 4958
rect 208348 4274 208404 4284
rect 208236 3726 208238 3778
rect 208290 3726 208292 3778
rect 208236 3714 208292 3726
rect 208236 3556 208292 3566
rect 208124 3554 208292 3556
rect 208124 3502 208238 3554
rect 208290 3502 208292 3554
rect 208124 3500 208292 3502
rect 208236 3490 208292 3500
rect 208460 3444 208516 5742
rect 208908 5796 208964 5806
rect 209356 5796 209412 7308
rect 209468 7298 209524 7308
rect 209468 7140 209524 7150
rect 209468 6130 209524 7084
rect 210476 6132 210532 7980
rect 210588 7970 210644 7980
rect 209468 6078 209470 6130
rect 209522 6078 209524 6130
rect 209468 5908 209524 6078
rect 209468 5842 209524 5852
rect 210252 6076 210532 6132
rect 210588 6804 210644 6814
rect 208908 5794 209412 5796
rect 208908 5742 208910 5794
rect 208962 5742 209412 5794
rect 208908 5740 209412 5742
rect 209804 5794 209860 5806
rect 209804 5742 209806 5794
rect 209858 5742 209860 5794
rect 208796 5572 208852 5582
rect 208796 5122 208852 5516
rect 208796 5070 208798 5122
rect 208850 5070 208852 5122
rect 208796 5058 208852 5070
rect 208908 4900 208964 5740
rect 209468 5124 209524 5134
rect 209468 5030 209524 5068
rect 208908 4834 208964 4844
rect 209580 5010 209636 5022
rect 209580 4958 209582 5010
rect 209634 4958 209636 5010
rect 209580 4564 209636 4958
rect 209132 4508 209636 4564
rect 208796 4340 208852 4350
rect 209020 4340 209076 4350
rect 208796 4338 209020 4340
rect 208796 4286 208798 4338
rect 208850 4286 209020 4338
rect 208796 4284 209020 4286
rect 208796 4274 208852 4284
rect 208684 3778 208740 3790
rect 208684 3726 208686 3778
rect 208738 3726 208740 3778
rect 208684 3666 208740 3726
rect 208684 3614 208686 3666
rect 208738 3614 208740 3666
rect 208684 3602 208740 3614
rect 208460 3378 208516 3388
rect 209020 3442 209076 4284
rect 209132 3666 209188 4508
rect 209804 4452 209860 5742
rect 209916 5124 209972 5134
rect 209916 5010 209972 5068
rect 210252 5122 210308 6076
rect 210364 5908 210420 5918
rect 210588 5908 210644 6748
rect 210364 5814 210420 5852
rect 210476 5852 210644 5908
rect 210812 5906 210868 8372
rect 211148 8260 211204 8372
rect 211148 8166 211204 8204
rect 211260 8372 211428 8428
rect 211708 9156 211764 9166
rect 210924 8036 210980 8046
rect 211260 8036 211316 8372
rect 211708 8258 211764 9100
rect 212044 8428 212100 9774
rect 212492 9826 212548 9838
rect 212492 9774 212494 9826
rect 212546 9774 212548 9826
rect 212492 9604 212548 9774
rect 212492 9538 212548 9548
rect 212716 9042 212772 9054
rect 212716 8990 212718 9042
rect 212770 8990 212772 9042
rect 211708 8206 211710 8258
rect 211762 8206 211764 8258
rect 211708 8194 211764 8206
rect 211932 8372 212100 8428
rect 212268 8482 212324 8494
rect 212268 8430 212270 8482
rect 212322 8430 212324 8482
rect 212156 8372 212212 8382
rect 211372 8148 211428 8158
rect 211372 8054 211428 8092
rect 210924 8034 211260 8036
rect 210924 7982 210926 8034
rect 210978 7982 211260 8034
rect 210924 7980 211260 7982
rect 210924 7970 210980 7980
rect 211260 7942 211316 7980
rect 211932 8036 211988 8372
rect 211932 7942 211988 7980
rect 212156 8034 212212 8316
rect 212156 7982 212158 8034
rect 212210 7982 212212 8034
rect 212156 7924 212212 7982
rect 212156 7858 212212 7868
rect 211596 7588 211652 7598
rect 211596 7494 211652 7532
rect 210924 7476 210980 7486
rect 210924 7382 210980 7420
rect 210812 5854 210814 5906
rect 210866 5854 210868 5906
rect 210476 5346 210532 5852
rect 210812 5842 210868 5854
rect 211260 5908 211316 5918
rect 211260 5814 211316 5852
rect 211372 5906 211428 5918
rect 211372 5854 211374 5906
rect 211426 5854 211428 5906
rect 210476 5294 210478 5346
rect 210530 5294 210532 5346
rect 210476 5282 210532 5294
rect 210588 5682 210644 5694
rect 210588 5630 210590 5682
rect 210642 5630 210644 5682
rect 210252 5070 210254 5122
rect 210306 5070 210308 5122
rect 210252 5058 210308 5070
rect 209916 4958 209918 5010
rect 209970 4958 209972 5010
rect 209916 4946 209972 4958
rect 209132 3614 209134 3666
rect 209186 3614 209188 3666
rect 209132 3602 209188 3614
rect 209468 4396 209804 4452
rect 209468 3554 209524 4396
rect 209804 4386 209860 4396
rect 210252 4900 210308 4910
rect 210028 4340 210084 4350
rect 210028 4246 210084 4284
rect 210252 4338 210308 4844
rect 210252 4286 210254 4338
rect 210306 4286 210308 4338
rect 210252 4274 210308 4286
rect 210364 4226 210420 4238
rect 210364 4174 210366 4226
rect 210418 4174 210420 4226
rect 209468 3502 209470 3554
rect 209522 3502 209524 3554
rect 209468 3490 209524 3502
rect 210028 3554 210084 3566
rect 210028 3502 210030 3554
rect 210082 3502 210084 3554
rect 209020 3390 209022 3442
rect 209074 3390 209076 3442
rect 209020 3378 209076 3390
rect 209132 3444 209188 3454
rect 209132 3220 209188 3388
rect 209244 3442 209300 3454
rect 209244 3390 209246 3442
rect 209298 3390 209300 3442
rect 209244 3332 209300 3390
rect 209804 3442 209860 3454
rect 209804 3390 209806 3442
rect 209858 3390 209860 3442
rect 209804 3332 209860 3390
rect 210028 3444 210084 3502
rect 210028 3378 210084 3388
rect 209244 3276 209860 3332
rect 208012 3154 208068 3164
rect 209020 3164 209188 3220
rect 207396 2604 207508 2660
rect 207340 2594 207396 2604
rect 206892 1026 206948 1036
rect 209020 800 209076 3164
rect 210364 1540 210420 4174
rect 210588 3780 210644 5630
rect 210700 5572 210756 5582
rect 210700 5122 210756 5516
rect 210700 5070 210702 5122
rect 210754 5070 210756 5122
rect 210700 5058 210756 5070
rect 211036 4898 211092 4910
rect 211036 4846 211038 4898
rect 211090 4846 211092 4898
rect 211036 4788 211092 4846
rect 211036 4722 211092 4732
rect 210812 4452 210868 4462
rect 210812 4358 210868 4396
rect 210476 3724 210644 3780
rect 211148 4340 211204 4350
rect 210476 2212 210532 3724
rect 210588 3556 210644 3566
rect 210588 3462 210644 3500
rect 211148 3442 211204 4284
rect 211372 3666 211428 5854
rect 211596 5794 211652 5806
rect 211596 5742 211598 5794
rect 211650 5742 211652 5794
rect 211596 5460 211652 5742
rect 211596 5394 211652 5404
rect 212268 5122 212324 8430
rect 212380 8260 212436 8270
rect 212380 8166 212436 8204
rect 212716 8036 212772 8990
rect 212828 8148 212884 55412
rect 217308 11844 217364 56142
rect 217532 56082 217588 56364
rect 222124 56306 222180 56590
rect 222124 56254 222126 56306
rect 222178 56254 222180 56306
rect 222124 56242 222180 56254
rect 223020 56642 223076 56654
rect 223020 56590 223022 56642
rect 223074 56590 223076 56642
rect 223020 56306 223076 56590
rect 223020 56254 223022 56306
rect 223074 56254 223076 56306
rect 223020 56242 223076 56254
rect 227836 56420 227892 59200
rect 227836 56364 228340 56420
rect 227836 56306 227892 56364
rect 227836 56254 227838 56306
rect 227890 56254 227892 56306
rect 227836 56242 227892 56254
rect 217532 56030 217534 56082
rect 217586 56030 217588 56082
rect 217532 56018 217588 56030
rect 222684 56194 222740 56206
rect 222684 56142 222686 56194
rect 222738 56142 222740 56194
rect 219516 55692 219780 55702
rect 219572 55636 219620 55692
rect 219676 55636 219724 55692
rect 219516 55626 219780 55636
rect 220668 54628 220724 54638
rect 219516 54124 219780 54134
rect 219572 54068 219620 54124
rect 219676 54068 219724 54124
rect 219516 54058 219780 54068
rect 219516 52556 219780 52566
rect 219572 52500 219620 52556
rect 219676 52500 219724 52556
rect 219516 52490 219780 52500
rect 219516 50988 219780 50998
rect 219572 50932 219620 50988
rect 219676 50932 219724 50988
rect 219516 50922 219780 50932
rect 219516 49420 219780 49430
rect 219572 49364 219620 49420
rect 219676 49364 219724 49420
rect 219516 49354 219780 49364
rect 219516 47852 219780 47862
rect 219572 47796 219620 47852
rect 219676 47796 219724 47852
rect 219516 47786 219780 47796
rect 219516 46284 219780 46294
rect 219572 46228 219620 46284
rect 219676 46228 219724 46284
rect 219516 46218 219780 46228
rect 219516 44716 219780 44726
rect 219572 44660 219620 44716
rect 219676 44660 219724 44716
rect 219516 44650 219780 44660
rect 219516 43148 219780 43158
rect 219572 43092 219620 43148
rect 219676 43092 219724 43148
rect 219516 43082 219780 43092
rect 219516 41580 219780 41590
rect 219572 41524 219620 41580
rect 219676 41524 219724 41580
rect 219516 41514 219780 41524
rect 219516 40012 219780 40022
rect 219572 39956 219620 40012
rect 219676 39956 219724 40012
rect 219516 39946 219780 39956
rect 219516 38444 219780 38454
rect 219572 38388 219620 38444
rect 219676 38388 219724 38444
rect 219516 38378 219780 38388
rect 219516 36876 219780 36886
rect 219572 36820 219620 36876
rect 219676 36820 219724 36876
rect 219516 36810 219780 36820
rect 219516 35308 219780 35318
rect 219572 35252 219620 35308
rect 219676 35252 219724 35308
rect 219516 35242 219780 35252
rect 219516 33740 219780 33750
rect 219572 33684 219620 33740
rect 219676 33684 219724 33740
rect 219516 33674 219780 33684
rect 219516 32172 219780 32182
rect 219572 32116 219620 32172
rect 219676 32116 219724 32172
rect 219516 32106 219780 32116
rect 219516 30604 219780 30614
rect 219572 30548 219620 30604
rect 219676 30548 219724 30604
rect 219516 30538 219780 30548
rect 219516 29036 219780 29046
rect 219572 28980 219620 29036
rect 219676 28980 219724 29036
rect 219516 28970 219780 28980
rect 219516 27468 219780 27478
rect 219572 27412 219620 27468
rect 219676 27412 219724 27468
rect 219516 27402 219780 27412
rect 219516 25900 219780 25910
rect 219572 25844 219620 25900
rect 219676 25844 219724 25900
rect 219516 25834 219780 25844
rect 219516 24332 219780 24342
rect 219572 24276 219620 24332
rect 219676 24276 219724 24332
rect 219516 24266 219780 24276
rect 219516 22764 219780 22774
rect 219572 22708 219620 22764
rect 219676 22708 219724 22764
rect 219516 22698 219780 22708
rect 219516 21196 219780 21206
rect 219572 21140 219620 21196
rect 219676 21140 219724 21196
rect 219516 21130 219780 21140
rect 220668 20188 220724 54572
rect 220668 20132 220948 20188
rect 219516 19628 219780 19638
rect 219572 19572 219620 19628
rect 219676 19572 219724 19628
rect 219516 19562 219780 19572
rect 219516 18060 219780 18070
rect 219572 18004 219620 18060
rect 219676 18004 219724 18060
rect 219516 17994 219780 18004
rect 219516 16492 219780 16502
rect 219572 16436 219620 16492
rect 219676 16436 219724 16492
rect 219516 16426 219780 16436
rect 219516 14924 219780 14934
rect 219572 14868 219620 14924
rect 219676 14868 219724 14924
rect 219516 14858 219780 14868
rect 219516 13356 219780 13366
rect 219572 13300 219620 13356
rect 219676 13300 219724 13356
rect 219516 13290 219780 13300
rect 217308 11778 217364 11788
rect 217420 12964 217476 12974
rect 213612 10388 213668 10398
rect 213388 9156 213444 9166
rect 213388 9042 213444 9100
rect 213388 8990 213390 9042
rect 213442 8990 213444 9042
rect 213388 8978 213444 8990
rect 213612 8428 213668 10332
rect 217420 9940 217476 12908
rect 219516 11788 219780 11798
rect 219572 11732 219620 11788
rect 219676 11732 219724 11788
rect 219516 11722 219780 11732
rect 219516 10220 219780 10230
rect 219572 10164 219620 10220
rect 219676 10164 219724 10220
rect 219516 10154 219780 10164
rect 217196 9938 217476 9940
rect 217196 9886 217422 9938
rect 217474 9886 217476 9938
rect 217196 9884 217476 9886
rect 216748 9604 216804 9614
rect 216748 9266 216804 9548
rect 216748 9214 216750 9266
rect 216802 9214 216804 9266
rect 216748 9202 216804 9214
rect 217196 9154 217252 9884
rect 217420 9874 217476 9884
rect 220556 10052 220612 10062
rect 218316 9828 218372 9838
rect 217196 9102 217198 9154
rect 217250 9102 217252 9154
rect 217196 9090 217252 9102
rect 217532 9604 217588 9614
rect 213836 9044 213892 9054
rect 213836 8950 213892 8988
rect 216524 9044 216580 9054
rect 216524 8950 216580 8988
rect 216972 9042 217028 9054
rect 216972 8990 216974 9042
rect 217026 8990 217028 9042
rect 216412 8932 216468 8942
rect 216188 8930 216468 8932
rect 216188 8878 216414 8930
rect 216466 8878 216468 8930
rect 216188 8876 216468 8878
rect 213388 8372 213668 8428
rect 215740 8596 215796 8606
rect 213388 8260 213444 8372
rect 213388 8166 213444 8204
rect 212828 8054 212884 8092
rect 212716 7970 212772 7980
rect 215740 7698 215796 8540
rect 215740 7646 215742 7698
rect 215794 7646 215796 7698
rect 215740 7634 215796 7646
rect 214060 7588 214116 7598
rect 214060 7474 214116 7532
rect 214732 7588 214788 7598
rect 214060 7422 214062 7474
rect 214114 7422 214116 7474
rect 214060 7410 214116 7422
rect 214508 7474 214564 7486
rect 214508 7422 214510 7474
rect 214562 7422 214564 7474
rect 214508 7364 214564 7422
rect 214508 7298 214564 7308
rect 213836 6916 213892 6926
rect 213836 6690 213892 6860
rect 213836 6638 213838 6690
rect 213890 6638 213892 6690
rect 213836 6626 213892 6638
rect 214620 6916 214676 6926
rect 212268 5070 212270 5122
rect 212322 5070 212324 5122
rect 212268 5058 212324 5070
rect 213612 6468 213668 6478
rect 212380 5010 212436 5022
rect 212380 4958 212382 5010
rect 212434 4958 212436 5010
rect 211820 4898 211876 4910
rect 211820 4846 211822 4898
rect 211874 4846 211876 4898
rect 211372 3614 211374 3666
rect 211426 3614 211428 3666
rect 211372 3602 211428 3614
rect 211596 4452 211652 4462
rect 211596 3554 211652 4396
rect 211596 3502 211598 3554
rect 211650 3502 211652 3554
rect 211596 3490 211652 3502
rect 211148 3390 211150 3442
rect 211202 3390 211204 3442
rect 211148 3378 211204 3390
rect 211372 3444 211428 3454
rect 211372 3350 211428 3388
rect 211820 2324 211876 4846
rect 212380 4564 212436 4958
rect 212604 5010 212660 5022
rect 212604 4958 212606 5010
rect 212658 4958 212660 5010
rect 212380 4498 212436 4508
rect 212492 4788 212548 4798
rect 212492 4562 212548 4732
rect 212492 4510 212494 4562
rect 212546 4510 212548 4562
rect 212492 4498 212548 4510
rect 212604 4562 212660 4958
rect 212604 4510 212606 4562
rect 212658 4510 212660 4562
rect 212604 4498 212660 4510
rect 212828 5010 212884 5022
rect 212828 4958 212830 5010
rect 212882 4958 212884 5010
rect 211932 4452 211988 4462
rect 211932 4338 211988 4396
rect 211932 4286 211934 4338
rect 211986 4286 211988 4338
rect 211932 4274 211988 4286
rect 212268 4338 212324 4350
rect 212268 4286 212270 4338
rect 212322 4286 212324 4338
rect 212044 3556 212100 3566
rect 212044 3462 212100 3500
rect 212268 3556 212324 4286
rect 212828 3780 212884 4958
rect 213612 5012 213668 6412
rect 214620 6132 214676 6860
rect 214284 6130 214676 6132
rect 214284 6078 214622 6130
rect 214674 6078 214676 6130
rect 214284 6076 214676 6078
rect 214284 5122 214340 6076
rect 214620 6066 214676 6076
rect 214284 5070 214286 5122
rect 214338 5070 214340 5122
rect 214284 5058 214340 5070
rect 214732 5236 214788 7532
rect 216188 7474 216244 8876
rect 216412 8866 216468 8876
rect 216972 8372 217028 8990
rect 216972 7812 217028 8316
rect 216972 7746 217028 7756
rect 217308 8484 217364 8494
rect 216188 7422 216190 7474
rect 216242 7422 216244 7474
rect 216188 7410 216244 7422
rect 216412 7476 216468 7486
rect 216412 7382 216468 7420
rect 216524 7474 216580 7486
rect 216524 7422 216526 7474
rect 216578 7422 216580 7474
rect 214956 6020 215012 6030
rect 214956 6018 215236 6020
rect 214956 5966 214958 6018
rect 215010 5966 215236 6018
rect 214956 5964 215236 5966
rect 214956 5954 215012 5964
rect 214732 5124 214788 5180
rect 214732 5122 214900 5124
rect 214732 5070 214734 5122
rect 214786 5070 214900 5122
rect 214732 5068 214900 5070
rect 214732 5058 214788 5068
rect 213612 4946 213668 4956
rect 214508 4898 214564 4910
rect 214508 4846 214510 4898
rect 214562 4846 214564 4898
rect 214508 4676 214564 4846
rect 214508 4610 214564 4620
rect 214844 4338 214900 5068
rect 215180 5122 215236 5964
rect 215292 5908 215348 5918
rect 215292 5234 215348 5852
rect 216188 5906 216244 5918
rect 216188 5854 216190 5906
rect 216242 5854 216244 5906
rect 215852 5796 215908 5806
rect 216188 5796 216244 5854
rect 215908 5740 216244 5796
rect 215852 5702 215908 5740
rect 216188 5572 216244 5740
rect 216412 5906 216468 5918
rect 216412 5854 216414 5906
rect 216466 5854 216468 5906
rect 216412 5796 216468 5854
rect 216412 5730 216468 5740
rect 216524 5794 216580 7422
rect 216748 7362 216804 7374
rect 216748 7310 216750 7362
rect 216802 7310 216804 7362
rect 216748 7028 216804 7310
rect 216748 6962 216804 6972
rect 217196 7364 217252 7374
rect 217196 6804 217252 7308
rect 217196 6690 217252 6748
rect 217196 6638 217198 6690
rect 217250 6638 217252 6690
rect 217196 6626 217252 6638
rect 216524 5742 216526 5794
rect 216578 5742 216580 5794
rect 216524 5730 216580 5742
rect 216636 6018 216692 6030
rect 216636 5966 216638 6018
rect 216690 5966 216692 6018
rect 216188 5516 216580 5572
rect 215964 5348 216020 5358
rect 215292 5182 215294 5234
rect 215346 5182 215348 5234
rect 215292 5170 215348 5182
rect 215628 5236 215684 5246
rect 215180 5070 215182 5122
rect 215234 5070 215236 5122
rect 215180 5012 215236 5070
rect 215628 5122 215684 5180
rect 215628 5070 215630 5122
rect 215682 5070 215684 5122
rect 215628 5058 215684 5070
rect 215180 4946 215236 4956
rect 215404 4900 215460 4910
rect 215404 4898 215572 4900
rect 215404 4846 215406 4898
rect 215458 4846 215572 4898
rect 215404 4844 215572 4846
rect 215404 4834 215460 4844
rect 215292 4676 215348 4686
rect 215292 4562 215348 4620
rect 215292 4510 215294 4562
rect 215346 4510 215348 4562
rect 215292 4498 215348 4510
rect 215404 4564 215460 4574
rect 215516 4564 215572 4844
rect 215964 4788 216020 5292
rect 216188 5124 216244 5134
rect 216188 5030 216244 5068
rect 216076 5012 216132 5022
rect 216076 4918 216132 4956
rect 216300 4900 216356 4910
rect 216300 4806 216356 4844
rect 215964 4732 216132 4788
rect 215964 4564 216020 4574
rect 215516 4508 215964 4564
rect 215404 4470 215460 4508
rect 215964 4470 216020 4508
rect 214844 4286 214846 4338
rect 214898 4286 214900 4338
rect 214844 4274 214900 4286
rect 215516 4340 215572 4350
rect 216076 4340 216132 4732
rect 215516 4338 216132 4340
rect 215516 4286 215518 4338
rect 215570 4286 216132 4338
rect 215516 4284 216132 4286
rect 216524 4340 216580 5516
rect 216636 5012 216692 5966
rect 217084 5796 217140 5806
rect 217084 5702 217140 5740
rect 217308 5234 217364 8428
rect 217532 8258 217588 9548
rect 217756 9268 217812 9278
rect 217756 9154 217812 9212
rect 217756 9102 217758 9154
rect 217810 9102 217812 9154
rect 217756 9090 217812 9102
rect 217980 9044 218036 9054
rect 217980 9042 218148 9044
rect 217980 8990 217982 9042
rect 218034 8990 218148 9042
rect 217980 8988 218148 8990
rect 217980 8978 218036 8988
rect 217868 8820 217924 8830
rect 217868 8818 218036 8820
rect 217868 8766 217870 8818
rect 217922 8766 218036 8818
rect 217868 8764 218036 8766
rect 217868 8754 217924 8764
rect 217532 8206 217534 8258
rect 217586 8206 217588 8258
rect 217532 8194 217588 8206
rect 217756 8148 217812 8158
rect 217756 8054 217812 8092
rect 217756 7476 217812 7486
rect 217756 6802 217812 7420
rect 217756 6750 217758 6802
rect 217810 6750 217812 6802
rect 217756 6738 217812 6750
rect 217644 6468 217700 6478
rect 217644 6374 217700 6412
rect 217868 6466 217924 6478
rect 217868 6414 217870 6466
rect 217922 6414 217924 6466
rect 217868 6132 217924 6414
rect 217868 6066 217924 6076
rect 217308 5182 217310 5234
rect 217362 5182 217364 5234
rect 217308 5170 217364 5182
rect 216636 4946 216692 4956
rect 216860 5122 216916 5134
rect 216860 5070 216862 5122
rect 216914 5070 216916 5122
rect 216860 4900 216916 5070
rect 217756 5124 217812 5134
rect 216748 4452 216804 4462
rect 216748 4358 216804 4396
rect 215516 4274 215572 4284
rect 212828 3714 212884 3724
rect 215404 3778 215460 3790
rect 215404 3726 215406 3778
rect 215458 3726 215460 3778
rect 215404 3666 215460 3726
rect 215404 3614 215406 3666
rect 215458 3614 215460 3666
rect 215404 3602 215460 3614
rect 212268 3490 212324 3500
rect 213052 3554 213108 3566
rect 213052 3502 213054 3554
rect 213106 3502 213108 3554
rect 211820 2258 211876 2268
rect 212604 3442 212660 3454
rect 212604 3390 212606 3442
rect 212658 3390 212660 3442
rect 212604 3220 212660 3390
rect 212828 3444 212884 3454
rect 212828 3350 212884 3388
rect 213052 3220 213108 3502
rect 215852 3330 215908 4284
rect 216524 4246 216580 4284
rect 215852 3278 215854 3330
rect 215906 3278 215908 3330
rect 215852 3266 215908 3278
rect 216188 3778 216244 3790
rect 216188 3726 216190 3778
rect 216242 3726 216244 3778
rect 216188 3556 216244 3726
rect 216860 3780 216916 4844
rect 217084 5012 217140 5022
rect 217084 4562 217140 4956
rect 217420 5010 217476 5022
rect 217420 4958 217422 5010
rect 217474 4958 217476 5010
rect 217084 4510 217086 4562
rect 217138 4510 217140 4562
rect 217084 4498 217140 4510
rect 217308 4564 217364 4574
rect 217308 4470 217364 4508
rect 217420 4226 217476 4958
rect 217756 5010 217812 5068
rect 217980 5122 218036 8764
rect 218092 8148 218148 8988
rect 218204 9042 218260 9054
rect 218204 8990 218206 9042
rect 218258 8990 218260 9042
rect 218204 8372 218260 8990
rect 218204 8306 218260 8316
rect 218092 8082 218148 8092
rect 218204 6804 218260 6814
rect 218204 6690 218260 6748
rect 218204 6638 218206 6690
rect 218258 6638 218260 6690
rect 218204 6626 218260 6638
rect 218316 5346 218372 9772
rect 218428 9716 218484 9726
rect 218428 9154 218484 9660
rect 219548 9716 219604 9726
rect 219100 9268 219156 9278
rect 219100 9174 219156 9212
rect 219548 9266 219604 9660
rect 220220 9324 220500 9380
rect 219548 9214 219550 9266
rect 219602 9214 219604 9266
rect 219548 9202 219604 9214
rect 219996 9268 220052 9278
rect 220220 9268 220276 9324
rect 218428 9102 218430 9154
rect 218482 9102 218484 9154
rect 218428 9090 218484 9102
rect 219996 9154 220052 9212
rect 219996 9102 219998 9154
rect 220050 9102 220052 9154
rect 219996 9090 220052 9102
rect 220108 9212 220276 9268
rect 220444 9266 220500 9324
rect 220444 9214 220446 9266
rect 220498 9214 220500 9266
rect 218764 9044 218820 9054
rect 218764 8950 218820 8988
rect 219516 8652 219780 8662
rect 219572 8596 219620 8652
rect 219676 8596 219724 8652
rect 219516 8586 219780 8596
rect 220108 7924 220164 9212
rect 220444 9202 220500 9214
rect 220332 9156 220388 9166
rect 220220 9042 220276 9054
rect 220220 8990 220222 9042
rect 220274 8990 220276 9042
rect 220220 8148 220276 8990
rect 220332 8372 220388 9100
rect 220556 9044 220612 9996
rect 220892 9940 220948 20132
rect 220668 9938 220948 9940
rect 220668 9886 220894 9938
rect 220946 9886 220948 9938
rect 220668 9884 220948 9886
rect 220668 9154 220724 9884
rect 220892 9874 220948 9884
rect 221788 11284 221844 11294
rect 221788 9716 221844 11228
rect 222684 10388 222740 56142
rect 228060 56194 228116 56206
rect 228060 56142 228062 56194
rect 228114 56142 228116 56194
rect 225932 53956 225988 53966
rect 222684 10322 222740 10332
rect 224252 53844 224308 53854
rect 221788 9650 221844 9660
rect 220668 9102 220670 9154
rect 220722 9102 220724 9154
rect 220668 9090 220724 9102
rect 221228 9268 221284 9278
rect 221228 9154 221284 9212
rect 221228 9102 221230 9154
rect 221282 9102 221284 9154
rect 221228 9090 221284 9102
rect 221900 9268 221956 9278
rect 221900 9154 221956 9212
rect 222348 9268 222404 9278
rect 222348 9174 222404 9212
rect 224252 9268 224308 53788
rect 224252 9202 224308 9212
rect 221900 9102 221902 9154
rect 221954 9102 221956 9154
rect 221900 9090 221956 9102
rect 220444 8988 220612 9044
rect 221452 9044 221508 9054
rect 221452 9042 221620 9044
rect 221452 8990 221454 9042
rect 221506 8990 221620 9042
rect 221452 8988 221620 8990
rect 220444 8484 220500 8988
rect 221452 8978 221508 8988
rect 220556 8820 220612 8830
rect 220556 8818 221284 8820
rect 220556 8766 220558 8818
rect 220610 8766 221284 8818
rect 220556 8764 221284 8766
rect 220556 8754 220612 8764
rect 220444 8428 220948 8484
rect 220332 8316 220724 8372
rect 220668 8260 220724 8316
rect 220780 8260 220836 8270
rect 220668 8258 220836 8260
rect 220668 8206 220782 8258
rect 220834 8206 220836 8258
rect 220668 8204 220836 8206
rect 220780 8194 220836 8204
rect 220220 8082 220276 8092
rect 220220 7924 220276 7934
rect 220108 7868 220220 7924
rect 220220 7858 220276 7868
rect 220780 7812 220836 7822
rect 220668 7700 220724 7710
rect 220556 7644 220668 7700
rect 219516 7084 219780 7094
rect 219572 7028 219620 7084
rect 219676 7028 219724 7084
rect 219516 7018 219780 7028
rect 218316 5294 218318 5346
rect 218370 5294 218372 5346
rect 218316 5282 218372 5294
rect 218540 6466 218596 6478
rect 218540 6414 218542 6466
rect 218594 6414 218596 6466
rect 217980 5070 217982 5122
rect 218034 5070 218036 5122
rect 217980 5058 218036 5070
rect 218540 5236 218596 6414
rect 218540 5122 218596 5180
rect 218540 5070 218542 5122
rect 218594 5070 218596 5122
rect 218540 5058 218596 5070
rect 218876 6468 218932 6478
rect 217756 4958 217758 5010
rect 217810 4958 217812 5010
rect 217756 4946 217812 4958
rect 218876 5010 218932 6412
rect 219100 6466 219156 6478
rect 219100 6414 219102 6466
rect 219154 6414 219156 6466
rect 219100 6132 219156 6414
rect 219100 6066 219156 6076
rect 219548 5794 219604 5806
rect 219548 5742 219550 5794
rect 219602 5742 219604 5794
rect 219548 5684 219604 5742
rect 219324 5628 219604 5684
rect 218988 5124 219044 5134
rect 218988 5030 219044 5068
rect 218876 4958 218878 5010
rect 218930 4958 218932 5010
rect 218876 4946 218932 4958
rect 219100 4898 219156 4910
rect 219100 4846 219102 4898
rect 219154 4846 219156 4898
rect 217532 4452 217588 4462
rect 217532 4358 217588 4396
rect 217980 4340 218036 4350
rect 217980 4246 218036 4284
rect 217420 4174 217422 4226
rect 217474 4174 217476 4226
rect 217420 4162 217476 4174
rect 219100 4228 219156 4846
rect 219324 4788 219380 5628
rect 219516 5516 219780 5526
rect 219572 5460 219620 5516
rect 219676 5460 219724 5516
rect 219516 5450 219780 5460
rect 219772 5122 219828 5134
rect 219772 5070 219774 5122
rect 219826 5070 219828 5122
rect 219772 4788 219828 5070
rect 220556 5122 220612 7644
rect 220668 7634 220724 7644
rect 220780 5346 220836 7756
rect 220780 5294 220782 5346
rect 220834 5294 220836 5346
rect 220780 5282 220836 5294
rect 220892 5346 220948 8428
rect 221228 8260 221284 8764
rect 221116 8204 221284 8260
rect 221340 8482 221396 8494
rect 221340 8430 221342 8482
rect 221394 8430 221396 8482
rect 221004 8148 221060 8158
rect 221004 8054 221060 8092
rect 220892 5294 220894 5346
rect 220946 5294 220948 5346
rect 220892 5282 220948 5294
rect 220556 5070 220558 5122
rect 220610 5070 220612 5122
rect 220556 5058 220612 5070
rect 221116 5122 221172 8204
rect 221228 8034 221284 8046
rect 221228 7982 221230 8034
rect 221282 7982 221284 8034
rect 221228 7924 221284 7982
rect 221228 7858 221284 7868
rect 221116 5070 221118 5122
rect 221170 5070 221172 5122
rect 221116 5058 221172 5070
rect 219100 4162 219156 4172
rect 219212 4732 219828 4788
rect 219996 5010 220052 5022
rect 219996 4958 219998 5010
rect 220050 4958 220052 5010
rect 216860 3714 216916 3724
rect 216636 3556 216692 3566
rect 216188 3554 216692 3556
rect 216188 3502 216638 3554
rect 216690 3502 216692 3554
rect 216188 3500 216692 3502
rect 212604 3164 213108 3220
rect 210476 2146 210532 2156
rect 210364 1474 210420 1484
rect 212604 800 212660 3164
rect 216188 800 216244 3500
rect 216636 3490 216692 3500
rect 216412 3332 216468 3342
rect 216412 3238 216468 3276
rect 219100 2772 219156 2782
rect 219212 2772 219268 4732
rect 219548 4452 219604 4462
rect 219548 4338 219604 4396
rect 219548 4286 219550 4338
rect 219602 4286 219604 4338
rect 219324 4228 219380 4238
rect 219324 4134 219380 4172
rect 219548 4116 219604 4286
rect 219548 4050 219604 4060
rect 219884 4338 219940 4350
rect 219884 4286 219886 4338
rect 219938 4286 219940 4338
rect 219516 3948 219780 3958
rect 219572 3892 219620 3948
rect 219676 3892 219724 3948
rect 219516 3882 219780 3892
rect 219324 3444 219380 3454
rect 219548 3444 219604 3454
rect 219324 3442 219604 3444
rect 219324 3390 219326 3442
rect 219378 3390 219550 3442
rect 219602 3390 219604 3442
rect 219324 3388 219604 3390
rect 219884 3442 219940 4286
rect 219996 4226 220052 4958
rect 220220 5010 220276 5022
rect 220220 4958 220222 5010
rect 220274 4958 220276 5010
rect 220108 4788 220164 4798
rect 220108 4562 220164 4732
rect 220108 4510 220110 4562
rect 220162 4510 220164 4562
rect 220108 4498 220164 4510
rect 219996 4174 219998 4226
rect 220050 4174 220052 4226
rect 219996 4162 220052 4174
rect 220108 4228 220164 4238
rect 220220 4228 220276 4958
rect 220668 4900 220724 4910
rect 220556 4788 220612 4798
rect 220332 4228 220388 4238
rect 220220 4172 220332 4228
rect 219884 3390 219886 3442
rect 219938 3390 219940 3442
rect 219324 3378 219380 3388
rect 219548 3332 219828 3388
rect 219884 3378 219940 3390
rect 219156 2716 219268 2772
rect 219100 2706 219156 2716
rect 219772 800 219828 3332
rect 220108 2772 220164 4172
rect 220332 4162 220388 4172
rect 220220 4004 220276 4014
rect 220220 3554 220276 3948
rect 220556 3668 220612 4732
rect 220668 4452 220724 4844
rect 220668 4358 220724 4396
rect 220780 4340 220836 4350
rect 220780 3778 220836 4284
rect 221340 4338 221396 8430
rect 221452 8372 221508 8382
rect 221452 8258 221508 8316
rect 221452 8206 221454 8258
rect 221506 8206 221508 8258
rect 221452 8194 221508 8206
rect 221564 8148 221620 8988
rect 221564 8082 221620 8092
rect 221676 9042 221732 9054
rect 221676 8990 221678 9042
rect 221730 8990 221732 9042
rect 221676 7924 221732 8990
rect 221676 7858 221732 7868
rect 221788 8818 221844 8830
rect 221788 8766 221790 8818
rect 221842 8766 221844 8818
rect 221788 7700 221844 8766
rect 222012 8372 222068 8382
rect 222012 8278 222068 8316
rect 225932 8372 225988 53900
rect 228060 53844 228116 56142
rect 228284 56082 228340 56364
rect 233212 56308 233268 59200
rect 234876 56476 235140 56486
rect 234932 56420 234980 56476
rect 235036 56420 235084 56476
rect 234876 56410 235140 56420
rect 233548 56308 233604 56318
rect 233212 56252 233548 56308
rect 233548 56214 233604 56252
rect 234220 56308 234276 56318
rect 228284 56030 228286 56082
rect 228338 56030 228340 56082
rect 228284 56018 228340 56030
rect 233996 56194 234052 56206
rect 233996 56142 233998 56194
rect 234050 56142 234052 56194
rect 233996 53956 234052 56142
rect 234220 56082 234276 56252
rect 238588 56308 238644 59200
rect 238812 56308 238868 56318
rect 238588 56306 238868 56308
rect 238588 56254 238590 56306
rect 238642 56254 238814 56306
rect 238866 56254 238868 56306
rect 238588 56252 238868 56254
rect 238588 56242 238644 56252
rect 238812 56242 238868 56252
rect 243964 56308 244020 59200
rect 244188 56308 244244 56318
rect 243964 56306 244244 56308
rect 243964 56254 243966 56306
rect 244018 56254 244190 56306
rect 244242 56254 244244 56306
rect 243964 56252 244244 56254
rect 243964 56242 244020 56252
rect 244188 56242 244244 56252
rect 248780 56308 248836 56318
rect 249340 56308 249396 59200
rect 249564 56308 249620 56318
rect 248780 56306 249620 56308
rect 248780 56254 248782 56306
rect 248834 56254 249566 56306
rect 249618 56254 249620 56306
rect 248780 56252 249620 56254
rect 248780 56242 248836 56252
rect 249564 56242 249620 56252
rect 254716 56308 254772 59200
rect 254716 56306 254996 56308
rect 254716 56254 254718 56306
rect 254770 56254 254996 56306
rect 254716 56252 254996 56254
rect 254716 56242 254772 56252
rect 234220 56030 234222 56082
rect 234274 56030 234276 56082
rect 234220 56018 234276 56030
rect 254940 56082 254996 56252
rect 254940 56030 254942 56082
rect 254994 56030 254996 56082
rect 254940 56018 254996 56030
rect 260092 56306 260148 59200
rect 260092 56254 260094 56306
rect 260146 56254 260148 56306
rect 260092 56084 260148 56254
rect 265468 56308 265524 59200
rect 270844 57090 270900 59200
rect 270844 57038 270846 57090
rect 270898 57038 270900 57090
rect 270844 57026 270900 57038
rect 271516 57090 271572 57102
rect 271516 57038 271518 57090
rect 271570 57038 271572 57090
rect 265596 56476 265860 56486
rect 265652 56420 265700 56476
rect 265756 56420 265804 56476
rect 265596 56410 265860 56420
rect 265468 56306 265748 56308
rect 265468 56254 265470 56306
rect 265522 56254 265748 56306
rect 265468 56252 265748 56254
rect 265468 56242 265524 56252
rect 260092 56018 260148 56028
rect 260764 56084 260820 56094
rect 260764 55990 260820 56028
rect 265692 56082 265748 56252
rect 265692 56030 265694 56082
rect 265746 56030 265748 56082
rect 265692 56018 265748 56030
rect 271516 56306 271572 57038
rect 271516 56254 271518 56306
rect 271570 56254 271572 56306
rect 271516 56084 271572 56254
rect 276220 56308 276276 59200
rect 276220 56306 276500 56308
rect 276220 56254 276222 56306
rect 276274 56254 276500 56306
rect 276220 56252 276500 56254
rect 276220 56242 276276 56252
rect 271516 56018 271572 56028
rect 272188 56084 272244 56094
rect 272188 55990 272244 56028
rect 276444 56082 276500 56252
rect 276444 56030 276446 56082
rect 276498 56030 276500 56082
rect 276444 56018 276500 56030
rect 281596 56084 281652 59200
rect 286860 56308 286916 56318
rect 286972 56308 287028 59200
rect 287308 56308 287364 56318
rect 286860 56306 287364 56308
rect 286860 56254 286862 56306
rect 286914 56254 287310 56306
rect 287362 56254 287364 56306
rect 286860 56252 287364 56254
rect 286860 56242 286916 56252
rect 287308 56242 287364 56252
rect 292348 56308 292404 59200
rect 296316 56476 296580 56486
rect 296372 56420 296420 56476
rect 296476 56420 296524 56476
rect 296316 56410 296580 56420
rect 292572 56308 292628 56318
rect 292348 56306 292628 56308
rect 292348 56254 292350 56306
rect 292402 56254 292574 56306
rect 292626 56254 292628 56306
rect 292348 56252 292628 56254
rect 292348 56242 292404 56252
rect 292572 56242 292628 56252
rect 281596 56018 281652 56028
rect 282716 56084 282772 56094
rect 282716 55990 282772 56028
rect 283612 56084 283668 56094
rect 283612 55990 283668 56028
rect 239260 55970 239316 55982
rect 239260 55918 239262 55970
rect 239314 55918 239316 55970
rect 234876 54908 235140 54918
rect 234932 54852 234980 54908
rect 235036 54852 235084 54908
rect 234876 54842 235140 54852
rect 239260 54628 239316 55918
rect 239260 54562 239316 54572
rect 244748 55970 244804 55982
rect 244748 55918 244750 55970
rect 244802 55918 244804 55970
rect 233996 53890 234052 53900
rect 228060 53778 228116 53788
rect 234876 53340 235140 53350
rect 234932 53284 234980 53340
rect 235036 53284 235084 53340
rect 234876 53274 235140 53284
rect 234876 51772 235140 51782
rect 234932 51716 234980 51772
rect 235036 51716 235084 51772
rect 234876 51706 235140 51716
rect 234876 50204 235140 50214
rect 234932 50148 234980 50204
rect 235036 50148 235084 50204
rect 234876 50138 235140 50148
rect 234876 48636 235140 48646
rect 234932 48580 234980 48636
rect 235036 48580 235084 48636
rect 234876 48570 235140 48580
rect 234876 47068 235140 47078
rect 234932 47012 234980 47068
rect 235036 47012 235084 47068
rect 234876 47002 235140 47012
rect 234876 45500 235140 45510
rect 234932 45444 234980 45500
rect 235036 45444 235084 45500
rect 234876 45434 235140 45444
rect 234876 43932 235140 43942
rect 234932 43876 234980 43932
rect 235036 43876 235084 43932
rect 234876 43866 235140 43876
rect 234876 42364 235140 42374
rect 234932 42308 234980 42364
rect 235036 42308 235084 42364
rect 234876 42298 235140 42308
rect 234876 40796 235140 40806
rect 234932 40740 234980 40796
rect 235036 40740 235084 40796
rect 234876 40730 235140 40740
rect 234876 39228 235140 39238
rect 234932 39172 234980 39228
rect 235036 39172 235084 39228
rect 234876 39162 235140 39172
rect 234876 37660 235140 37670
rect 234932 37604 234980 37660
rect 235036 37604 235084 37660
rect 234876 37594 235140 37604
rect 234876 36092 235140 36102
rect 234932 36036 234980 36092
rect 235036 36036 235084 36092
rect 234876 36026 235140 36036
rect 234876 34524 235140 34534
rect 234932 34468 234980 34524
rect 235036 34468 235084 34524
rect 234876 34458 235140 34468
rect 234876 32956 235140 32966
rect 234932 32900 234980 32956
rect 235036 32900 235084 32956
rect 234876 32890 235140 32900
rect 234876 31388 235140 31398
rect 234932 31332 234980 31388
rect 235036 31332 235084 31388
rect 234876 31322 235140 31332
rect 234876 29820 235140 29830
rect 234932 29764 234980 29820
rect 235036 29764 235084 29820
rect 234876 29754 235140 29764
rect 234876 28252 235140 28262
rect 234932 28196 234980 28252
rect 235036 28196 235084 28252
rect 234876 28186 235140 28196
rect 234876 26684 235140 26694
rect 234932 26628 234980 26684
rect 235036 26628 235084 26684
rect 234876 26618 235140 26628
rect 234876 25116 235140 25126
rect 234932 25060 234980 25116
rect 235036 25060 235084 25116
rect 234876 25050 235140 25060
rect 234876 23548 235140 23558
rect 234932 23492 234980 23548
rect 235036 23492 235084 23548
rect 234876 23482 235140 23492
rect 234876 21980 235140 21990
rect 234932 21924 234980 21980
rect 235036 21924 235084 21980
rect 234876 21914 235140 21924
rect 234876 20412 235140 20422
rect 234932 20356 234980 20412
rect 235036 20356 235084 20412
rect 234876 20346 235140 20356
rect 234876 18844 235140 18854
rect 234932 18788 234980 18844
rect 235036 18788 235084 18844
rect 234876 18778 235140 18788
rect 234876 17276 235140 17286
rect 234932 17220 234980 17276
rect 235036 17220 235084 17276
rect 234876 17210 235140 17220
rect 234876 15708 235140 15718
rect 234932 15652 234980 15708
rect 235036 15652 235084 15708
rect 234876 15642 235140 15652
rect 234876 14140 235140 14150
rect 234932 14084 234980 14140
rect 235036 14084 235084 14140
rect 234876 14074 235140 14084
rect 234876 12572 235140 12582
rect 234932 12516 234980 12572
rect 235036 12516 235084 12572
rect 234876 12506 235140 12516
rect 244748 11284 244804 55918
rect 250124 55970 250180 55982
rect 250124 55918 250126 55970
rect 250178 55918 250180 55970
rect 250124 12964 250180 55918
rect 256060 55970 256116 55982
rect 256060 55918 256062 55970
rect 256114 55918 256116 55970
rect 250236 55692 250500 55702
rect 250292 55636 250340 55692
rect 250396 55636 250444 55692
rect 250236 55626 250500 55636
rect 250236 54124 250500 54134
rect 250292 54068 250340 54124
rect 250396 54068 250444 54124
rect 250236 54058 250500 54068
rect 250236 52556 250500 52566
rect 250292 52500 250340 52556
rect 250396 52500 250444 52556
rect 250236 52490 250500 52500
rect 250236 50988 250500 50998
rect 250292 50932 250340 50988
rect 250396 50932 250444 50988
rect 250236 50922 250500 50932
rect 250236 49420 250500 49430
rect 250292 49364 250340 49420
rect 250396 49364 250444 49420
rect 250236 49354 250500 49364
rect 250236 47852 250500 47862
rect 250292 47796 250340 47852
rect 250396 47796 250444 47852
rect 250236 47786 250500 47796
rect 250236 46284 250500 46294
rect 250292 46228 250340 46284
rect 250396 46228 250444 46284
rect 250236 46218 250500 46228
rect 250236 44716 250500 44726
rect 250292 44660 250340 44716
rect 250396 44660 250444 44716
rect 250236 44650 250500 44660
rect 250236 43148 250500 43158
rect 250292 43092 250340 43148
rect 250396 43092 250444 43148
rect 250236 43082 250500 43092
rect 250236 41580 250500 41590
rect 250292 41524 250340 41580
rect 250396 41524 250444 41580
rect 250236 41514 250500 41524
rect 250236 40012 250500 40022
rect 250292 39956 250340 40012
rect 250396 39956 250444 40012
rect 250236 39946 250500 39956
rect 250236 38444 250500 38454
rect 250292 38388 250340 38444
rect 250396 38388 250444 38444
rect 250236 38378 250500 38388
rect 250236 36876 250500 36886
rect 250292 36820 250340 36876
rect 250396 36820 250444 36876
rect 250236 36810 250500 36820
rect 250236 35308 250500 35318
rect 250292 35252 250340 35308
rect 250396 35252 250444 35308
rect 250236 35242 250500 35252
rect 250236 33740 250500 33750
rect 250292 33684 250340 33740
rect 250396 33684 250444 33740
rect 250236 33674 250500 33684
rect 250236 32172 250500 32182
rect 250292 32116 250340 32172
rect 250396 32116 250444 32172
rect 250236 32106 250500 32116
rect 250236 30604 250500 30614
rect 250292 30548 250340 30604
rect 250396 30548 250444 30604
rect 250236 30538 250500 30548
rect 250236 29036 250500 29046
rect 250292 28980 250340 29036
rect 250396 28980 250444 29036
rect 250236 28970 250500 28980
rect 250236 27468 250500 27478
rect 250292 27412 250340 27468
rect 250396 27412 250444 27468
rect 250236 27402 250500 27412
rect 250236 25900 250500 25910
rect 250292 25844 250340 25900
rect 250396 25844 250444 25900
rect 250236 25834 250500 25844
rect 250236 24332 250500 24342
rect 250292 24276 250340 24332
rect 250396 24276 250444 24332
rect 250236 24266 250500 24276
rect 250236 22764 250500 22774
rect 250292 22708 250340 22764
rect 250396 22708 250444 22764
rect 250236 22698 250500 22708
rect 250236 21196 250500 21206
rect 250292 21140 250340 21196
rect 250396 21140 250444 21196
rect 250236 21130 250500 21140
rect 250236 19628 250500 19638
rect 250292 19572 250340 19628
rect 250396 19572 250444 19628
rect 250236 19562 250500 19572
rect 250236 18060 250500 18070
rect 250292 18004 250340 18060
rect 250396 18004 250444 18060
rect 250236 17994 250500 18004
rect 250236 16492 250500 16502
rect 250292 16436 250340 16492
rect 250396 16436 250444 16492
rect 250236 16426 250500 16436
rect 250236 14924 250500 14934
rect 250292 14868 250340 14924
rect 250396 14868 250444 14924
rect 250236 14858 250500 14868
rect 256060 14308 256116 55918
rect 256060 14242 256116 14252
rect 261772 55970 261828 55982
rect 261772 55918 261774 55970
rect 261826 55918 261828 55970
rect 250236 13356 250500 13366
rect 250292 13300 250340 13356
rect 250396 13300 250444 13356
rect 250236 13290 250500 13300
rect 250124 12898 250180 12908
rect 250236 11788 250500 11798
rect 250292 11732 250340 11788
rect 250396 11732 250444 11788
rect 250236 11722 250500 11732
rect 244748 11218 244804 11228
rect 261772 11172 261828 55918
rect 264572 55972 264628 55982
rect 264572 15988 264628 55916
rect 266364 55972 266420 55982
rect 266364 55878 266420 55916
rect 273196 55970 273252 55982
rect 273196 55918 273198 55970
rect 273250 55918 273252 55970
rect 265596 54908 265860 54918
rect 265652 54852 265700 54908
rect 265756 54852 265804 54908
rect 265596 54842 265860 54852
rect 265596 53340 265860 53350
rect 265652 53284 265700 53340
rect 265756 53284 265804 53340
rect 265596 53274 265860 53284
rect 265596 51772 265860 51782
rect 265652 51716 265700 51772
rect 265756 51716 265804 51772
rect 265596 51706 265860 51716
rect 265596 50204 265860 50214
rect 265652 50148 265700 50204
rect 265756 50148 265804 50204
rect 265596 50138 265860 50148
rect 265596 48636 265860 48646
rect 265652 48580 265700 48636
rect 265756 48580 265804 48636
rect 265596 48570 265860 48580
rect 265596 47068 265860 47078
rect 265652 47012 265700 47068
rect 265756 47012 265804 47068
rect 265596 47002 265860 47012
rect 265596 45500 265860 45510
rect 265652 45444 265700 45500
rect 265756 45444 265804 45500
rect 265596 45434 265860 45444
rect 265596 43932 265860 43942
rect 265652 43876 265700 43932
rect 265756 43876 265804 43932
rect 265596 43866 265860 43876
rect 265596 42364 265860 42374
rect 265652 42308 265700 42364
rect 265756 42308 265804 42364
rect 265596 42298 265860 42308
rect 265596 40796 265860 40806
rect 265652 40740 265700 40796
rect 265756 40740 265804 40796
rect 265596 40730 265860 40740
rect 265596 39228 265860 39238
rect 265652 39172 265700 39228
rect 265756 39172 265804 39228
rect 265596 39162 265860 39172
rect 265596 37660 265860 37670
rect 265652 37604 265700 37660
rect 265756 37604 265804 37660
rect 265596 37594 265860 37604
rect 265596 36092 265860 36102
rect 265652 36036 265700 36092
rect 265756 36036 265804 36092
rect 265596 36026 265860 36036
rect 265596 34524 265860 34534
rect 265652 34468 265700 34524
rect 265756 34468 265804 34524
rect 265596 34458 265860 34468
rect 265596 32956 265860 32966
rect 265652 32900 265700 32956
rect 265756 32900 265804 32956
rect 265596 32890 265860 32900
rect 265596 31388 265860 31398
rect 265652 31332 265700 31388
rect 265756 31332 265804 31388
rect 265596 31322 265860 31332
rect 265596 29820 265860 29830
rect 265652 29764 265700 29820
rect 265756 29764 265804 29820
rect 265596 29754 265860 29764
rect 265596 28252 265860 28262
rect 265652 28196 265700 28252
rect 265756 28196 265804 28252
rect 265596 28186 265860 28196
rect 265596 26684 265860 26694
rect 265652 26628 265700 26684
rect 265756 26628 265804 26684
rect 265596 26618 265860 26628
rect 265596 25116 265860 25126
rect 265652 25060 265700 25116
rect 265756 25060 265804 25116
rect 265596 25050 265860 25060
rect 265596 23548 265860 23558
rect 265652 23492 265700 23548
rect 265756 23492 265804 23548
rect 265596 23482 265860 23492
rect 265596 21980 265860 21990
rect 265652 21924 265700 21980
rect 265756 21924 265804 21980
rect 265596 21914 265860 21924
rect 265596 20412 265860 20422
rect 265652 20356 265700 20412
rect 265756 20356 265804 20412
rect 265596 20346 265860 20356
rect 265596 18844 265860 18854
rect 265652 18788 265700 18844
rect 265756 18788 265804 18844
rect 265596 18778 265860 18788
rect 265596 17276 265860 17286
rect 265652 17220 265700 17276
rect 265756 17220 265804 17276
rect 265596 17210 265860 17220
rect 264572 15922 264628 15932
rect 265596 15708 265860 15718
rect 265652 15652 265700 15708
rect 265756 15652 265804 15708
rect 265596 15642 265860 15652
rect 265596 14140 265860 14150
rect 265652 14084 265700 14140
rect 265756 14084 265804 14140
rect 265596 14074 265860 14084
rect 273196 12852 273252 55918
rect 277228 55972 277284 55982
rect 277228 55878 277284 55916
rect 279692 55972 279748 55982
rect 273196 12786 273252 12796
rect 279692 12740 279748 55916
rect 281820 55972 281876 55982
rect 281820 55878 281876 55916
rect 288092 55858 288148 55870
rect 288092 55806 288094 55858
rect 288146 55806 288148 55858
rect 280956 55692 281220 55702
rect 281012 55636 281060 55692
rect 281116 55636 281164 55692
rect 280956 55626 281220 55636
rect 280956 54124 281220 54134
rect 281012 54068 281060 54124
rect 281116 54068 281164 54124
rect 280956 54058 281220 54068
rect 280956 52556 281220 52566
rect 281012 52500 281060 52556
rect 281116 52500 281164 52556
rect 280956 52490 281220 52500
rect 280956 50988 281220 50998
rect 281012 50932 281060 50988
rect 281116 50932 281164 50988
rect 280956 50922 281220 50932
rect 280956 49420 281220 49430
rect 281012 49364 281060 49420
rect 281116 49364 281164 49420
rect 280956 49354 281220 49364
rect 280956 47852 281220 47862
rect 281012 47796 281060 47852
rect 281116 47796 281164 47852
rect 280956 47786 281220 47796
rect 280956 46284 281220 46294
rect 281012 46228 281060 46284
rect 281116 46228 281164 46284
rect 280956 46218 281220 46228
rect 280956 44716 281220 44726
rect 281012 44660 281060 44716
rect 281116 44660 281164 44716
rect 280956 44650 281220 44660
rect 280956 43148 281220 43158
rect 281012 43092 281060 43148
rect 281116 43092 281164 43148
rect 280956 43082 281220 43092
rect 280956 41580 281220 41590
rect 281012 41524 281060 41580
rect 281116 41524 281164 41580
rect 280956 41514 281220 41524
rect 280956 40012 281220 40022
rect 281012 39956 281060 40012
rect 281116 39956 281164 40012
rect 280956 39946 281220 39956
rect 280956 38444 281220 38454
rect 281012 38388 281060 38444
rect 281116 38388 281164 38444
rect 280956 38378 281220 38388
rect 280956 36876 281220 36886
rect 281012 36820 281060 36876
rect 281116 36820 281164 36876
rect 280956 36810 281220 36820
rect 280956 35308 281220 35318
rect 281012 35252 281060 35308
rect 281116 35252 281164 35308
rect 280956 35242 281220 35252
rect 280956 33740 281220 33750
rect 281012 33684 281060 33740
rect 281116 33684 281164 33740
rect 280956 33674 281220 33684
rect 280956 32172 281220 32182
rect 281012 32116 281060 32172
rect 281116 32116 281164 32172
rect 280956 32106 281220 32116
rect 280956 30604 281220 30614
rect 281012 30548 281060 30604
rect 281116 30548 281164 30604
rect 280956 30538 281220 30548
rect 280956 29036 281220 29046
rect 281012 28980 281060 29036
rect 281116 28980 281164 29036
rect 280956 28970 281220 28980
rect 288092 27748 288148 55806
rect 288092 27682 288148 27692
rect 293356 55858 293412 55870
rect 293356 55806 293358 55858
rect 293410 55806 293412 55858
rect 280956 27468 281220 27478
rect 281012 27412 281060 27468
rect 281116 27412 281164 27468
rect 280956 27402 281220 27412
rect 280956 25900 281220 25910
rect 281012 25844 281060 25900
rect 281116 25844 281164 25900
rect 280956 25834 281220 25844
rect 280956 24332 281220 24342
rect 281012 24276 281060 24332
rect 281116 24276 281164 24332
rect 280956 24266 281220 24276
rect 280956 22764 281220 22774
rect 281012 22708 281060 22764
rect 281116 22708 281164 22764
rect 280956 22698 281220 22708
rect 280956 21196 281220 21206
rect 281012 21140 281060 21196
rect 281116 21140 281164 21196
rect 280956 21130 281220 21140
rect 293356 21028 293412 55806
rect 296316 54908 296580 54918
rect 296372 54852 296420 54908
rect 296476 54852 296524 54908
rect 296316 54842 296580 54852
rect 296316 53340 296580 53350
rect 296372 53284 296420 53340
rect 296476 53284 296524 53340
rect 296316 53274 296580 53284
rect 296316 51772 296580 51782
rect 296372 51716 296420 51772
rect 296476 51716 296524 51772
rect 296316 51706 296580 51716
rect 296316 50204 296580 50214
rect 296372 50148 296420 50204
rect 296476 50148 296524 50204
rect 296316 50138 296580 50148
rect 296316 48636 296580 48646
rect 296372 48580 296420 48636
rect 296476 48580 296524 48636
rect 296316 48570 296580 48580
rect 296316 47068 296580 47078
rect 296372 47012 296420 47068
rect 296476 47012 296524 47068
rect 296316 47002 296580 47012
rect 296316 45500 296580 45510
rect 296372 45444 296420 45500
rect 296476 45444 296524 45500
rect 296316 45434 296580 45444
rect 296316 43932 296580 43942
rect 296372 43876 296420 43932
rect 296476 43876 296524 43932
rect 296316 43866 296580 43876
rect 296316 42364 296580 42374
rect 296372 42308 296420 42364
rect 296476 42308 296524 42364
rect 296316 42298 296580 42308
rect 296316 40796 296580 40806
rect 296372 40740 296420 40796
rect 296476 40740 296524 40796
rect 296316 40730 296580 40740
rect 296316 39228 296580 39238
rect 296372 39172 296420 39228
rect 296476 39172 296524 39228
rect 296316 39162 296580 39172
rect 296316 37660 296580 37670
rect 296372 37604 296420 37660
rect 296476 37604 296524 37660
rect 296316 37594 296580 37604
rect 296316 36092 296580 36102
rect 296372 36036 296420 36092
rect 296476 36036 296524 36092
rect 296316 36026 296580 36036
rect 296316 34524 296580 34534
rect 296372 34468 296420 34524
rect 296476 34468 296524 34524
rect 296316 34458 296580 34468
rect 296316 32956 296580 32966
rect 296372 32900 296420 32956
rect 296476 32900 296524 32956
rect 296316 32890 296580 32900
rect 296316 31388 296580 31398
rect 296372 31332 296420 31388
rect 296476 31332 296524 31388
rect 296316 31322 296580 31332
rect 296316 29820 296580 29830
rect 296372 29764 296420 29820
rect 296476 29764 296524 29820
rect 296316 29754 296580 29764
rect 296316 28252 296580 28262
rect 296372 28196 296420 28252
rect 296476 28196 296524 28252
rect 296316 28186 296580 28196
rect 296316 26684 296580 26694
rect 296372 26628 296420 26684
rect 296476 26628 296524 26684
rect 296316 26618 296580 26628
rect 296316 25116 296580 25126
rect 296372 25060 296420 25116
rect 296476 25060 296524 25116
rect 296316 25050 296580 25060
rect 296316 23548 296580 23558
rect 296372 23492 296420 23548
rect 296476 23492 296524 23548
rect 296316 23482 296580 23492
rect 296316 21980 296580 21990
rect 296372 21924 296420 21980
rect 296476 21924 296524 21980
rect 296316 21914 296580 21924
rect 293356 20962 293412 20972
rect 296316 20412 296580 20422
rect 296372 20356 296420 20412
rect 296476 20356 296524 20412
rect 296316 20346 296580 20356
rect 280956 19628 281220 19638
rect 281012 19572 281060 19628
rect 281116 19572 281164 19628
rect 280956 19562 281220 19572
rect 296316 18844 296580 18854
rect 296372 18788 296420 18844
rect 296476 18788 296524 18844
rect 296316 18778 296580 18788
rect 280956 18060 281220 18070
rect 281012 18004 281060 18060
rect 281116 18004 281164 18060
rect 280956 17994 281220 18004
rect 296316 17276 296580 17286
rect 296372 17220 296420 17276
rect 296476 17220 296524 17276
rect 296316 17210 296580 17220
rect 280956 16492 281220 16502
rect 281012 16436 281060 16492
rect 281116 16436 281164 16492
rect 280956 16426 281220 16436
rect 296316 15708 296580 15718
rect 296372 15652 296420 15708
rect 296476 15652 296524 15708
rect 296316 15642 296580 15652
rect 280956 14924 281220 14934
rect 281012 14868 281060 14924
rect 281116 14868 281164 14924
rect 280956 14858 281220 14868
rect 296316 14140 296580 14150
rect 296372 14084 296420 14140
rect 296476 14084 296524 14140
rect 296316 14074 296580 14084
rect 280956 13356 281220 13366
rect 281012 13300 281060 13356
rect 281116 13300 281164 13356
rect 280956 13290 281220 13300
rect 279692 12674 279748 12684
rect 265596 12572 265860 12582
rect 265652 12516 265700 12572
rect 265756 12516 265804 12572
rect 265596 12506 265860 12516
rect 296316 12572 296580 12582
rect 296372 12516 296420 12572
rect 296476 12516 296524 12572
rect 296316 12506 296580 12516
rect 280956 11788 281220 11798
rect 281012 11732 281060 11788
rect 281116 11732 281164 11788
rect 280956 11722 281220 11732
rect 261772 11106 261828 11116
rect 234876 11004 235140 11014
rect 234932 10948 234980 11004
rect 235036 10948 235084 11004
rect 234876 10938 235140 10948
rect 265596 11004 265860 11014
rect 265652 10948 265700 11004
rect 265756 10948 265804 11004
rect 265596 10938 265860 10948
rect 296316 11004 296580 11014
rect 296372 10948 296420 11004
rect 296476 10948 296524 11004
rect 296316 10938 296580 10948
rect 250236 10220 250500 10230
rect 250292 10164 250340 10220
rect 250396 10164 250444 10220
rect 250236 10154 250500 10164
rect 280956 10220 281220 10230
rect 281012 10164 281060 10220
rect 281116 10164 281164 10220
rect 280956 10154 281220 10164
rect 270620 9940 270676 9950
rect 234876 9436 235140 9446
rect 234932 9380 234980 9436
rect 235036 9380 235084 9436
rect 234876 9370 235140 9380
rect 265596 9436 265860 9446
rect 265652 9380 265700 9436
rect 265756 9380 265804 9436
rect 265596 9370 265860 9380
rect 250236 8652 250500 8662
rect 250292 8596 250340 8652
rect 250396 8596 250444 8652
rect 250236 8586 250500 8596
rect 225932 8306 225988 8316
rect 234876 7868 235140 7878
rect 234932 7812 234980 7868
rect 235036 7812 235084 7868
rect 234876 7802 235140 7812
rect 265596 7868 265860 7878
rect 265652 7812 265700 7868
rect 265756 7812 265804 7868
rect 265596 7802 265860 7812
rect 221788 7634 221844 7644
rect 250236 7084 250500 7094
rect 250292 7028 250340 7084
rect 250396 7028 250444 7084
rect 250236 7018 250500 7028
rect 234876 6300 235140 6310
rect 234932 6244 234980 6300
rect 235036 6244 235084 6300
rect 234876 6234 235140 6244
rect 265596 6300 265860 6310
rect 265652 6244 265700 6300
rect 265756 6244 265804 6300
rect 265596 6234 265860 6244
rect 263004 6132 263060 6142
rect 223580 5794 223636 5806
rect 223580 5742 223582 5794
rect 223634 5742 223636 5794
rect 222572 5236 222628 5246
rect 221564 5124 221620 5134
rect 221564 5030 221620 5068
rect 221788 5122 221844 5134
rect 221788 5070 221790 5122
rect 221842 5070 221844 5122
rect 221340 4286 221342 4338
rect 221394 4286 221396 4338
rect 221340 4274 221396 4286
rect 221676 5010 221732 5022
rect 221676 4958 221678 5010
rect 221730 4958 221732 5010
rect 221116 4114 221172 4126
rect 221116 4062 221118 4114
rect 221170 4062 221172 4114
rect 220780 3726 220782 3778
rect 220834 3726 220836 3778
rect 220780 3714 220836 3726
rect 220892 4004 220948 4014
rect 220220 3502 220222 3554
rect 220274 3502 220276 3554
rect 220220 3490 220276 3502
rect 220444 3556 220500 3566
rect 220444 3442 220500 3500
rect 220444 3390 220446 3442
rect 220498 3390 220500 3442
rect 220444 3378 220500 3390
rect 220556 3444 220612 3612
rect 220892 3554 220948 3948
rect 220892 3502 220894 3554
rect 220946 3502 220948 3554
rect 220892 3490 220948 3502
rect 220668 3444 220724 3454
rect 220556 3442 220724 3444
rect 220556 3390 220670 3442
rect 220722 3390 220724 3442
rect 220556 3388 220724 3390
rect 220668 3378 220724 3388
rect 220108 2706 220164 2716
rect 221116 2100 221172 4062
rect 221564 3780 221620 3790
rect 221676 3780 221732 4958
rect 221788 4900 221844 5070
rect 222572 5122 222628 5180
rect 222572 5070 222574 5122
rect 222626 5070 222628 5122
rect 222124 4900 222180 4910
rect 221788 4834 221844 4844
rect 221900 4844 222124 4900
rect 221900 4564 221956 4844
rect 222124 4834 222180 4844
rect 221788 4508 221956 4564
rect 221788 4450 221844 4508
rect 221788 4398 221790 4450
rect 221842 4398 221844 4450
rect 221788 4386 221844 4398
rect 221900 4340 221956 4350
rect 221900 4246 221956 4284
rect 222012 4338 222068 4350
rect 222012 4286 222014 4338
rect 222066 4286 222068 4338
rect 221564 3778 221732 3780
rect 221564 3726 221566 3778
rect 221618 3726 221732 3778
rect 221564 3724 221732 3726
rect 221564 3714 221620 3724
rect 221452 3668 221508 3678
rect 221228 3444 221284 3482
rect 221228 3378 221284 3388
rect 221452 3442 221508 3612
rect 221452 3390 221454 3442
rect 221506 3390 221508 3442
rect 221452 3378 221508 3390
rect 222012 3666 222068 4286
rect 222572 4338 222628 5070
rect 223468 5236 223524 5246
rect 223468 5122 223524 5180
rect 223468 5070 223470 5122
rect 223522 5070 223524 5122
rect 223468 5058 223524 5070
rect 222572 4286 222574 4338
rect 222626 4286 222628 4338
rect 222572 4274 222628 4286
rect 223020 4898 223076 4910
rect 223020 4846 223022 4898
rect 223074 4846 223076 4898
rect 223020 4788 223076 4846
rect 223132 4900 223188 4910
rect 223132 4806 223188 4844
rect 223244 4900 223300 4910
rect 223580 4900 223636 5742
rect 234332 5796 234388 5806
rect 224028 5124 224084 5134
rect 224028 5030 224084 5068
rect 223244 4898 223636 4900
rect 223244 4846 223246 4898
rect 223298 4846 223636 4898
rect 223244 4844 223636 4846
rect 223916 4898 223972 4910
rect 223916 4846 223918 4898
rect 223970 4846 223972 4898
rect 223244 4834 223300 4844
rect 223020 4338 223076 4732
rect 223020 4286 223022 4338
rect 223074 4286 223076 4338
rect 223020 4274 223076 4286
rect 223244 4340 223300 4350
rect 223244 4246 223300 4284
rect 223132 4228 223188 4238
rect 223132 4134 223188 4172
rect 223356 4116 223412 4844
rect 223916 4788 223972 4846
rect 224140 4900 224196 4910
rect 224700 4900 224756 4910
rect 224140 4898 224756 4900
rect 224140 4846 224142 4898
rect 224194 4846 224702 4898
rect 224754 4846 224756 4898
rect 224140 4844 224756 4846
rect 224140 4834 224196 4844
rect 223916 4722 223972 4732
rect 223692 4340 223748 4350
rect 223692 4246 223748 4284
rect 223356 4050 223412 4060
rect 222012 3614 222014 3666
rect 222066 3614 222068 3666
rect 222012 2884 222068 3614
rect 224700 3668 224756 4844
rect 230748 4564 230804 4574
rect 224700 3602 224756 3612
rect 228508 4452 228564 4462
rect 223804 3556 223860 3566
rect 222012 2818 222068 2828
rect 223356 3554 223860 3556
rect 223356 3502 223806 3554
rect 223858 3502 223860 3554
rect 223356 3500 223860 3502
rect 223356 3442 223412 3500
rect 223804 3490 223860 3500
rect 223916 3556 223972 3566
rect 223356 3390 223358 3442
rect 223410 3390 223412 3442
rect 221116 2034 221172 2044
rect 223356 800 223412 3390
rect 223580 3332 223636 3342
rect 223916 3332 223972 3500
rect 223580 3330 223972 3332
rect 223580 3278 223582 3330
rect 223634 3278 223972 3330
rect 223580 3276 223972 3278
rect 225932 3556 225988 3566
rect 227388 3556 227444 3566
rect 223580 3266 223636 3276
rect 225932 2996 225988 3500
rect 225932 2930 225988 2940
rect 226940 3554 227444 3556
rect 226940 3502 227390 3554
rect 227442 3502 227444 3554
rect 226940 3500 227444 3502
rect 226940 3442 226996 3500
rect 227388 3490 227444 3500
rect 226940 3390 226942 3442
rect 226994 3390 226996 3442
rect 226940 800 226996 3390
rect 227164 3332 227220 3342
rect 227164 3238 227220 3276
rect 228508 2548 228564 4396
rect 228508 2482 228564 2492
rect 230524 3442 230580 3454
rect 230524 3390 230526 3442
rect 230578 3390 230580 3442
rect 230524 3108 230580 3390
rect 230748 3330 230804 4508
rect 230748 3278 230750 3330
rect 230802 3278 230804 3330
rect 230748 3266 230804 3278
rect 230972 3554 231028 3566
rect 230972 3502 230974 3554
rect 231026 3502 231028 3554
rect 230972 3108 231028 3502
rect 230524 3052 231028 3108
rect 233548 3442 233604 3454
rect 233548 3390 233550 3442
rect 233602 3390 233604 3442
rect 230524 800 230580 3052
rect 233548 2212 233604 3390
rect 234332 3330 234388 5740
rect 250236 5516 250500 5526
rect 250292 5460 250340 5516
rect 250396 5460 250444 5516
rect 250236 5450 250500 5460
rect 245420 5236 245476 5246
rect 241612 5012 241668 5022
rect 234876 4732 235140 4742
rect 234932 4676 234980 4732
rect 235036 4676 235084 4732
rect 234876 4666 235140 4676
rect 237916 3780 237972 3790
rect 234332 3278 234334 3330
rect 234386 3278 234388 3330
rect 234332 3266 234388 3278
rect 234556 3554 234612 3566
rect 234556 3502 234558 3554
rect 234610 3502 234612 3554
rect 234556 2212 234612 3502
rect 237356 3442 237412 3454
rect 237356 3390 237358 3442
rect 237410 3390 237412 3442
rect 234876 3164 235140 3174
rect 234932 3108 234980 3164
rect 235036 3108 235084 3164
rect 234876 3098 235140 3108
rect 233548 2156 234612 2212
rect 237356 2212 237412 3390
rect 237916 3330 237972 3724
rect 237916 3278 237918 3330
rect 237970 3278 237972 3330
rect 237916 3266 237972 3278
rect 238140 3554 238196 3566
rect 238140 3502 238142 3554
rect 238194 3502 238196 3554
rect 238140 2212 238196 3502
rect 241164 3444 241220 3454
rect 241164 3442 241332 3444
rect 241164 3390 241166 3442
rect 241218 3390 241332 3442
rect 241164 3388 241332 3390
rect 241164 3378 241220 3388
rect 237356 2156 238196 2212
rect 241276 3108 241332 3388
rect 241612 3330 241668 4956
rect 241612 3278 241614 3330
rect 241666 3278 241668 3330
rect 241612 3266 241668 3278
rect 241836 3554 241892 3566
rect 241836 3502 241838 3554
rect 241890 3502 241892 3554
rect 241836 3108 241892 3502
rect 244972 3444 245028 3454
rect 241276 3052 241892 3108
rect 244860 3388 244972 3444
rect 234108 800 234164 2156
rect 237692 800 237748 2156
rect 241276 800 241332 3052
rect 244860 800 244916 3388
rect 244972 3350 245028 3388
rect 245420 3442 245476 5180
rect 249228 4340 249284 4350
rect 245420 3390 245422 3442
rect 245474 3390 245476 3442
rect 245420 3378 245476 3390
rect 245644 3554 245700 3566
rect 245644 3502 245646 3554
rect 245698 3502 245700 3554
rect 245644 3444 245700 3502
rect 248780 3444 248836 3454
rect 245644 3378 245700 3388
rect 248444 3388 248780 3444
rect 248444 800 248500 3388
rect 248780 3350 248836 3388
rect 249228 3442 249284 4284
rect 253036 4116 253092 4126
rect 250236 3948 250500 3958
rect 250292 3892 250340 3948
rect 250396 3892 250444 3948
rect 250236 3882 250500 3892
rect 249228 3390 249230 3442
rect 249282 3390 249284 3442
rect 249228 3378 249284 3390
rect 249340 3668 249396 3678
rect 249340 1316 249396 3612
rect 249452 3554 249508 3566
rect 249452 3502 249454 3554
rect 249506 3502 249508 3554
rect 249452 3444 249508 3502
rect 249452 3378 249508 3388
rect 252588 3442 252644 3454
rect 252588 3390 252590 3442
rect 252642 3390 252644 3442
rect 252588 3108 252644 3390
rect 253036 3330 253092 4060
rect 255836 3780 255892 3790
rect 253036 3278 253038 3330
rect 253090 3278 253092 3330
rect 253036 3266 253092 3278
rect 253260 3554 253316 3566
rect 253260 3502 253262 3554
rect 253314 3502 253316 3554
rect 253260 3108 253316 3502
rect 252588 3052 253316 3108
rect 255612 3442 255668 3454
rect 255612 3390 255614 3442
rect 255666 3390 255668 3442
rect 255612 3108 255668 3390
rect 255836 3330 255892 3724
rect 255836 3278 255838 3330
rect 255890 3278 255892 3330
rect 255836 3266 255892 3278
rect 256060 3554 256116 3566
rect 259644 3556 259700 3566
rect 256060 3502 256062 3554
rect 256114 3502 256116 3554
rect 256060 3108 256116 3502
rect 255612 3052 256116 3108
rect 259196 3554 259700 3556
rect 259196 3502 259646 3554
rect 259698 3502 259700 3554
rect 259196 3500 259700 3502
rect 259196 3442 259252 3500
rect 259644 3490 259700 3500
rect 259196 3390 259198 3442
rect 259250 3390 259252 3442
rect 252588 2212 252644 3052
rect 249340 1250 249396 1260
rect 252028 2156 252644 2212
rect 252028 800 252084 2156
rect 255612 800 255668 3052
rect 259196 800 259252 3390
rect 262780 3442 262836 3454
rect 262780 3390 262782 3442
rect 262834 3390 262836 3442
rect 259420 3330 259476 3342
rect 259420 3278 259422 3330
rect 259474 3278 259476 3330
rect 259420 2772 259476 3278
rect 259420 2706 259476 2716
rect 262780 3108 262836 3390
rect 263004 3330 263060 6076
rect 265596 4732 265860 4742
rect 265652 4676 265700 4732
rect 265756 4676 265804 4732
rect 265596 4666 265860 4676
rect 267036 3666 267092 3678
rect 267036 3614 267038 3666
rect 267090 3614 267092 3666
rect 263004 3278 263006 3330
rect 263058 3278 263060 3330
rect 263004 3266 263060 3278
rect 263228 3554 263284 3566
rect 263228 3502 263230 3554
rect 263282 3502 263284 3554
rect 263228 3108 263284 3502
rect 262780 3052 263284 3108
rect 265356 3444 265412 3454
rect 262780 800 262836 3052
rect 265356 1652 265412 3388
rect 266364 3444 266420 3454
rect 266588 3444 266644 3454
rect 266364 3442 266644 3444
rect 266364 3390 266366 3442
rect 266418 3390 266590 3442
rect 266642 3390 266644 3442
rect 266364 3388 266644 3390
rect 265596 3164 265860 3174
rect 265652 3108 265700 3164
rect 265756 3108 265804 3164
rect 265596 3098 265860 3108
rect 265356 1586 265412 1596
rect 266364 800 266420 3388
rect 266588 3378 266644 3388
rect 267036 3444 267092 3614
rect 270620 3666 270676 9884
rect 296316 9436 296580 9446
rect 296372 9380 296420 9436
rect 296476 9380 296524 9436
rect 296316 9370 296580 9380
rect 280956 8652 281220 8662
rect 281012 8596 281060 8652
rect 281116 8596 281164 8652
rect 280956 8586 281220 8596
rect 296316 7868 296580 7878
rect 296372 7812 296420 7868
rect 296476 7812 296524 7868
rect 296316 7802 296580 7812
rect 280956 7084 281220 7094
rect 281012 7028 281060 7084
rect 281116 7028 281164 7084
rect 280956 7018 281220 7028
rect 296316 6300 296580 6310
rect 296372 6244 296420 6300
rect 296476 6244 296524 6300
rect 296316 6234 296580 6244
rect 292124 6020 292180 6030
rect 280956 5516 281220 5526
rect 281012 5460 281060 5516
rect 281116 5460 281164 5516
rect 280956 5450 281220 5460
rect 288540 4452 288596 4462
rect 280956 3948 281220 3958
rect 281012 3892 281060 3948
rect 281116 3892 281164 3948
rect 280956 3882 281220 3892
rect 270620 3614 270622 3666
rect 270674 3614 270676 3666
rect 270620 3602 270676 3614
rect 281372 3780 281428 3790
rect 281372 3666 281428 3724
rect 281372 3614 281374 3666
rect 281426 3614 281428 3666
rect 281372 3602 281428 3614
rect 288540 3666 288596 4396
rect 288540 3614 288542 3666
rect 288594 3614 288596 3666
rect 288540 3602 288596 3614
rect 292124 3666 292180 5964
rect 296316 4732 296580 4742
rect 296372 4676 296420 4732
rect 296476 4676 296524 4732
rect 296316 4666 296580 4676
rect 292124 3614 292126 3666
rect 292178 3614 292180 3666
rect 292124 3602 292180 3614
rect 285068 3556 285124 3566
rect 285068 3462 285124 3500
rect 267036 3378 267092 3388
rect 269948 3444 270004 3454
rect 270172 3444 270228 3454
rect 269948 3442 270228 3444
rect 269948 3390 269950 3442
rect 270002 3390 270174 3442
rect 270226 3390 270228 3442
rect 269948 3388 270228 3390
rect 269948 800 270004 3388
rect 270172 3378 270228 3388
rect 273532 3444 273588 3454
rect 273756 3444 273812 3454
rect 273532 3442 273812 3444
rect 273532 3390 273534 3442
rect 273586 3390 273758 3442
rect 273810 3390 273812 3442
rect 273532 3388 273812 3390
rect 273532 800 273588 3388
rect 273756 3378 273812 3388
rect 274316 3442 274372 3454
rect 274316 3390 274318 3442
rect 274370 3390 274372 3442
rect 274316 1428 274372 3390
rect 274316 1362 274372 1372
rect 277116 3444 277172 3454
rect 277340 3444 277396 3454
rect 277116 3442 277396 3444
rect 277116 3390 277118 3442
rect 277170 3390 277342 3442
rect 277394 3390 277396 3442
rect 277116 3388 277396 3390
rect 277116 800 277172 3388
rect 277340 3378 277396 3388
rect 277900 3442 277956 3454
rect 277900 3390 277902 3442
rect 277954 3390 277956 3442
rect 277900 3332 277956 3390
rect 277900 3266 277956 3276
rect 280700 3444 280756 3454
rect 280924 3444 280980 3454
rect 280700 3442 280980 3444
rect 280700 3390 280702 3442
rect 280754 3390 280926 3442
rect 280978 3390 280980 3442
rect 280700 3388 280980 3390
rect 280700 800 280756 3388
rect 280924 3378 280980 3388
rect 284284 3444 284340 3454
rect 284508 3444 284564 3454
rect 284284 3442 284564 3444
rect 284284 3390 284286 3442
rect 284338 3390 284510 3442
rect 284562 3390 284564 3442
rect 284284 3388 284564 3390
rect 284284 800 284340 3388
rect 284508 3378 284564 3388
rect 287868 3444 287924 3454
rect 288092 3444 288148 3454
rect 287868 3442 288148 3444
rect 287868 3390 287870 3442
rect 287922 3390 288094 3442
rect 288146 3390 288148 3442
rect 287868 3388 288148 3390
rect 287868 800 287924 3388
rect 288092 3378 288148 3388
rect 291452 3444 291508 3454
rect 291676 3444 291732 3454
rect 291452 3442 291732 3444
rect 291452 3390 291454 3442
rect 291506 3390 291678 3442
rect 291730 3390 291732 3442
rect 291452 3388 291732 3390
rect 291452 800 291508 3388
rect 291676 3378 291732 3388
rect 296316 3164 296580 3174
rect 296372 3108 296420 3164
rect 296476 3108 296524 3164
rect 296316 3098 296580 3108
rect 98252 700 98644 756
rect 101472 0 101584 800
rect 105056 0 105168 800
rect 108640 0 108752 800
rect 112224 0 112336 800
rect 115808 0 115920 800
rect 119392 0 119504 800
rect 122976 0 123088 800
rect 126560 0 126672 800
rect 130144 0 130256 800
rect 133728 0 133840 800
rect 137312 0 137424 800
rect 140896 0 141008 800
rect 144480 0 144592 800
rect 148064 0 148176 800
rect 151648 0 151760 800
rect 155232 0 155344 800
rect 158816 0 158928 800
rect 162400 0 162512 800
rect 165984 0 166096 800
rect 169568 0 169680 800
rect 173152 0 173264 800
rect 176736 0 176848 800
rect 180320 0 180432 800
rect 183904 0 184016 800
rect 187488 0 187600 800
rect 191072 0 191184 800
rect 194656 0 194768 800
rect 198240 0 198352 800
rect 201824 0 201936 800
rect 205408 0 205520 800
rect 208992 0 209104 800
rect 212576 0 212688 800
rect 216160 0 216272 800
rect 219744 0 219856 800
rect 223328 0 223440 800
rect 226912 0 227024 800
rect 230496 0 230608 800
rect 234080 0 234192 800
rect 237664 0 237776 800
rect 241248 0 241360 800
rect 244832 0 244944 800
rect 248416 0 248528 800
rect 252000 0 252112 800
rect 255584 0 255696 800
rect 259168 0 259280 800
rect 262752 0 262864 800
rect 266336 0 266448 800
rect 269920 0 270032 800
rect 273504 0 273616 800
rect 277088 0 277200 800
rect 280672 0 280784 800
rect 284256 0 284368 800
rect 287840 0 287952 800
rect 291424 0 291536 800
<< via2 >>
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 7420 51996 7476 52052
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 19180 56306 19236 56308
rect 19180 56254 19182 56306
rect 19182 56254 19234 56306
rect 19234 56254 19236 56306
rect 19180 56252 19236 56254
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35084 19292 35140 19348
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 40460 15932 40516 15988
rect 43820 24444 43876 24500
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 29708 9212 29764 9268
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 25116 7532 25172 7588
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 8316 3388 8372 3444
rect 10108 3442 10164 3444
rect 10108 3390 10110 3442
rect 10110 3390 10162 3442
rect 10162 3390 10164 3442
rect 10108 3388 10164 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 43036 3612 43092 3668
rect 51772 55970 51828 55972
rect 51772 55918 51774 55970
rect 51774 55918 51826 55970
rect 51826 55918 51828 55970
rect 51772 55916 51828 55918
rect 52892 55916 52948 55972
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 45836 20972 45892 21028
rect 47628 26012 47684 26068
rect 43820 3666 43876 3668
rect 43820 3614 43822 3666
rect 43822 3614 43874 3666
rect 43874 3614 43876 3666
rect 43820 3612 43876 3614
rect 46844 3612 46900 3668
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 52892 22876 52948 22932
rect 54348 41132 54404 41188
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 69356 55916 69412 55972
rect 70476 55970 70532 55972
rect 70476 55918 70478 55970
rect 70478 55918 70530 55970
rect 70530 55918 70532 55970
rect 70476 55916 70532 55918
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 61964 55468 62020 55524
rect 73052 55916 73108 55972
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 68236 36204 68292 36260
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 60956 32732 61012 32788
rect 56588 5852 56644 5908
rect 57260 31052 57316 31108
rect 47628 3666 47684 3668
rect 47628 3614 47630 3666
rect 47630 3614 47682 3666
rect 47682 3614 47684 3666
rect 47628 3612 47684 3614
rect 50540 3554 50596 3556
rect 50540 3502 50542 3554
rect 50542 3502 50594 3554
rect 50594 3502 50596 3554
rect 50540 3500 50596 3502
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 59612 29372 59668 29428
rect 59612 3500 59668 3556
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 62076 3612 62132 3668
rect 62860 3666 62916 3668
rect 62860 3614 62862 3666
rect 62862 3614 62914 3666
rect 62914 3614 62916 3666
rect 62860 3612 62916 3614
rect 65212 3612 65268 3668
rect 65772 3666 65828 3668
rect 65772 3614 65774 3666
rect 65774 3614 65826 3666
rect 65826 3614 65828 3666
rect 65772 3612 65828 3614
rect 65660 3388 65716 3444
rect 69580 34636 69636 34692
rect 68236 3612 68292 3668
rect 69244 3612 69300 3668
rect 68908 3554 68964 3556
rect 68908 3502 68910 3554
rect 68910 3502 68962 3554
rect 68962 3502 68964 3554
rect 68908 3500 68964 3502
rect 66668 3388 66724 3444
rect 81276 56474 81332 56476
rect 81276 56422 81278 56474
rect 81278 56422 81330 56474
rect 81330 56422 81332 56474
rect 81276 56420 81332 56422
rect 81380 56474 81436 56476
rect 81380 56422 81382 56474
rect 81382 56422 81434 56474
rect 81434 56422 81436 56474
rect 81380 56420 81436 56422
rect 81484 56474 81540 56476
rect 81484 56422 81486 56474
rect 81486 56422 81538 56474
rect 81538 56422 81540 56474
rect 81484 56420 81540 56422
rect 80444 55916 80500 55972
rect 81004 55970 81060 55972
rect 81004 55918 81006 55970
rect 81006 55918 81058 55970
rect 81058 55918 81060 55970
rect 81004 55916 81060 55918
rect 84924 56082 84980 56084
rect 84924 56030 84926 56082
rect 84926 56030 84978 56082
rect 84978 56030 84980 56082
rect 84924 56028 84980 56030
rect 85708 56082 85764 56084
rect 85708 56030 85710 56082
rect 85710 56030 85762 56082
rect 85762 56030 85764 56082
rect 85708 56028 85764 56030
rect 83132 55916 83188 55972
rect 81276 54906 81332 54908
rect 81276 54854 81278 54906
rect 81278 54854 81330 54906
rect 81330 54854 81332 54906
rect 81276 54852 81332 54854
rect 81380 54906 81436 54908
rect 81380 54854 81382 54906
rect 81382 54854 81434 54906
rect 81434 54854 81436 54906
rect 81380 54852 81436 54854
rect 81484 54906 81540 54908
rect 81484 54854 81486 54906
rect 81486 54854 81538 54906
rect 81538 54854 81540 54906
rect 81484 54852 81540 54854
rect 81276 53338 81332 53340
rect 81276 53286 81278 53338
rect 81278 53286 81330 53338
rect 81330 53286 81332 53338
rect 81276 53284 81332 53286
rect 81380 53338 81436 53340
rect 81380 53286 81382 53338
rect 81382 53286 81434 53338
rect 81434 53286 81436 53338
rect 81380 53284 81436 53286
rect 81484 53338 81540 53340
rect 81484 53286 81486 53338
rect 81486 53286 81538 53338
rect 81538 53286 81540 53338
rect 81484 53284 81540 53286
rect 81276 51770 81332 51772
rect 81276 51718 81278 51770
rect 81278 51718 81330 51770
rect 81330 51718 81332 51770
rect 81276 51716 81332 51718
rect 81380 51770 81436 51772
rect 81380 51718 81382 51770
rect 81382 51718 81434 51770
rect 81434 51718 81436 51770
rect 81380 51716 81436 51718
rect 81484 51770 81540 51772
rect 81484 51718 81486 51770
rect 81486 51718 81538 51770
rect 81538 51718 81540 51770
rect 81484 51716 81540 51718
rect 81276 50202 81332 50204
rect 81276 50150 81278 50202
rect 81278 50150 81330 50202
rect 81330 50150 81332 50202
rect 81276 50148 81332 50150
rect 81380 50202 81436 50204
rect 81380 50150 81382 50202
rect 81382 50150 81434 50202
rect 81434 50150 81436 50202
rect 81380 50148 81436 50150
rect 81484 50202 81540 50204
rect 81484 50150 81486 50202
rect 81486 50150 81538 50202
rect 81538 50150 81540 50202
rect 81484 50148 81540 50150
rect 81276 48634 81332 48636
rect 81276 48582 81278 48634
rect 81278 48582 81330 48634
rect 81330 48582 81332 48634
rect 81276 48580 81332 48582
rect 81380 48634 81436 48636
rect 81380 48582 81382 48634
rect 81382 48582 81434 48634
rect 81434 48582 81436 48634
rect 81380 48580 81436 48582
rect 81484 48634 81540 48636
rect 81484 48582 81486 48634
rect 81486 48582 81538 48634
rect 81538 48582 81540 48634
rect 81484 48580 81540 48582
rect 81276 47066 81332 47068
rect 81276 47014 81278 47066
rect 81278 47014 81330 47066
rect 81330 47014 81332 47066
rect 81276 47012 81332 47014
rect 81380 47066 81436 47068
rect 81380 47014 81382 47066
rect 81382 47014 81434 47066
rect 81434 47014 81436 47066
rect 81380 47012 81436 47014
rect 81484 47066 81540 47068
rect 81484 47014 81486 47066
rect 81486 47014 81538 47066
rect 81538 47014 81540 47066
rect 81484 47012 81540 47014
rect 81276 45498 81332 45500
rect 81276 45446 81278 45498
rect 81278 45446 81330 45498
rect 81330 45446 81332 45498
rect 81276 45444 81332 45446
rect 81380 45498 81436 45500
rect 81380 45446 81382 45498
rect 81382 45446 81434 45498
rect 81434 45446 81436 45498
rect 81380 45444 81436 45446
rect 81484 45498 81540 45500
rect 81484 45446 81486 45498
rect 81486 45446 81538 45498
rect 81538 45446 81540 45498
rect 81484 45444 81540 45446
rect 81276 43930 81332 43932
rect 81276 43878 81278 43930
rect 81278 43878 81330 43930
rect 81330 43878 81332 43930
rect 81276 43876 81332 43878
rect 81380 43930 81436 43932
rect 81380 43878 81382 43930
rect 81382 43878 81434 43930
rect 81434 43878 81436 43930
rect 81380 43876 81436 43878
rect 81484 43930 81540 43932
rect 81484 43878 81486 43930
rect 81486 43878 81538 43930
rect 81538 43878 81540 43930
rect 81484 43876 81540 43878
rect 81276 42362 81332 42364
rect 81276 42310 81278 42362
rect 81278 42310 81330 42362
rect 81330 42310 81332 42362
rect 81276 42308 81332 42310
rect 81380 42362 81436 42364
rect 81380 42310 81382 42362
rect 81382 42310 81434 42362
rect 81434 42310 81436 42362
rect 81380 42308 81436 42310
rect 81484 42362 81540 42364
rect 81484 42310 81486 42362
rect 81486 42310 81538 42362
rect 81538 42310 81540 42362
rect 81484 42308 81540 42310
rect 81276 40794 81332 40796
rect 81276 40742 81278 40794
rect 81278 40742 81330 40794
rect 81330 40742 81332 40794
rect 81276 40740 81332 40742
rect 81380 40794 81436 40796
rect 81380 40742 81382 40794
rect 81382 40742 81434 40794
rect 81434 40742 81436 40794
rect 81380 40740 81436 40742
rect 81484 40794 81540 40796
rect 81484 40742 81486 40794
rect 81486 40742 81538 40794
rect 81538 40742 81540 40794
rect 81484 40740 81540 40742
rect 81276 39226 81332 39228
rect 81276 39174 81278 39226
rect 81278 39174 81330 39226
rect 81330 39174 81332 39226
rect 81276 39172 81332 39174
rect 81380 39226 81436 39228
rect 81380 39174 81382 39226
rect 81382 39174 81434 39226
rect 81434 39174 81436 39226
rect 81380 39172 81436 39174
rect 81484 39226 81540 39228
rect 81484 39174 81486 39226
rect 81486 39174 81538 39226
rect 81538 39174 81540 39226
rect 81484 39172 81540 39174
rect 81276 37658 81332 37660
rect 81276 37606 81278 37658
rect 81278 37606 81330 37658
rect 81330 37606 81332 37658
rect 81276 37604 81332 37606
rect 81380 37658 81436 37660
rect 81380 37606 81382 37658
rect 81382 37606 81434 37658
rect 81434 37606 81436 37658
rect 81380 37604 81436 37606
rect 81484 37658 81540 37660
rect 81484 37606 81486 37658
rect 81486 37606 81538 37658
rect 81538 37606 81540 37658
rect 81484 37604 81540 37606
rect 81276 36090 81332 36092
rect 81276 36038 81278 36090
rect 81278 36038 81330 36090
rect 81330 36038 81332 36090
rect 81276 36036 81332 36038
rect 81380 36090 81436 36092
rect 81380 36038 81382 36090
rect 81382 36038 81434 36090
rect 81434 36038 81436 36090
rect 81380 36036 81436 36038
rect 81484 36090 81540 36092
rect 81484 36038 81486 36090
rect 81486 36038 81538 36090
rect 81538 36038 81540 36090
rect 81484 36036 81540 36038
rect 81276 34522 81332 34524
rect 81276 34470 81278 34522
rect 81278 34470 81330 34522
rect 81330 34470 81332 34522
rect 81276 34468 81332 34470
rect 81380 34522 81436 34524
rect 81380 34470 81382 34522
rect 81382 34470 81434 34522
rect 81434 34470 81436 34522
rect 81380 34468 81436 34470
rect 81484 34522 81540 34524
rect 81484 34470 81486 34522
rect 81486 34470 81538 34522
rect 81538 34470 81540 34522
rect 81484 34468 81540 34470
rect 81276 32954 81332 32956
rect 81276 32902 81278 32954
rect 81278 32902 81330 32954
rect 81330 32902 81332 32954
rect 81276 32900 81332 32902
rect 81380 32954 81436 32956
rect 81380 32902 81382 32954
rect 81382 32902 81434 32954
rect 81434 32902 81436 32954
rect 81380 32900 81436 32902
rect 81484 32954 81540 32956
rect 81484 32902 81486 32954
rect 81486 32902 81538 32954
rect 81538 32902 81540 32954
rect 81484 32900 81540 32902
rect 81276 31386 81332 31388
rect 81276 31334 81278 31386
rect 81278 31334 81330 31386
rect 81330 31334 81332 31386
rect 81276 31332 81332 31334
rect 81380 31386 81436 31388
rect 81380 31334 81382 31386
rect 81382 31334 81434 31386
rect 81434 31334 81436 31386
rect 81380 31332 81436 31334
rect 81484 31386 81540 31388
rect 81484 31334 81486 31386
rect 81486 31334 81538 31386
rect 81538 31334 81540 31386
rect 81484 31332 81540 31334
rect 81276 29818 81332 29820
rect 81276 29766 81278 29818
rect 81278 29766 81330 29818
rect 81330 29766 81332 29818
rect 81276 29764 81332 29766
rect 81380 29818 81436 29820
rect 81380 29766 81382 29818
rect 81382 29766 81434 29818
rect 81434 29766 81436 29818
rect 81380 29764 81436 29766
rect 81484 29818 81540 29820
rect 81484 29766 81486 29818
rect 81486 29766 81538 29818
rect 81538 29766 81540 29818
rect 81484 29764 81540 29766
rect 81276 28250 81332 28252
rect 81276 28198 81278 28250
rect 81278 28198 81330 28250
rect 81330 28198 81332 28250
rect 81276 28196 81332 28198
rect 81380 28250 81436 28252
rect 81380 28198 81382 28250
rect 81382 28198 81434 28250
rect 81434 28198 81436 28250
rect 81380 28196 81436 28198
rect 81484 28250 81540 28252
rect 81484 28198 81486 28250
rect 81486 28198 81538 28250
rect 81538 28198 81540 28250
rect 81484 28196 81540 28198
rect 81276 26682 81332 26684
rect 81276 26630 81278 26682
rect 81278 26630 81330 26682
rect 81330 26630 81332 26682
rect 81276 26628 81332 26630
rect 81380 26682 81436 26684
rect 81380 26630 81382 26682
rect 81382 26630 81434 26682
rect 81434 26630 81436 26682
rect 81380 26628 81436 26630
rect 81484 26682 81540 26684
rect 81484 26630 81486 26682
rect 81486 26630 81538 26682
rect 81538 26630 81540 26682
rect 81484 26628 81540 26630
rect 81276 25114 81332 25116
rect 81276 25062 81278 25114
rect 81278 25062 81330 25114
rect 81330 25062 81332 25114
rect 81276 25060 81332 25062
rect 81380 25114 81436 25116
rect 81380 25062 81382 25114
rect 81382 25062 81434 25114
rect 81434 25062 81436 25114
rect 81380 25060 81436 25062
rect 81484 25114 81540 25116
rect 81484 25062 81486 25114
rect 81486 25062 81538 25114
rect 81538 25062 81540 25114
rect 81484 25060 81540 25062
rect 81276 23546 81332 23548
rect 81276 23494 81278 23546
rect 81278 23494 81330 23546
rect 81330 23494 81332 23546
rect 81276 23492 81332 23494
rect 81380 23546 81436 23548
rect 81380 23494 81382 23546
rect 81382 23494 81434 23546
rect 81434 23494 81436 23546
rect 81380 23492 81436 23494
rect 81484 23546 81540 23548
rect 81484 23494 81486 23546
rect 81486 23494 81538 23546
rect 81538 23494 81540 23546
rect 81484 23492 81540 23494
rect 81276 21978 81332 21980
rect 81276 21926 81278 21978
rect 81278 21926 81330 21978
rect 81330 21926 81332 21978
rect 81276 21924 81332 21926
rect 81380 21978 81436 21980
rect 81380 21926 81382 21978
rect 81382 21926 81434 21978
rect 81434 21926 81436 21978
rect 81380 21924 81436 21926
rect 81484 21978 81540 21980
rect 81484 21926 81486 21978
rect 81486 21926 81538 21978
rect 81538 21926 81540 21978
rect 81484 21924 81540 21926
rect 81276 20410 81332 20412
rect 81276 20358 81278 20410
rect 81278 20358 81330 20410
rect 81330 20358 81332 20410
rect 81276 20356 81332 20358
rect 81380 20410 81436 20412
rect 81380 20358 81382 20410
rect 81382 20358 81434 20410
rect 81434 20358 81436 20410
rect 81380 20356 81436 20358
rect 81484 20410 81540 20412
rect 81484 20358 81486 20410
rect 81486 20358 81538 20410
rect 81538 20358 81540 20410
rect 81484 20356 81540 20358
rect 75180 14252 75236 14308
rect 78652 19292 78708 19348
rect 73052 12684 73108 12740
rect 73388 11228 73444 11284
rect 71148 7532 71204 7588
rect 70476 3666 70532 3668
rect 70476 3614 70478 3666
rect 70478 3614 70530 3666
rect 70530 3614 70532 3666
rect 70476 3612 70532 3614
rect 69580 3500 69636 3556
rect 74844 9212 74900 9268
rect 75404 4284 75460 4340
rect 76636 4338 76692 4340
rect 76636 4286 76638 4338
rect 76638 4286 76690 4338
rect 76690 4286 76692 4338
rect 76636 4284 76692 4286
rect 71708 3500 71764 3556
rect 76412 4060 76468 4116
rect 74060 3554 74116 3556
rect 74060 3502 74062 3554
rect 74062 3502 74114 3554
rect 74114 3502 74116 3554
rect 74060 3500 74116 3502
rect 72940 3388 72996 3444
rect 75628 3442 75684 3444
rect 75628 3390 75630 3442
rect 75630 3390 75682 3442
rect 75682 3390 75684 3442
rect 75628 3388 75684 3390
rect 77644 4114 77700 4116
rect 77644 4062 77646 4114
rect 77646 4062 77698 4114
rect 77698 4062 77700 4114
rect 77644 4060 77700 4062
rect 81276 18842 81332 18844
rect 81276 18790 81278 18842
rect 81278 18790 81330 18842
rect 81330 18790 81332 18842
rect 81276 18788 81332 18790
rect 81380 18842 81436 18844
rect 81380 18790 81382 18842
rect 81382 18790 81434 18842
rect 81434 18790 81436 18842
rect 81380 18788 81436 18790
rect 81484 18842 81540 18844
rect 81484 18790 81486 18842
rect 81486 18790 81538 18842
rect 81538 18790 81540 18842
rect 81484 18788 81540 18790
rect 83132 17612 83188 17668
rect 85036 20972 85092 21028
rect 81276 17274 81332 17276
rect 81276 17222 81278 17274
rect 81278 17222 81330 17274
rect 81330 17222 81332 17274
rect 81276 17220 81332 17222
rect 81380 17274 81436 17276
rect 81380 17222 81382 17274
rect 81382 17222 81434 17274
rect 81434 17222 81436 17274
rect 81380 17220 81436 17222
rect 81484 17274 81540 17276
rect 81484 17222 81486 17274
rect 81486 17222 81538 17274
rect 81538 17222 81540 17274
rect 81484 17220 81540 17222
rect 83132 15932 83188 15988
rect 81276 15706 81332 15708
rect 81276 15654 81278 15706
rect 81278 15654 81330 15706
rect 81330 15654 81332 15706
rect 81276 15652 81332 15654
rect 81380 15706 81436 15708
rect 81380 15654 81382 15706
rect 81382 15654 81434 15706
rect 81434 15654 81436 15706
rect 81380 15652 81436 15654
rect 81484 15706 81540 15708
rect 81484 15654 81486 15706
rect 81486 15654 81538 15706
rect 81538 15654 81540 15706
rect 81484 15652 81540 15654
rect 81276 14138 81332 14140
rect 81276 14086 81278 14138
rect 81278 14086 81330 14138
rect 81330 14086 81332 14138
rect 81276 14084 81332 14086
rect 81380 14138 81436 14140
rect 81380 14086 81382 14138
rect 81382 14086 81434 14138
rect 81434 14086 81436 14138
rect 81380 14084 81436 14086
rect 81484 14138 81540 14140
rect 81484 14086 81486 14138
rect 81486 14086 81538 14138
rect 81538 14086 81540 14138
rect 81484 14084 81540 14086
rect 81276 12570 81332 12572
rect 81276 12518 81278 12570
rect 81278 12518 81330 12570
rect 81330 12518 81332 12570
rect 81276 12516 81332 12518
rect 81380 12570 81436 12572
rect 81380 12518 81382 12570
rect 81382 12518 81434 12570
rect 81434 12518 81436 12570
rect 81380 12516 81436 12518
rect 81484 12570 81540 12572
rect 81484 12518 81486 12570
rect 81486 12518 81538 12570
rect 81538 12518 81540 12570
rect 81484 12516 81540 12518
rect 81276 11002 81332 11004
rect 81276 10950 81278 11002
rect 81278 10950 81330 11002
rect 81330 10950 81332 11002
rect 81276 10948 81332 10950
rect 81380 11002 81436 11004
rect 81380 10950 81382 11002
rect 81382 10950 81434 11002
rect 81434 10950 81436 11002
rect 81380 10948 81436 10950
rect 81484 11002 81540 11004
rect 81484 10950 81486 11002
rect 81486 10950 81538 11002
rect 81538 10950 81540 11002
rect 81484 10948 81540 10950
rect 81276 9434 81332 9436
rect 81276 9382 81278 9434
rect 81278 9382 81330 9434
rect 81330 9382 81332 9434
rect 81276 9380 81332 9382
rect 81380 9434 81436 9436
rect 81380 9382 81382 9434
rect 81382 9382 81434 9434
rect 81434 9382 81436 9434
rect 81380 9380 81436 9382
rect 81484 9434 81540 9436
rect 81484 9382 81486 9434
rect 81486 9382 81538 9434
rect 81538 9382 81540 9434
rect 81484 9380 81540 9382
rect 81276 7866 81332 7868
rect 81276 7814 81278 7866
rect 81278 7814 81330 7866
rect 81330 7814 81332 7866
rect 81276 7812 81332 7814
rect 81380 7866 81436 7868
rect 81380 7814 81382 7866
rect 81382 7814 81434 7866
rect 81434 7814 81436 7866
rect 81380 7812 81436 7814
rect 81484 7866 81540 7868
rect 81484 7814 81486 7866
rect 81486 7814 81538 7866
rect 81538 7814 81540 7866
rect 81484 7812 81540 7814
rect 81276 6298 81332 6300
rect 81276 6246 81278 6298
rect 81278 6246 81330 6298
rect 81330 6246 81332 6298
rect 81276 6244 81332 6246
rect 81380 6298 81436 6300
rect 81380 6246 81382 6298
rect 81382 6246 81434 6298
rect 81434 6246 81436 6298
rect 81380 6244 81436 6246
rect 81484 6298 81540 6300
rect 81484 6246 81486 6298
rect 81486 6246 81538 6298
rect 81538 6246 81540 6298
rect 81484 6244 81540 6246
rect 81276 4730 81332 4732
rect 81276 4678 81278 4730
rect 81278 4678 81330 4730
rect 81330 4678 81332 4730
rect 81276 4676 81332 4678
rect 81380 4730 81436 4732
rect 81380 4678 81382 4730
rect 81382 4678 81434 4730
rect 81434 4678 81436 4730
rect 81380 4676 81436 4678
rect 81484 4730 81540 4732
rect 81484 4678 81486 4730
rect 81486 4678 81538 4730
rect 81538 4678 81540 4730
rect 81484 4676 81540 4678
rect 79996 4060 80052 4116
rect 81228 4114 81284 4116
rect 81228 4062 81230 4114
rect 81230 4062 81282 4114
rect 81282 4062 81284 4114
rect 81228 4060 81284 4062
rect 88060 55916 88116 55972
rect 89516 55970 89572 55972
rect 89516 55918 89518 55970
rect 89518 55918 89570 55970
rect 89570 55918 89572 55970
rect 89516 55916 89572 55918
rect 91644 55468 91700 55524
rect 85708 11116 85764 11172
rect 88732 22876 88788 22932
rect 85036 4396 85092 4452
rect 86716 4450 86772 4452
rect 86716 4398 86718 4450
rect 86718 4398 86770 4450
rect 86770 4398 86772 4450
rect 86716 4396 86772 4398
rect 83580 4060 83636 4116
rect 81276 3162 81332 3164
rect 81276 3110 81278 3162
rect 81278 3110 81330 3162
rect 81330 3110 81332 3162
rect 81276 3108 81332 3110
rect 81380 3162 81436 3164
rect 81380 3110 81382 3162
rect 81382 3110 81434 3162
rect 81434 3110 81436 3162
rect 81380 3108 81436 3110
rect 81484 3162 81540 3164
rect 81484 3110 81486 3162
rect 81486 3110 81538 3162
rect 81538 3110 81540 3162
rect 81484 3108 81540 3110
rect 84812 4114 84868 4116
rect 84812 4062 84814 4114
rect 84814 4062 84866 4114
rect 84866 4062 84868 4114
rect 84812 4060 84868 4062
rect 87052 4284 87108 4340
rect 87948 4338 88004 4340
rect 87948 4286 87950 4338
rect 87950 4286 88002 4338
rect 88002 4286 88004 4338
rect 87948 4284 88004 4286
rect 87164 4172 87220 4228
rect 96236 55916 96292 55972
rect 97132 55970 97188 55972
rect 97132 55918 97134 55970
rect 97134 55918 97186 55970
rect 97186 55918 97188 55970
rect 97132 55916 97188 55918
rect 96636 55690 96692 55692
rect 96636 55638 96638 55690
rect 96638 55638 96690 55690
rect 96690 55638 96692 55690
rect 96636 55636 96692 55638
rect 96740 55690 96796 55692
rect 96740 55638 96742 55690
rect 96742 55638 96794 55690
rect 96794 55638 96796 55690
rect 96740 55636 96796 55638
rect 96844 55690 96900 55692
rect 96844 55638 96846 55690
rect 96846 55638 96898 55690
rect 96898 55638 96900 55690
rect 96844 55636 96900 55638
rect 98812 55356 98868 55412
rect 99932 55916 99988 55972
rect 111996 56474 112052 56476
rect 111996 56422 111998 56474
rect 111998 56422 112050 56474
rect 112050 56422 112052 56474
rect 111996 56420 112052 56422
rect 112100 56474 112156 56476
rect 112100 56422 112102 56474
rect 112102 56422 112154 56474
rect 112154 56422 112156 56474
rect 112100 56420 112156 56422
rect 112204 56474 112260 56476
rect 112204 56422 112206 56474
rect 112206 56422 112258 56474
rect 112258 56422 112260 56474
rect 112204 56420 112260 56422
rect 126252 56194 126308 56196
rect 126252 56142 126254 56194
rect 126254 56142 126306 56194
rect 126306 56142 126308 56194
rect 126252 56140 126308 56142
rect 127820 56140 127876 56196
rect 96636 54122 96692 54124
rect 96636 54070 96638 54122
rect 96638 54070 96690 54122
rect 96690 54070 96692 54122
rect 96636 54068 96692 54070
rect 96740 54122 96796 54124
rect 96740 54070 96742 54122
rect 96742 54070 96794 54122
rect 96794 54070 96796 54122
rect 96740 54068 96796 54070
rect 96844 54122 96900 54124
rect 96844 54070 96846 54122
rect 96846 54070 96898 54122
rect 96898 54070 96900 54122
rect 96844 54068 96900 54070
rect 96636 52554 96692 52556
rect 96636 52502 96638 52554
rect 96638 52502 96690 52554
rect 96690 52502 96692 52554
rect 96636 52500 96692 52502
rect 96740 52554 96796 52556
rect 96740 52502 96742 52554
rect 96742 52502 96794 52554
rect 96794 52502 96796 52554
rect 96740 52500 96796 52502
rect 96844 52554 96900 52556
rect 96844 52502 96846 52554
rect 96846 52502 96898 52554
rect 96898 52502 96900 52554
rect 96844 52500 96900 52502
rect 96636 50986 96692 50988
rect 96636 50934 96638 50986
rect 96638 50934 96690 50986
rect 96690 50934 96692 50986
rect 96636 50932 96692 50934
rect 96740 50986 96796 50988
rect 96740 50934 96742 50986
rect 96742 50934 96794 50986
rect 96794 50934 96796 50986
rect 96740 50932 96796 50934
rect 96844 50986 96900 50988
rect 96844 50934 96846 50986
rect 96846 50934 96898 50986
rect 96898 50934 96900 50986
rect 96844 50932 96900 50934
rect 96636 49418 96692 49420
rect 96636 49366 96638 49418
rect 96638 49366 96690 49418
rect 96690 49366 96692 49418
rect 96636 49364 96692 49366
rect 96740 49418 96796 49420
rect 96740 49366 96742 49418
rect 96742 49366 96794 49418
rect 96794 49366 96796 49418
rect 96740 49364 96796 49366
rect 96844 49418 96900 49420
rect 96844 49366 96846 49418
rect 96846 49366 96898 49418
rect 96898 49366 96900 49418
rect 96844 49364 96900 49366
rect 96636 47850 96692 47852
rect 96636 47798 96638 47850
rect 96638 47798 96690 47850
rect 96690 47798 96692 47850
rect 96636 47796 96692 47798
rect 96740 47850 96796 47852
rect 96740 47798 96742 47850
rect 96742 47798 96794 47850
rect 96794 47798 96796 47850
rect 96740 47796 96796 47798
rect 96844 47850 96900 47852
rect 96844 47798 96846 47850
rect 96846 47798 96898 47850
rect 96898 47798 96900 47850
rect 96844 47796 96900 47798
rect 96636 46282 96692 46284
rect 96636 46230 96638 46282
rect 96638 46230 96690 46282
rect 96690 46230 96692 46282
rect 96636 46228 96692 46230
rect 96740 46282 96796 46284
rect 96740 46230 96742 46282
rect 96742 46230 96794 46282
rect 96794 46230 96796 46282
rect 96740 46228 96796 46230
rect 96844 46282 96900 46284
rect 96844 46230 96846 46282
rect 96846 46230 96898 46282
rect 96898 46230 96900 46282
rect 96844 46228 96900 46230
rect 96636 44714 96692 44716
rect 96636 44662 96638 44714
rect 96638 44662 96690 44714
rect 96690 44662 96692 44714
rect 96636 44660 96692 44662
rect 96740 44714 96796 44716
rect 96740 44662 96742 44714
rect 96742 44662 96794 44714
rect 96794 44662 96796 44714
rect 96740 44660 96796 44662
rect 96844 44714 96900 44716
rect 96844 44662 96846 44714
rect 96846 44662 96898 44714
rect 96898 44662 96900 44714
rect 96844 44660 96900 44662
rect 96636 43146 96692 43148
rect 96636 43094 96638 43146
rect 96638 43094 96690 43146
rect 96690 43094 96692 43146
rect 96636 43092 96692 43094
rect 96740 43146 96796 43148
rect 96740 43094 96742 43146
rect 96742 43094 96794 43146
rect 96794 43094 96796 43146
rect 96740 43092 96796 43094
rect 96844 43146 96900 43148
rect 96844 43094 96846 43146
rect 96846 43094 96898 43146
rect 96898 43094 96900 43146
rect 96844 43092 96900 43094
rect 96636 41578 96692 41580
rect 96636 41526 96638 41578
rect 96638 41526 96690 41578
rect 96690 41526 96692 41578
rect 96636 41524 96692 41526
rect 96740 41578 96796 41580
rect 96740 41526 96742 41578
rect 96742 41526 96794 41578
rect 96794 41526 96796 41578
rect 96740 41524 96796 41526
rect 96844 41578 96900 41580
rect 96844 41526 96846 41578
rect 96846 41526 96898 41578
rect 96898 41526 96900 41578
rect 96844 41524 96900 41526
rect 96636 40010 96692 40012
rect 96636 39958 96638 40010
rect 96638 39958 96690 40010
rect 96690 39958 96692 40010
rect 96636 39956 96692 39958
rect 96740 40010 96796 40012
rect 96740 39958 96742 40010
rect 96742 39958 96794 40010
rect 96794 39958 96796 40010
rect 96740 39956 96796 39958
rect 96844 40010 96900 40012
rect 96844 39958 96846 40010
rect 96846 39958 96898 40010
rect 96898 39958 96900 40010
rect 96844 39956 96900 39958
rect 96636 38442 96692 38444
rect 96636 38390 96638 38442
rect 96638 38390 96690 38442
rect 96690 38390 96692 38442
rect 96636 38388 96692 38390
rect 96740 38442 96796 38444
rect 96740 38390 96742 38442
rect 96742 38390 96794 38442
rect 96794 38390 96796 38442
rect 96740 38388 96796 38390
rect 96844 38442 96900 38444
rect 96844 38390 96846 38442
rect 96846 38390 96898 38442
rect 96898 38390 96900 38442
rect 96844 38388 96900 38390
rect 96636 36874 96692 36876
rect 96636 36822 96638 36874
rect 96638 36822 96690 36874
rect 96690 36822 96692 36874
rect 96636 36820 96692 36822
rect 96740 36874 96796 36876
rect 96740 36822 96742 36874
rect 96742 36822 96794 36874
rect 96794 36822 96796 36874
rect 96740 36820 96796 36822
rect 96844 36874 96900 36876
rect 96844 36822 96846 36874
rect 96846 36822 96898 36874
rect 96898 36822 96900 36874
rect 96844 36820 96900 36822
rect 96636 35306 96692 35308
rect 96636 35254 96638 35306
rect 96638 35254 96690 35306
rect 96690 35254 96692 35306
rect 96636 35252 96692 35254
rect 96740 35306 96796 35308
rect 96740 35254 96742 35306
rect 96742 35254 96794 35306
rect 96794 35254 96796 35306
rect 96740 35252 96796 35254
rect 96844 35306 96900 35308
rect 96844 35254 96846 35306
rect 96846 35254 96898 35306
rect 96898 35254 96900 35306
rect 96844 35252 96900 35254
rect 96636 33738 96692 33740
rect 96636 33686 96638 33738
rect 96638 33686 96690 33738
rect 96690 33686 96692 33738
rect 96636 33684 96692 33686
rect 96740 33738 96796 33740
rect 96740 33686 96742 33738
rect 96742 33686 96794 33738
rect 96794 33686 96796 33738
rect 96740 33684 96796 33686
rect 96844 33738 96900 33740
rect 96844 33686 96846 33738
rect 96846 33686 96898 33738
rect 96898 33686 96900 33738
rect 96844 33684 96900 33686
rect 96636 32170 96692 32172
rect 96636 32118 96638 32170
rect 96638 32118 96690 32170
rect 96690 32118 96692 32170
rect 96636 32116 96692 32118
rect 96740 32170 96796 32172
rect 96740 32118 96742 32170
rect 96742 32118 96794 32170
rect 96794 32118 96796 32170
rect 96740 32116 96796 32118
rect 96844 32170 96900 32172
rect 96844 32118 96846 32170
rect 96846 32118 96898 32170
rect 96898 32118 96900 32170
rect 96844 32116 96900 32118
rect 96636 30602 96692 30604
rect 96636 30550 96638 30602
rect 96638 30550 96690 30602
rect 96690 30550 96692 30602
rect 96636 30548 96692 30550
rect 96740 30602 96796 30604
rect 96740 30550 96742 30602
rect 96742 30550 96794 30602
rect 96794 30550 96796 30602
rect 96740 30548 96796 30550
rect 96844 30602 96900 30604
rect 96844 30550 96846 30602
rect 96846 30550 96898 30602
rect 96898 30550 96900 30602
rect 96844 30548 96900 30550
rect 96636 29034 96692 29036
rect 96636 28982 96638 29034
rect 96638 28982 96690 29034
rect 96690 28982 96692 29034
rect 96636 28980 96692 28982
rect 96740 29034 96796 29036
rect 96740 28982 96742 29034
rect 96742 28982 96794 29034
rect 96794 28982 96796 29034
rect 96740 28980 96796 28982
rect 96844 29034 96900 29036
rect 96844 28982 96846 29034
rect 96846 28982 96898 29034
rect 96898 28982 96900 29034
rect 96844 28980 96900 28982
rect 96636 27466 96692 27468
rect 96636 27414 96638 27466
rect 96638 27414 96690 27466
rect 96690 27414 96692 27466
rect 96636 27412 96692 27414
rect 96740 27466 96796 27468
rect 96740 27414 96742 27466
rect 96742 27414 96794 27466
rect 96794 27414 96796 27466
rect 96740 27412 96796 27414
rect 96844 27466 96900 27468
rect 96844 27414 96846 27466
rect 96846 27414 96898 27466
rect 96898 27414 96900 27466
rect 96844 27412 96900 27414
rect 96636 25898 96692 25900
rect 96636 25846 96638 25898
rect 96638 25846 96690 25898
rect 96690 25846 96692 25898
rect 96636 25844 96692 25846
rect 96740 25898 96796 25900
rect 96740 25846 96742 25898
rect 96742 25846 96794 25898
rect 96794 25846 96796 25898
rect 96740 25844 96796 25846
rect 96844 25898 96900 25900
rect 96844 25846 96846 25898
rect 96846 25846 96898 25898
rect 96898 25846 96900 25898
rect 96844 25844 96900 25846
rect 96636 24330 96692 24332
rect 96636 24278 96638 24330
rect 96638 24278 96690 24330
rect 96690 24278 96692 24330
rect 96636 24276 96692 24278
rect 96740 24330 96796 24332
rect 96740 24278 96742 24330
rect 96742 24278 96794 24330
rect 96794 24278 96796 24330
rect 96740 24276 96796 24278
rect 96844 24330 96900 24332
rect 96844 24278 96846 24330
rect 96846 24278 96898 24330
rect 96898 24278 96900 24330
rect 96844 24276 96900 24278
rect 96636 22762 96692 22764
rect 96636 22710 96638 22762
rect 96638 22710 96690 22762
rect 96690 22710 96692 22762
rect 96636 22708 96692 22710
rect 96740 22762 96796 22764
rect 96740 22710 96742 22762
rect 96742 22710 96794 22762
rect 96794 22710 96796 22762
rect 96740 22708 96796 22710
rect 96844 22762 96900 22764
rect 96844 22710 96846 22762
rect 96846 22710 96898 22762
rect 96898 22710 96900 22762
rect 96844 22708 96900 22710
rect 96636 21194 96692 21196
rect 96636 21142 96638 21194
rect 96638 21142 96690 21194
rect 96690 21142 96692 21194
rect 96636 21140 96692 21142
rect 96740 21194 96796 21196
rect 96740 21142 96742 21194
rect 96742 21142 96794 21194
rect 96794 21142 96796 21194
rect 96740 21140 96796 21142
rect 96844 21194 96900 21196
rect 96844 21142 96846 21194
rect 96846 21142 96898 21194
rect 96898 21142 96900 21194
rect 96844 21140 96900 21142
rect 92428 20972 92484 21028
rect 96636 19626 96692 19628
rect 96636 19574 96638 19626
rect 96638 19574 96690 19626
rect 96690 19574 96692 19626
rect 96636 19572 96692 19574
rect 96740 19626 96796 19628
rect 96740 19574 96742 19626
rect 96742 19574 96794 19626
rect 96794 19574 96796 19626
rect 96740 19572 96796 19574
rect 96844 19626 96900 19628
rect 96844 19574 96846 19626
rect 96846 19574 96898 19626
rect 96898 19574 96900 19626
rect 96844 19572 96900 19574
rect 96636 18058 96692 18060
rect 96636 18006 96638 18058
rect 96638 18006 96690 18058
rect 96690 18006 96692 18058
rect 96636 18004 96692 18006
rect 96740 18058 96796 18060
rect 96740 18006 96742 18058
rect 96742 18006 96794 18058
rect 96794 18006 96796 18058
rect 96740 18004 96796 18006
rect 96844 18058 96900 18060
rect 96844 18006 96846 18058
rect 96846 18006 96898 18058
rect 96898 18006 96900 18058
rect 96844 18004 96900 18006
rect 96636 16490 96692 16492
rect 96636 16438 96638 16490
rect 96638 16438 96690 16490
rect 96690 16438 96692 16490
rect 96636 16436 96692 16438
rect 96740 16490 96796 16492
rect 96740 16438 96742 16490
rect 96742 16438 96794 16490
rect 96794 16438 96796 16490
rect 96740 16436 96796 16438
rect 96844 16490 96900 16492
rect 96844 16438 96846 16490
rect 96846 16438 96898 16490
rect 96898 16438 96900 16490
rect 96844 16436 96900 16438
rect 96636 14922 96692 14924
rect 96636 14870 96638 14922
rect 96638 14870 96690 14922
rect 96690 14870 96692 14922
rect 96636 14868 96692 14870
rect 96740 14922 96796 14924
rect 96740 14870 96742 14922
rect 96742 14870 96794 14922
rect 96794 14870 96796 14922
rect 96740 14868 96796 14870
rect 96844 14922 96900 14924
rect 96844 14870 96846 14922
rect 96846 14870 96898 14922
rect 96898 14870 96900 14922
rect 96844 14868 96900 14870
rect 96636 13354 96692 13356
rect 96636 13302 96638 13354
rect 96638 13302 96690 13354
rect 96690 13302 96692 13354
rect 96636 13300 96692 13302
rect 96740 13354 96796 13356
rect 96740 13302 96742 13354
rect 96742 13302 96794 13354
rect 96794 13302 96796 13354
rect 96740 13300 96796 13302
rect 96844 13354 96900 13356
rect 96844 13302 96846 13354
rect 96846 13302 96898 13354
rect 96898 13302 96900 13354
rect 96844 13300 96900 13302
rect 96636 11786 96692 11788
rect 96636 11734 96638 11786
rect 96638 11734 96690 11786
rect 96690 11734 96692 11786
rect 96636 11732 96692 11734
rect 96740 11786 96796 11788
rect 96740 11734 96742 11786
rect 96742 11734 96794 11786
rect 96794 11734 96796 11786
rect 96740 11732 96796 11734
rect 96844 11786 96900 11788
rect 96844 11734 96846 11786
rect 96846 11734 96898 11786
rect 96898 11734 96900 11786
rect 96844 11732 96900 11734
rect 96636 10218 96692 10220
rect 96636 10166 96638 10218
rect 96638 10166 96690 10218
rect 96690 10166 96692 10218
rect 96636 10164 96692 10166
rect 96740 10218 96796 10220
rect 96740 10166 96742 10218
rect 96742 10166 96794 10218
rect 96794 10166 96796 10218
rect 96740 10164 96796 10166
rect 96844 10218 96900 10220
rect 96844 10166 96846 10218
rect 96846 10166 96898 10218
rect 96898 10166 96900 10218
rect 96844 10164 96900 10166
rect 100044 55410 100100 55412
rect 100044 55358 100046 55410
rect 100046 55358 100098 55410
rect 100098 55358 100100 55410
rect 100044 55356 100100 55358
rect 102508 49532 102564 49588
rect 110348 55132 110404 55188
rect 111996 54906 112052 54908
rect 111996 54854 111998 54906
rect 111998 54854 112050 54906
rect 112050 54854 112052 54906
rect 111996 54852 112052 54854
rect 112100 54906 112156 54908
rect 112100 54854 112102 54906
rect 112102 54854 112154 54906
rect 112154 54854 112156 54906
rect 112100 54852 112156 54854
rect 112204 54906 112260 54908
rect 112204 54854 112206 54906
rect 112206 54854 112258 54906
rect 112258 54854 112260 54906
rect 112204 54852 112260 54854
rect 111996 53338 112052 53340
rect 111996 53286 111998 53338
rect 111998 53286 112050 53338
rect 112050 53286 112052 53338
rect 111996 53284 112052 53286
rect 112100 53338 112156 53340
rect 112100 53286 112102 53338
rect 112102 53286 112154 53338
rect 112154 53286 112156 53338
rect 112100 53284 112156 53286
rect 112204 53338 112260 53340
rect 112204 53286 112206 53338
rect 112206 53286 112258 53338
rect 112258 53286 112260 53338
rect 112204 53284 112260 53286
rect 121100 55970 121156 55972
rect 121100 55918 121102 55970
rect 121102 55918 121154 55970
rect 121154 55918 121156 55970
rect 121100 55916 121156 55918
rect 127356 55690 127412 55692
rect 127356 55638 127358 55690
rect 127358 55638 127410 55690
rect 127410 55638 127412 55690
rect 127356 55636 127412 55638
rect 127460 55690 127516 55692
rect 127460 55638 127462 55690
rect 127462 55638 127514 55690
rect 127514 55638 127516 55690
rect 127460 55636 127516 55638
rect 127564 55690 127620 55692
rect 127564 55638 127566 55690
rect 127566 55638 127618 55690
rect 127618 55638 127620 55690
rect 127564 55636 127620 55638
rect 127356 54122 127412 54124
rect 127356 54070 127358 54122
rect 127358 54070 127410 54122
rect 127410 54070 127412 54122
rect 127356 54068 127412 54070
rect 127460 54122 127516 54124
rect 127460 54070 127462 54122
rect 127462 54070 127514 54122
rect 127514 54070 127516 54122
rect 127460 54068 127516 54070
rect 127564 54122 127620 54124
rect 127564 54070 127566 54122
rect 127566 54070 127618 54122
rect 127618 54070 127620 54122
rect 127564 54068 127620 54070
rect 135772 56140 135828 56196
rect 130284 54348 130340 54404
rect 132972 55244 133028 55300
rect 135100 55298 135156 55300
rect 135100 55246 135102 55298
rect 135102 55246 135154 55298
rect 135154 55246 135156 55298
rect 135100 55244 135156 55246
rect 136668 56194 136724 56196
rect 136668 56142 136670 56194
rect 136670 56142 136722 56194
rect 136722 56142 136724 56194
rect 136668 56140 136724 56142
rect 142716 56474 142772 56476
rect 142716 56422 142718 56474
rect 142718 56422 142770 56474
rect 142770 56422 142772 56474
rect 142716 56420 142772 56422
rect 142820 56474 142876 56476
rect 142820 56422 142822 56474
rect 142822 56422 142874 56474
rect 142874 56422 142876 56474
rect 142820 56420 142876 56422
rect 142924 56474 142980 56476
rect 142924 56422 142926 56474
rect 142926 56422 142978 56474
rect 142978 56422 142980 56474
rect 142924 56420 142980 56422
rect 142156 56140 142212 56196
rect 141260 55410 141316 55412
rect 141260 55358 141262 55410
rect 141262 55358 141314 55410
rect 141314 55358 141316 55410
rect 141260 55356 141316 55358
rect 138348 55298 138404 55300
rect 138348 55246 138350 55298
rect 138350 55246 138402 55298
rect 138402 55246 138404 55298
rect 138348 55244 138404 55246
rect 140476 55298 140532 55300
rect 140476 55246 140478 55298
rect 140478 55246 140530 55298
rect 140530 55246 140532 55298
rect 140476 55244 140532 55246
rect 142828 56140 142884 56196
rect 142604 55356 142660 55412
rect 143836 55298 143892 55300
rect 143836 55246 143838 55298
rect 143838 55246 143890 55298
rect 143890 55246 143892 55298
rect 143836 55244 143892 55246
rect 142716 54906 142772 54908
rect 142716 54854 142718 54906
rect 142718 54854 142770 54906
rect 142770 54854 142772 54906
rect 142716 54852 142772 54854
rect 142820 54906 142876 54908
rect 142820 54854 142822 54906
rect 142822 54854 142874 54906
rect 142874 54854 142876 54906
rect 142820 54852 142876 54854
rect 142924 54906 142980 54908
rect 142924 54854 142926 54906
rect 142926 54854 142978 54906
rect 142978 54854 142980 54906
rect 142924 54852 142980 54854
rect 131740 54402 131796 54404
rect 131740 54350 131742 54402
rect 131742 54350 131794 54402
rect 131794 54350 131796 54402
rect 131740 54348 131796 54350
rect 145964 54348 146020 54404
rect 127820 52780 127876 52836
rect 127356 52554 127412 52556
rect 127356 52502 127358 52554
rect 127358 52502 127410 52554
rect 127410 52502 127412 52554
rect 127356 52500 127412 52502
rect 127460 52554 127516 52556
rect 127460 52502 127462 52554
rect 127462 52502 127514 52554
rect 127514 52502 127516 52554
rect 127460 52500 127516 52502
rect 127564 52554 127620 52556
rect 127564 52502 127566 52554
rect 127566 52502 127618 52554
rect 127618 52502 127620 52554
rect 127564 52500 127620 52502
rect 116508 52108 116564 52164
rect 111996 51770 112052 51772
rect 111996 51718 111998 51770
rect 111998 51718 112050 51770
rect 112050 51718 112052 51770
rect 111996 51716 112052 51718
rect 112100 51770 112156 51772
rect 112100 51718 112102 51770
rect 112102 51718 112154 51770
rect 112154 51718 112156 51770
rect 112100 51716 112156 51718
rect 112204 51770 112260 51772
rect 112204 51718 112206 51770
rect 112206 51718 112258 51770
rect 112258 51718 112260 51770
rect 112204 51716 112260 51718
rect 127356 50986 127412 50988
rect 127356 50934 127358 50986
rect 127358 50934 127410 50986
rect 127410 50934 127412 50986
rect 127356 50932 127412 50934
rect 127460 50986 127516 50988
rect 127460 50934 127462 50986
rect 127462 50934 127514 50986
rect 127514 50934 127516 50986
rect 127460 50932 127516 50934
rect 127564 50986 127620 50988
rect 127564 50934 127566 50986
rect 127566 50934 127618 50986
rect 127618 50934 127620 50986
rect 127564 50932 127620 50934
rect 111996 50202 112052 50204
rect 111996 50150 111998 50202
rect 111998 50150 112050 50202
rect 112050 50150 112052 50202
rect 111996 50148 112052 50150
rect 112100 50202 112156 50204
rect 112100 50150 112102 50202
rect 112102 50150 112154 50202
rect 112154 50150 112156 50202
rect 112100 50148 112156 50150
rect 112204 50202 112260 50204
rect 112204 50150 112206 50202
rect 112206 50150 112258 50202
rect 112258 50150 112260 50202
rect 112204 50148 112260 50150
rect 127356 49418 127412 49420
rect 127356 49366 127358 49418
rect 127358 49366 127410 49418
rect 127410 49366 127412 49418
rect 127356 49364 127412 49366
rect 127460 49418 127516 49420
rect 127460 49366 127462 49418
rect 127462 49366 127514 49418
rect 127514 49366 127516 49418
rect 127460 49364 127516 49366
rect 127564 49418 127620 49420
rect 127564 49366 127566 49418
rect 127566 49366 127618 49418
rect 127618 49366 127620 49418
rect 127564 49364 127620 49366
rect 111996 48634 112052 48636
rect 111996 48582 111998 48634
rect 111998 48582 112050 48634
rect 112050 48582 112052 48634
rect 111996 48580 112052 48582
rect 112100 48634 112156 48636
rect 112100 48582 112102 48634
rect 112102 48582 112154 48634
rect 112154 48582 112156 48634
rect 112100 48580 112156 48582
rect 112204 48634 112260 48636
rect 112204 48582 112206 48634
rect 112206 48582 112258 48634
rect 112258 48582 112260 48634
rect 112204 48580 112260 48582
rect 127356 47850 127412 47852
rect 127356 47798 127358 47850
rect 127358 47798 127410 47850
rect 127410 47798 127412 47850
rect 127356 47796 127412 47798
rect 127460 47850 127516 47852
rect 127460 47798 127462 47850
rect 127462 47798 127514 47850
rect 127514 47798 127516 47850
rect 127460 47796 127516 47798
rect 127564 47850 127620 47852
rect 127564 47798 127566 47850
rect 127566 47798 127618 47850
rect 127618 47798 127620 47850
rect 127564 47796 127620 47798
rect 111996 47066 112052 47068
rect 111996 47014 111998 47066
rect 111998 47014 112050 47066
rect 112050 47014 112052 47066
rect 111996 47012 112052 47014
rect 112100 47066 112156 47068
rect 112100 47014 112102 47066
rect 112102 47014 112154 47066
rect 112154 47014 112156 47066
rect 112100 47012 112156 47014
rect 112204 47066 112260 47068
rect 112204 47014 112206 47066
rect 112206 47014 112258 47066
rect 112258 47014 112260 47066
rect 112204 47012 112260 47014
rect 127356 46282 127412 46284
rect 127356 46230 127358 46282
rect 127358 46230 127410 46282
rect 127410 46230 127412 46282
rect 127356 46228 127412 46230
rect 127460 46282 127516 46284
rect 127460 46230 127462 46282
rect 127462 46230 127514 46282
rect 127514 46230 127516 46282
rect 127460 46228 127516 46230
rect 127564 46282 127620 46284
rect 127564 46230 127566 46282
rect 127566 46230 127618 46282
rect 127618 46230 127620 46282
rect 127564 46228 127620 46230
rect 111996 45498 112052 45500
rect 111996 45446 111998 45498
rect 111998 45446 112050 45498
rect 112050 45446 112052 45498
rect 111996 45444 112052 45446
rect 112100 45498 112156 45500
rect 112100 45446 112102 45498
rect 112102 45446 112154 45498
rect 112154 45446 112156 45498
rect 112100 45444 112156 45446
rect 112204 45498 112260 45500
rect 112204 45446 112206 45498
rect 112206 45446 112258 45498
rect 112258 45446 112260 45498
rect 112204 45444 112260 45446
rect 127356 44714 127412 44716
rect 127356 44662 127358 44714
rect 127358 44662 127410 44714
rect 127410 44662 127412 44714
rect 127356 44660 127412 44662
rect 127460 44714 127516 44716
rect 127460 44662 127462 44714
rect 127462 44662 127514 44714
rect 127514 44662 127516 44714
rect 127460 44660 127516 44662
rect 127564 44714 127620 44716
rect 127564 44662 127566 44714
rect 127566 44662 127618 44714
rect 127618 44662 127620 44714
rect 127564 44660 127620 44662
rect 111996 43930 112052 43932
rect 111996 43878 111998 43930
rect 111998 43878 112050 43930
rect 112050 43878 112052 43930
rect 111996 43876 112052 43878
rect 112100 43930 112156 43932
rect 112100 43878 112102 43930
rect 112102 43878 112154 43930
rect 112154 43878 112156 43930
rect 112100 43876 112156 43878
rect 112204 43930 112260 43932
rect 112204 43878 112206 43930
rect 112206 43878 112258 43930
rect 112258 43878 112260 43930
rect 112204 43876 112260 43878
rect 127356 43146 127412 43148
rect 127356 43094 127358 43146
rect 127358 43094 127410 43146
rect 127410 43094 127412 43146
rect 127356 43092 127412 43094
rect 127460 43146 127516 43148
rect 127460 43094 127462 43146
rect 127462 43094 127514 43146
rect 127514 43094 127516 43146
rect 127460 43092 127516 43094
rect 127564 43146 127620 43148
rect 127564 43094 127566 43146
rect 127566 43094 127618 43146
rect 127618 43094 127620 43146
rect 127564 43092 127620 43094
rect 111996 42362 112052 42364
rect 111996 42310 111998 42362
rect 111998 42310 112050 42362
rect 112050 42310 112052 42362
rect 111996 42308 112052 42310
rect 112100 42362 112156 42364
rect 112100 42310 112102 42362
rect 112102 42310 112154 42362
rect 112154 42310 112156 42362
rect 112100 42308 112156 42310
rect 112204 42362 112260 42364
rect 112204 42310 112206 42362
rect 112206 42310 112258 42362
rect 112258 42310 112260 42362
rect 112204 42308 112260 42310
rect 127356 41578 127412 41580
rect 127356 41526 127358 41578
rect 127358 41526 127410 41578
rect 127410 41526 127412 41578
rect 127356 41524 127412 41526
rect 127460 41578 127516 41580
rect 127460 41526 127462 41578
rect 127462 41526 127514 41578
rect 127514 41526 127516 41578
rect 127460 41524 127516 41526
rect 127564 41578 127620 41580
rect 127564 41526 127566 41578
rect 127566 41526 127618 41578
rect 127618 41526 127620 41578
rect 127564 41524 127620 41526
rect 111996 40794 112052 40796
rect 111996 40742 111998 40794
rect 111998 40742 112050 40794
rect 112050 40742 112052 40794
rect 111996 40740 112052 40742
rect 112100 40794 112156 40796
rect 112100 40742 112102 40794
rect 112102 40742 112154 40794
rect 112154 40742 112156 40794
rect 112100 40740 112156 40742
rect 112204 40794 112260 40796
rect 112204 40742 112206 40794
rect 112206 40742 112258 40794
rect 112258 40742 112260 40794
rect 112204 40740 112260 40742
rect 127356 40010 127412 40012
rect 127356 39958 127358 40010
rect 127358 39958 127410 40010
rect 127410 39958 127412 40010
rect 127356 39956 127412 39958
rect 127460 40010 127516 40012
rect 127460 39958 127462 40010
rect 127462 39958 127514 40010
rect 127514 39958 127516 40010
rect 127460 39956 127516 39958
rect 127564 40010 127620 40012
rect 127564 39958 127566 40010
rect 127566 39958 127618 40010
rect 127618 39958 127620 40010
rect 127564 39956 127620 39958
rect 111996 39226 112052 39228
rect 111996 39174 111998 39226
rect 111998 39174 112050 39226
rect 112050 39174 112052 39226
rect 111996 39172 112052 39174
rect 112100 39226 112156 39228
rect 112100 39174 112102 39226
rect 112102 39174 112154 39226
rect 112154 39174 112156 39226
rect 112100 39172 112156 39174
rect 112204 39226 112260 39228
rect 112204 39174 112206 39226
rect 112206 39174 112258 39226
rect 112258 39174 112260 39226
rect 112204 39172 112260 39174
rect 127356 38442 127412 38444
rect 127356 38390 127358 38442
rect 127358 38390 127410 38442
rect 127410 38390 127412 38442
rect 127356 38388 127412 38390
rect 127460 38442 127516 38444
rect 127460 38390 127462 38442
rect 127462 38390 127514 38442
rect 127514 38390 127516 38442
rect 127460 38388 127516 38390
rect 127564 38442 127620 38444
rect 127564 38390 127566 38442
rect 127566 38390 127618 38442
rect 127618 38390 127620 38442
rect 127564 38388 127620 38390
rect 111996 37658 112052 37660
rect 111996 37606 111998 37658
rect 111998 37606 112050 37658
rect 112050 37606 112052 37658
rect 111996 37604 112052 37606
rect 112100 37658 112156 37660
rect 112100 37606 112102 37658
rect 112102 37606 112154 37658
rect 112154 37606 112156 37658
rect 112100 37604 112156 37606
rect 112204 37658 112260 37660
rect 112204 37606 112206 37658
rect 112206 37606 112258 37658
rect 112258 37606 112260 37658
rect 112204 37604 112260 37606
rect 127356 36874 127412 36876
rect 127356 36822 127358 36874
rect 127358 36822 127410 36874
rect 127410 36822 127412 36874
rect 127356 36820 127412 36822
rect 127460 36874 127516 36876
rect 127460 36822 127462 36874
rect 127462 36822 127514 36874
rect 127514 36822 127516 36874
rect 127460 36820 127516 36822
rect 127564 36874 127620 36876
rect 127564 36822 127566 36874
rect 127566 36822 127618 36874
rect 127618 36822 127620 36874
rect 127564 36820 127620 36822
rect 111996 36090 112052 36092
rect 111996 36038 111998 36090
rect 111998 36038 112050 36090
rect 112050 36038 112052 36090
rect 111996 36036 112052 36038
rect 112100 36090 112156 36092
rect 112100 36038 112102 36090
rect 112102 36038 112154 36090
rect 112154 36038 112156 36090
rect 112100 36036 112156 36038
rect 112204 36090 112260 36092
rect 112204 36038 112206 36090
rect 112206 36038 112258 36090
rect 112258 36038 112260 36090
rect 112204 36036 112260 36038
rect 127356 35306 127412 35308
rect 127356 35254 127358 35306
rect 127358 35254 127410 35306
rect 127410 35254 127412 35306
rect 127356 35252 127412 35254
rect 127460 35306 127516 35308
rect 127460 35254 127462 35306
rect 127462 35254 127514 35306
rect 127514 35254 127516 35306
rect 127460 35252 127516 35254
rect 127564 35306 127620 35308
rect 127564 35254 127566 35306
rect 127566 35254 127618 35306
rect 127618 35254 127620 35306
rect 127564 35252 127620 35254
rect 111996 34522 112052 34524
rect 111996 34470 111998 34522
rect 111998 34470 112050 34522
rect 112050 34470 112052 34522
rect 111996 34468 112052 34470
rect 112100 34522 112156 34524
rect 112100 34470 112102 34522
rect 112102 34470 112154 34522
rect 112154 34470 112156 34522
rect 112100 34468 112156 34470
rect 112204 34522 112260 34524
rect 112204 34470 112206 34522
rect 112206 34470 112258 34522
rect 112258 34470 112260 34522
rect 112204 34468 112260 34470
rect 127356 33738 127412 33740
rect 127356 33686 127358 33738
rect 127358 33686 127410 33738
rect 127410 33686 127412 33738
rect 127356 33684 127412 33686
rect 127460 33738 127516 33740
rect 127460 33686 127462 33738
rect 127462 33686 127514 33738
rect 127514 33686 127516 33738
rect 127460 33684 127516 33686
rect 127564 33738 127620 33740
rect 127564 33686 127566 33738
rect 127566 33686 127618 33738
rect 127618 33686 127620 33738
rect 127564 33684 127620 33686
rect 111996 32954 112052 32956
rect 111996 32902 111998 32954
rect 111998 32902 112050 32954
rect 112050 32902 112052 32954
rect 111996 32900 112052 32902
rect 112100 32954 112156 32956
rect 112100 32902 112102 32954
rect 112102 32902 112154 32954
rect 112154 32902 112156 32954
rect 112100 32900 112156 32902
rect 112204 32954 112260 32956
rect 112204 32902 112206 32954
rect 112206 32902 112258 32954
rect 112258 32902 112260 32954
rect 112204 32900 112260 32902
rect 127356 32170 127412 32172
rect 127356 32118 127358 32170
rect 127358 32118 127410 32170
rect 127410 32118 127412 32170
rect 127356 32116 127412 32118
rect 127460 32170 127516 32172
rect 127460 32118 127462 32170
rect 127462 32118 127514 32170
rect 127514 32118 127516 32170
rect 127460 32116 127516 32118
rect 127564 32170 127620 32172
rect 127564 32118 127566 32170
rect 127566 32118 127618 32170
rect 127618 32118 127620 32170
rect 127564 32116 127620 32118
rect 111996 31386 112052 31388
rect 111996 31334 111998 31386
rect 111998 31334 112050 31386
rect 112050 31334 112052 31386
rect 111996 31332 112052 31334
rect 112100 31386 112156 31388
rect 112100 31334 112102 31386
rect 112102 31334 112154 31386
rect 112154 31334 112156 31386
rect 112100 31332 112156 31334
rect 112204 31386 112260 31388
rect 112204 31334 112206 31386
rect 112206 31334 112258 31386
rect 112258 31334 112260 31386
rect 112204 31332 112260 31334
rect 127356 30602 127412 30604
rect 127356 30550 127358 30602
rect 127358 30550 127410 30602
rect 127410 30550 127412 30602
rect 127356 30548 127412 30550
rect 127460 30602 127516 30604
rect 127460 30550 127462 30602
rect 127462 30550 127514 30602
rect 127514 30550 127516 30602
rect 127460 30548 127516 30550
rect 127564 30602 127620 30604
rect 127564 30550 127566 30602
rect 127566 30550 127618 30602
rect 127618 30550 127620 30602
rect 127564 30548 127620 30550
rect 111996 29818 112052 29820
rect 111996 29766 111998 29818
rect 111998 29766 112050 29818
rect 112050 29766 112052 29818
rect 111996 29764 112052 29766
rect 112100 29818 112156 29820
rect 112100 29766 112102 29818
rect 112102 29766 112154 29818
rect 112154 29766 112156 29818
rect 112100 29764 112156 29766
rect 112204 29818 112260 29820
rect 112204 29766 112206 29818
rect 112206 29766 112258 29818
rect 112258 29766 112260 29818
rect 112204 29764 112260 29766
rect 127356 29034 127412 29036
rect 127356 28982 127358 29034
rect 127358 28982 127410 29034
rect 127410 28982 127412 29034
rect 127356 28980 127412 28982
rect 127460 29034 127516 29036
rect 127460 28982 127462 29034
rect 127462 28982 127514 29034
rect 127514 28982 127516 29034
rect 127460 28980 127516 28982
rect 127564 29034 127620 29036
rect 127564 28982 127566 29034
rect 127566 28982 127618 29034
rect 127618 28982 127620 29034
rect 127564 28980 127620 28982
rect 111996 28250 112052 28252
rect 111996 28198 111998 28250
rect 111998 28198 112050 28250
rect 112050 28198 112052 28250
rect 111996 28196 112052 28198
rect 112100 28250 112156 28252
rect 112100 28198 112102 28250
rect 112102 28198 112154 28250
rect 112154 28198 112156 28250
rect 112100 28196 112156 28198
rect 112204 28250 112260 28252
rect 112204 28198 112206 28250
rect 112206 28198 112258 28250
rect 112258 28198 112260 28250
rect 112204 28196 112260 28198
rect 127356 27466 127412 27468
rect 127356 27414 127358 27466
rect 127358 27414 127410 27466
rect 127410 27414 127412 27466
rect 127356 27412 127412 27414
rect 127460 27466 127516 27468
rect 127460 27414 127462 27466
rect 127462 27414 127514 27466
rect 127514 27414 127516 27466
rect 127460 27412 127516 27414
rect 127564 27466 127620 27468
rect 127564 27414 127566 27466
rect 127566 27414 127618 27466
rect 127618 27414 127620 27466
rect 127564 27412 127620 27414
rect 111996 26682 112052 26684
rect 111996 26630 111998 26682
rect 111998 26630 112050 26682
rect 112050 26630 112052 26682
rect 111996 26628 112052 26630
rect 112100 26682 112156 26684
rect 112100 26630 112102 26682
rect 112102 26630 112154 26682
rect 112154 26630 112156 26682
rect 112100 26628 112156 26630
rect 112204 26682 112260 26684
rect 112204 26630 112206 26682
rect 112206 26630 112258 26682
rect 112258 26630 112260 26682
rect 112204 26628 112260 26630
rect 127356 25898 127412 25900
rect 127356 25846 127358 25898
rect 127358 25846 127410 25898
rect 127410 25846 127412 25898
rect 127356 25844 127412 25846
rect 127460 25898 127516 25900
rect 127460 25846 127462 25898
rect 127462 25846 127514 25898
rect 127514 25846 127516 25898
rect 127460 25844 127516 25846
rect 127564 25898 127620 25900
rect 127564 25846 127566 25898
rect 127566 25846 127618 25898
rect 127618 25846 127620 25898
rect 127564 25844 127620 25846
rect 111996 25114 112052 25116
rect 111996 25062 111998 25114
rect 111998 25062 112050 25114
rect 112050 25062 112052 25114
rect 111996 25060 112052 25062
rect 112100 25114 112156 25116
rect 112100 25062 112102 25114
rect 112102 25062 112154 25114
rect 112154 25062 112156 25114
rect 112100 25060 112156 25062
rect 112204 25114 112260 25116
rect 112204 25062 112206 25114
rect 112206 25062 112258 25114
rect 112258 25062 112260 25114
rect 112204 25060 112260 25062
rect 147868 55244 147924 55300
rect 152684 55020 152740 55076
rect 148092 54684 148148 54740
rect 148652 54738 148708 54740
rect 148652 54686 148654 54738
rect 148654 54686 148706 54738
rect 148706 54686 148708 54738
rect 148652 54684 148708 54686
rect 150108 54738 150164 54740
rect 150108 54686 150110 54738
rect 150110 54686 150162 54738
rect 150162 54686 150164 54738
rect 150108 54684 150164 54686
rect 147420 54402 147476 54404
rect 147420 54350 147422 54402
rect 147422 54350 147474 54402
rect 147474 54350 147476 54402
rect 147420 54348 147476 54350
rect 151564 54348 151620 54404
rect 158076 55690 158132 55692
rect 158076 55638 158078 55690
rect 158078 55638 158130 55690
rect 158130 55638 158132 55690
rect 158076 55636 158132 55638
rect 158180 55690 158236 55692
rect 158180 55638 158182 55690
rect 158182 55638 158234 55690
rect 158234 55638 158236 55690
rect 158180 55636 158236 55638
rect 158284 55690 158340 55692
rect 158284 55638 158286 55690
rect 158286 55638 158338 55690
rect 158338 55638 158340 55690
rect 158284 55636 158340 55638
rect 173436 56474 173492 56476
rect 173436 56422 173438 56474
rect 173438 56422 173490 56474
rect 173490 56422 173492 56474
rect 173436 56420 173492 56422
rect 173540 56474 173596 56476
rect 173540 56422 173542 56474
rect 173542 56422 173594 56474
rect 173594 56422 173596 56474
rect 173540 56420 173596 56422
rect 173644 56474 173700 56476
rect 173644 56422 173646 56474
rect 173646 56422 173698 56474
rect 173698 56422 173700 56474
rect 173644 56420 173700 56422
rect 153916 55356 153972 55412
rect 153244 55074 153300 55076
rect 153244 55022 153246 55074
rect 153246 55022 153298 55074
rect 153298 55022 153300 55074
rect 153244 55020 153300 55022
rect 156268 55410 156324 55412
rect 156268 55358 156270 55410
rect 156270 55358 156322 55410
rect 156322 55358 156324 55410
rect 156268 55356 156324 55358
rect 156716 55356 156772 55412
rect 161868 55410 161924 55412
rect 161868 55358 161870 55410
rect 161870 55358 161922 55410
rect 161922 55358 161924 55410
rect 161868 55356 161924 55358
rect 162428 55356 162484 55412
rect 153916 54684 153972 54740
rect 162316 54738 162372 54740
rect 162316 54686 162318 54738
rect 162318 54686 162370 54738
rect 162370 54686 162372 54738
rect 162316 54684 162372 54686
rect 169708 55298 169764 55300
rect 169708 55246 169710 55298
rect 169710 55246 169762 55298
rect 169762 55246 169764 55298
rect 169708 55244 169764 55246
rect 170380 55298 170436 55300
rect 170380 55246 170382 55298
rect 170382 55246 170434 55298
rect 170434 55246 170436 55298
rect 170380 55244 170436 55246
rect 163212 54684 163268 54740
rect 166236 55020 166292 55076
rect 153132 54402 153188 54404
rect 153132 54350 153134 54402
rect 153134 54350 153186 54402
rect 153186 54350 153188 54402
rect 153132 54348 153188 54350
rect 142716 53338 142772 53340
rect 142716 53286 142718 53338
rect 142718 53286 142770 53338
rect 142770 53286 142772 53338
rect 142716 53284 142772 53286
rect 142820 53338 142876 53340
rect 142820 53286 142822 53338
rect 142822 53286 142874 53338
rect 142874 53286 142876 53338
rect 142820 53284 142876 53286
rect 142924 53338 142980 53340
rect 142924 53286 142926 53338
rect 142926 53286 142978 53338
rect 142978 53286 142980 53338
rect 142924 53284 142980 53286
rect 142716 51770 142772 51772
rect 142716 51718 142718 51770
rect 142718 51718 142770 51770
rect 142770 51718 142772 51770
rect 142716 51716 142772 51718
rect 142820 51770 142876 51772
rect 142820 51718 142822 51770
rect 142822 51718 142874 51770
rect 142874 51718 142876 51770
rect 142820 51716 142876 51718
rect 142924 51770 142980 51772
rect 142924 51718 142926 51770
rect 142926 51718 142978 51770
rect 142978 51718 142980 51770
rect 142924 51716 142980 51718
rect 142716 50202 142772 50204
rect 142716 50150 142718 50202
rect 142718 50150 142770 50202
rect 142770 50150 142772 50202
rect 142716 50148 142772 50150
rect 142820 50202 142876 50204
rect 142820 50150 142822 50202
rect 142822 50150 142874 50202
rect 142874 50150 142876 50202
rect 142820 50148 142876 50150
rect 142924 50202 142980 50204
rect 142924 50150 142926 50202
rect 142926 50150 142978 50202
rect 142978 50150 142980 50202
rect 142924 50148 142980 50150
rect 142716 48634 142772 48636
rect 142716 48582 142718 48634
rect 142718 48582 142770 48634
rect 142770 48582 142772 48634
rect 142716 48580 142772 48582
rect 142820 48634 142876 48636
rect 142820 48582 142822 48634
rect 142822 48582 142874 48634
rect 142874 48582 142876 48634
rect 142820 48580 142876 48582
rect 142924 48634 142980 48636
rect 142924 48582 142926 48634
rect 142926 48582 142978 48634
rect 142978 48582 142980 48634
rect 142924 48580 142980 48582
rect 142716 47066 142772 47068
rect 142716 47014 142718 47066
rect 142718 47014 142770 47066
rect 142770 47014 142772 47066
rect 142716 47012 142772 47014
rect 142820 47066 142876 47068
rect 142820 47014 142822 47066
rect 142822 47014 142874 47066
rect 142874 47014 142876 47066
rect 142820 47012 142876 47014
rect 142924 47066 142980 47068
rect 142924 47014 142926 47066
rect 142926 47014 142978 47066
rect 142978 47014 142980 47066
rect 142924 47012 142980 47014
rect 142716 45498 142772 45500
rect 142716 45446 142718 45498
rect 142718 45446 142770 45498
rect 142770 45446 142772 45498
rect 142716 45444 142772 45446
rect 142820 45498 142876 45500
rect 142820 45446 142822 45498
rect 142822 45446 142874 45498
rect 142874 45446 142876 45498
rect 142820 45444 142876 45446
rect 142924 45498 142980 45500
rect 142924 45446 142926 45498
rect 142926 45446 142978 45498
rect 142978 45446 142980 45498
rect 142924 45444 142980 45446
rect 142716 43930 142772 43932
rect 142716 43878 142718 43930
rect 142718 43878 142770 43930
rect 142770 43878 142772 43930
rect 142716 43876 142772 43878
rect 142820 43930 142876 43932
rect 142820 43878 142822 43930
rect 142822 43878 142874 43930
rect 142874 43878 142876 43930
rect 142820 43876 142876 43878
rect 142924 43930 142980 43932
rect 142924 43878 142926 43930
rect 142926 43878 142978 43930
rect 142978 43878 142980 43930
rect 142924 43876 142980 43878
rect 142716 42362 142772 42364
rect 142716 42310 142718 42362
rect 142718 42310 142770 42362
rect 142770 42310 142772 42362
rect 142716 42308 142772 42310
rect 142820 42362 142876 42364
rect 142820 42310 142822 42362
rect 142822 42310 142874 42362
rect 142874 42310 142876 42362
rect 142820 42308 142876 42310
rect 142924 42362 142980 42364
rect 142924 42310 142926 42362
rect 142926 42310 142978 42362
rect 142978 42310 142980 42362
rect 142924 42308 142980 42310
rect 145180 41132 145236 41188
rect 142716 40794 142772 40796
rect 142716 40742 142718 40794
rect 142718 40742 142770 40794
rect 142770 40742 142772 40794
rect 142716 40740 142772 40742
rect 142820 40794 142876 40796
rect 142820 40742 142822 40794
rect 142822 40742 142874 40794
rect 142874 40742 142876 40794
rect 142820 40740 142876 40742
rect 142924 40794 142980 40796
rect 142924 40742 142926 40794
rect 142926 40742 142978 40794
rect 142978 40742 142980 40794
rect 142924 40740 142980 40742
rect 142716 39226 142772 39228
rect 142716 39174 142718 39226
rect 142718 39174 142770 39226
rect 142770 39174 142772 39226
rect 142716 39172 142772 39174
rect 142820 39226 142876 39228
rect 142820 39174 142822 39226
rect 142822 39174 142874 39226
rect 142874 39174 142876 39226
rect 142820 39172 142876 39174
rect 142924 39226 142980 39228
rect 142924 39174 142926 39226
rect 142926 39174 142978 39226
rect 142978 39174 142980 39226
rect 142924 39172 142980 39174
rect 142716 37658 142772 37660
rect 142716 37606 142718 37658
rect 142718 37606 142770 37658
rect 142770 37606 142772 37658
rect 142716 37604 142772 37606
rect 142820 37658 142876 37660
rect 142820 37606 142822 37658
rect 142822 37606 142874 37658
rect 142874 37606 142876 37658
rect 142820 37604 142876 37606
rect 142924 37658 142980 37660
rect 142924 37606 142926 37658
rect 142926 37606 142978 37658
rect 142978 37606 142980 37658
rect 142924 37604 142980 37606
rect 142716 36090 142772 36092
rect 142716 36038 142718 36090
rect 142718 36038 142770 36090
rect 142770 36038 142772 36090
rect 142716 36036 142772 36038
rect 142820 36090 142876 36092
rect 142820 36038 142822 36090
rect 142822 36038 142874 36090
rect 142874 36038 142876 36090
rect 142820 36036 142876 36038
rect 142924 36090 142980 36092
rect 142924 36038 142926 36090
rect 142926 36038 142978 36090
rect 142978 36038 142980 36090
rect 142924 36036 142980 36038
rect 142716 34522 142772 34524
rect 142716 34470 142718 34522
rect 142718 34470 142770 34522
rect 142770 34470 142772 34522
rect 142716 34468 142772 34470
rect 142820 34522 142876 34524
rect 142820 34470 142822 34522
rect 142822 34470 142874 34522
rect 142874 34470 142876 34522
rect 142820 34468 142876 34470
rect 142924 34522 142980 34524
rect 142924 34470 142926 34522
rect 142926 34470 142978 34522
rect 142978 34470 142980 34522
rect 142924 34468 142980 34470
rect 142716 32954 142772 32956
rect 142716 32902 142718 32954
rect 142718 32902 142770 32954
rect 142770 32902 142772 32954
rect 142716 32900 142772 32902
rect 142820 32954 142876 32956
rect 142820 32902 142822 32954
rect 142822 32902 142874 32954
rect 142874 32902 142876 32954
rect 142820 32900 142876 32902
rect 142924 32954 142980 32956
rect 142924 32902 142926 32954
rect 142926 32902 142978 32954
rect 142978 32902 142980 32954
rect 142924 32900 142980 32902
rect 142716 31386 142772 31388
rect 142716 31334 142718 31386
rect 142718 31334 142770 31386
rect 142770 31334 142772 31386
rect 142716 31332 142772 31334
rect 142820 31386 142876 31388
rect 142820 31334 142822 31386
rect 142822 31334 142874 31386
rect 142874 31334 142876 31386
rect 142820 31332 142876 31334
rect 142924 31386 142980 31388
rect 142924 31334 142926 31386
rect 142926 31334 142978 31386
rect 142978 31334 142980 31386
rect 142924 31332 142980 31334
rect 158076 54122 158132 54124
rect 158076 54070 158078 54122
rect 158078 54070 158130 54122
rect 158130 54070 158132 54122
rect 158076 54068 158132 54070
rect 158180 54122 158236 54124
rect 158180 54070 158182 54122
rect 158182 54070 158234 54122
rect 158234 54070 158236 54122
rect 158180 54068 158236 54070
rect 158284 54122 158340 54124
rect 158284 54070 158286 54122
rect 158286 54070 158338 54122
rect 158338 54070 158340 54122
rect 158284 54068 158340 54070
rect 158076 52554 158132 52556
rect 158076 52502 158078 52554
rect 158078 52502 158130 52554
rect 158130 52502 158132 52554
rect 158076 52500 158132 52502
rect 158180 52554 158236 52556
rect 158180 52502 158182 52554
rect 158182 52502 158234 52554
rect 158234 52502 158236 52554
rect 158180 52500 158236 52502
rect 158284 52554 158340 52556
rect 158284 52502 158286 52554
rect 158286 52502 158338 52554
rect 158338 52502 158340 52554
rect 158284 52500 158340 52502
rect 158076 50986 158132 50988
rect 158076 50934 158078 50986
rect 158078 50934 158130 50986
rect 158130 50934 158132 50986
rect 158076 50932 158132 50934
rect 158180 50986 158236 50988
rect 158180 50934 158182 50986
rect 158182 50934 158234 50986
rect 158234 50934 158236 50986
rect 158180 50932 158236 50934
rect 158284 50986 158340 50988
rect 158284 50934 158286 50986
rect 158286 50934 158338 50986
rect 158338 50934 158340 50986
rect 158284 50932 158340 50934
rect 158076 49418 158132 49420
rect 158076 49366 158078 49418
rect 158078 49366 158130 49418
rect 158130 49366 158132 49418
rect 158076 49364 158132 49366
rect 158180 49418 158236 49420
rect 158180 49366 158182 49418
rect 158182 49366 158234 49418
rect 158234 49366 158236 49418
rect 158180 49364 158236 49366
rect 158284 49418 158340 49420
rect 158284 49366 158286 49418
rect 158286 49366 158338 49418
rect 158338 49366 158340 49418
rect 158284 49364 158340 49366
rect 158076 47850 158132 47852
rect 158076 47798 158078 47850
rect 158078 47798 158130 47850
rect 158130 47798 158132 47850
rect 158076 47796 158132 47798
rect 158180 47850 158236 47852
rect 158180 47798 158182 47850
rect 158182 47798 158234 47850
rect 158234 47798 158236 47850
rect 158180 47796 158236 47798
rect 158284 47850 158340 47852
rect 158284 47798 158286 47850
rect 158286 47798 158338 47850
rect 158338 47798 158340 47850
rect 158284 47796 158340 47798
rect 158076 46282 158132 46284
rect 158076 46230 158078 46282
rect 158078 46230 158130 46282
rect 158130 46230 158132 46282
rect 158076 46228 158132 46230
rect 158180 46282 158236 46284
rect 158180 46230 158182 46282
rect 158182 46230 158234 46282
rect 158234 46230 158236 46282
rect 158180 46228 158236 46230
rect 158284 46282 158340 46284
rect 158284 46230 158286 46282
rect 158286 46230 158338 46282
rect 158338 46230 158340 46282
rect 158284 46228 158340 46230
rect 158076 44714 158132 44716
rect 158076 44662 158078 44714
rect 158078 44662 158130 44714
rect 158130 44662 158132 44714
rect 158076 44660 158132 44662
rect 158180 44714 158236 44716
rect 158180 44662 158182 44714
rect 158182 44662 158234 44714
rect 158234 44662 158236 44714
rect 158180 44660 158236 44662
rect 158284 44714 158340 44716
rect 158284 44662 158286 44714
rect 158286 44662 158338 44714
rect 158338 44662 158340 44714
rect 158284 44660 158340 44662
rect 158076 43146 158132 43148
rect 158076 43094 158078 43146
rect 158078 43094 158130 43146
rect 158130 43094 158132 43146
rect 158076 43092 158132 43094
rect 158180 43146 158236 43148
rect 158180 43094 158182 43146
rect 158182 43094 158234 43146
rect 158234 43094 158236 43146
rect 158180 43092 158236 43094
rect 158284 43146 158340 43148
rect 158284 43094 158286 43146
rect 158286 43094 158338 43146
rect 158338 43094 158340 43146
rect 158284 43092 158340 43094
rect 158076 41578 158132 41580
rect 158076 41526 158078 41578
rect 158078 41526 158130 41578
rect 158130 41526 158132 41578
rect 158076 41524 158132 41526
rect 158180 41578 158236 41580
rect 158180 41526 158182 41578
rect 158182 41526 158234 41578
rect 158234 41526 158236 41578
rect 158180 41524 158236 41526
rect 158284 41578 158340 41580
rect 158284 41526 158286 41578
rect 158286 41526 158338 41578
rect 158338 41526 158340 41578
rect 158284 41524 158340 41526
rect 158076 40010 158132 40012
rect 158076 39958 158078 40010
rect 158078 39958 158130 40010
rect 158130 39958 158132 40010
rect 158076 39956 158132 39958
rect 158180 40010 158236 40012
rect 158180 39958 158182 40010
rect 158182 39958 158234 40010
rect 158234 39958 158236 40010
rect 158180 39956 158236 39958
rect 158284 40010 158340 40012
rect 158284 39958 158286 40010
rect 158286 39958 158338 40010
rect 158338 39958 158340 40010
rect 158284 39956 158340 39958
rect 158076 38442 158132 38444
rect 158076 38390 158078 38442
rect 158078 38390 158130 38442
rect 158130 38390 158132 38442
rect 158076 38388 158132 38390
rect 158180 38442 158236 38444
rect 158180 38390 158182 38442
rect 158182 38390 158234 38442
rect 158234 38390 158236 38442
rect 158180 38388 158236 38390
rect 158284 38442 158340 38444
rect 158284 38390 158286 38442
rect 158286 38390 158338 38442
rect 158338 38390 158340 38442
rect 158284 38388 158340 38390
rect 158076 36874 158132 36876
rect 158076 36822 158078 36874
rect 158078 36822 158130 36874
rect 158130 36822 158132 36874
rect 158076 36820 158132 36822
rect 158180 36874 158236 36876
rect 158180 36822 158182 36874
rect 158182 36822 158234 36874
rect 158234 36822 158236 36874
rect 158180 36820 158236 36822
rect 158284 36874 158340 36876
rect 158284 36822 158286 36874
rect 158286 36822 158338 36874
rect 158338 36822 158340 36874
rect 158284 36820 158340 36822
rect 167916 54738 167972 54740
rect 167916 54686 167918 54738
rect 167918 54686 167970 54738
rect 167970 54686 167972 54738
rect 167916 54684 167972 54686
rect 184044 56140 184100 56196
rect 183372 55804 183428 55860
rect 182364 55410 182420 55412
rect 182364 55358 182366 55410
rect 182366 55358 182418 55410
rect 182418 55358 182420 55410
rect 182364 55356 182420 55358
rect 174972 55298 175028 55300
rect 174972 55246 174974 55298
rect 174974 55246 175026 55298
rect 175026 55246 175028 55298
rect 174972 55244 175028 55246
rect 175532 55298 175588 55300
rect 175532 55246 175534 55298
rect 175534 55246 175586 55298
rect 175586 55246 175588 55298
rect 175532 55244 175588 55246
rect 179452 55298 179508 55300
rect 179452 55246 179454 55298
rect 179454 55246 179506 55298
rect 179506 55246 179508 55298
rect 179452 55244 179508 55246
rect 173436 54906 173492 54908
rect 173436 54854 173438 54906
rect 173438 54854 173490 54906
rect 173490 54854 173492 54906
rect 173436 54852 173492 54854
rect 173540 54906 173596 54908
rect 173540 54854 173542 54906
rect 173542 54854 173594 54906
rect 173594 54854 173596 54906
rect 173540 54852 173596 54854
rect 173644 54906 173700 54908
rect 173644 54854 173646 54906
rect 173646 54854 173698 54906
rect 173698 54854 173700 54906
rect 173644 54852 173700 54854
rect 168924 54684 168980 54740
rect 172732 54738 172788 54740
rect 172732 54686 172734 54738
rect 172734 54686 172786 54738
rect 172786 54686 172788 54738
rect 172732 54684 172788 54686
rect 174300 54684 174356 54740
rect 166236 53564 166292 53620
rect 161980 51996 162036 52052
rect 161532 36204 161588 36260
rect 158076 35306 158132 35308
rect 158076 35254 158078 35306
rect 158078 35254 158130 35306
rect 158130 35254 158132 35306
rect 158076 35252 158132 35254
rect 158180 35306 158236 35308
rect 158180 35254 158182 35306
rect 158182 35254 158234 35306
rect 158234 35254 158236 35306
rect 158180 35252 158236 35254
rect 158284 35306 158340 35308
rect 158284 35254 158286 35306
rect 158286 35254 158338 35306
rect 158338 35254 158340 35306
rect 158284 35252 158340 35254
rect 167468 53618 167524 53620
rect 167468 53566 167470 53618
rect 167470 53566 167522 53618
rect 167522 53566 167524 53618
rect 167468 53564 167524 53566
rect 167132 34636 167188 34692
rect 158076 33738 158132 33740
rect 158076 33686 158078 33738
rect 158078 33686 158130 33738
rect 158130 33686 158132 33738
rect 158076 33684 158132 33686
rect 158180 33738 158236 33740
rect 158180 33686 158182 33738
rect 158182 33686 158234 33738
rect 158234 33686 158236 33738
rect 158180 33684 158236 33686
rect 158284 33738 158340 33740
rect 158284 33686 158286 33738
rect 158286 33686 158338 33738
rect 158338 33686 158340 33738
rect 158284 33684 158340 33686
rect 156380 32732 156436 32788
rect 158076 32170 158132 32172
rect 158076 32118 158078 32170
rect 158078 32118 158130 32170
rect 158130 32118 158132 32170
rect 158076 32116 158132 32118
rect 158180 32170 158236 32172
rect 158180 32118 158182 32170
rect 158182 32118 158234 32170
rect 158234 32118 158236 32170
rect 158180 32116 158236 32118
rect 158284 32170 158340 32172
rect 158284 32118 158286 32170
rect 158286 32118 158338 32170
rect 158338 32118 158340 32170
rect 158284 32116 158340 32118
rect 150780 31052 150836 31108
rect 158076 30602 158132 30604
rect 158076 30550 158078 30602
rect 158078 30550 158130 30602
rect 158130 30550 158132 30602
rect 158076 30548 158132 30550
rect 158180 30602 158236 30604
rect 158180 30550 158182 30602
rect 158182 30550 158234 30602
rect 158234 30550 158236 30602
rect 158180 30548 158236 30550
rect 158284 30602 158340 30604
rect 158284 30550 158286 30602
rect 158286 30550 158338 30602
rect 158338 30550 158340 30602
rect 158284 30548 158340 30550
rect 142716 29818 142772 29820
rect 142716 29766 142718 29818
rect 142718 29766 142770 29818
rect 142770 29766 142772 29818
rect 142716 29764 142772 29766
rect 142820 29818 142876 29820
rect 142820 29766 142822 29818
rect 142822 29766 142874 29818
rect 142874 29766 142876 29818
rect 142820 29764 142876 29766
rect 142924 29818 142980 29820
rect 142924 29766 142926 29818
rect 142926 29766 142978 29818
rect 142978 29766 142980 29818
rect 142924 29764 142980 29766
rect 140252 29372 140308 29428
rect 158076 29034 158132 29036
rect 158076 28982 158078 29034
rect 158078 28982 158130 29034
rect 158130 28982 158132 29034
rect 158076 28980 158132 28982
rect 158180 29034 158236 29036
rect 158180 28982 158182 29034
rect 158182 28982 158234 29034
rect 158234 28982 158236 29034
rect 158180 28980 158236 28982
rect 158284 29034 158340 29036
rect 158284 28982 158286 29034
rect 158286 28982 158338 29034
rect 158338 28982 158340 29034
rect 158284 28980 158340 28982
rect 142716 28250 142772 28252
rect 142716 28198 142718 28250
rect 142718 28198 142770 28250
rect 142770 28198 142772 28250
rect 142716 28196 142772 28198
rect 142820 28250 142876 28252
rect 142820 28198 142822 28250
rect 142822 28198 142874 28250
rect 142874 28198 142876 28250
rect 142820 28196 142876 28198
rect 142924 28250 142980 28252
rect 142924 28198 142926 28250
rect 142926 28198 142978 28250
rect 142978 28198 142980 28250
rect 142924 28196 142980 28198
rect 158076 27466 158132 27468
rect 158076 27414 158078 27466
rect 158078 27414 158130 27466
rect 158130 27414 158132 27466
rect 158076 27412 158132 27414
rect 158180 27466 158236 27468
rect 158180 27414 158182 27466
rect 158182 27414 158234 27466
rect 158234 27414 158236 27466
rect 158180 27412 158236 27414
rect 158284 27466 158340 27468
rect 158284 27414 158286 27466
rect 158286 27414 158338 27466
rect 158338 27414 158340 27466
rect 158284 27412 158340 27414
rect 142716 26682 142772 26684
rect 142716 26630 142718 26682
rect 142718 26630 142770 26682
rect 142770 26630 142772 26682
rect 142716 26628 142772 26630
rect 142820 26682 142876 26684
rect 142820 26630 142822 26682
rect 142822 26630 142874 26682
rect 142874 26630 142876 26682
rect 142820 26628 142876 26630
rect 142924 26682 142980 26684
rect 142924 26630 142926 26682
rect 142926 26630 142978 26682
rect 142978 26630 142980 26682
rect 142924 26628 142980 26630
rect 134876 26012 134932 26068
rect 158076 25898 158132 25900
rect 158076 25846 158078 25898
rect 158078 25846 158130 25898
rect 158130 25846 158132 25898
rect 158076 25844 158132 25846
rect 158180 25898 158236 25900
rect 158180 25846 158182 25898
rect 158182 25846 158234 25898
rect 158234 25846 158236 25898
rect 158180 25844 158236 25846
rect 158284 25898 158340 25900
rect 158284 25846 158286 25898
rect 158286 25846 158338 25898
rect 158338 25846 158340 25898
rect 158284 25844 158340 25846
rect 142716 25114 142772 25116
rect 142716 25062 142718 25114
rect 142718 25062 142770 25114
rect 142770 25062 142772 25114
rect 142716 25060 142772 25062
rect 142820 25114 142876 25116
rect 142820 25062 142822 25114
rect 142822 25062 142874 25114
rect 142874 25062 142876 25114
rect 142820 25060 142876 25062
rect 142924 25114 142980 25116
rect 142924 25062 142926 25114
rect 142926 25062 142978 25114
rect 142978 25062 142980 25114
rect 142924 25060 142980 25062
rect 129388 24444 129444 24500
rect 127356 24330 127412 24332
rect 127356 24278 127358 24330
rect 127358 24278 127410 24330
rect 127410 24278 127412 24330
rect 127356 24276 127412 24278
rect 127460 24330 127516 24332
rect 127460 24278 127462 24330
rect 127462 24278 127514 24330
rect 127514 24278 127516 24330
rect 127460 24276 127516 24278
rect 127564 24330 127620 24332
rect 127564 24278 127566 24330
rect 127566 24278 127618 24330
rect 127618 24278 127620 24330
rect 127564 24276 127620 24278
rect 158076 24330 158132 24332
rect 158076 24278 158078 24330
rect 158078 24278 158130 24330
rect 158130 24278 158132 24330
rect 158076 24276 158132 24278
rect 158180 24330 158236 24332
rect 158180 24278 158182 24330
rect 158182 24278 158234 24330
rect 158234 24278 158236 24330
rect 158180 24276 158236 24278
rect 158284 24330 158340 24332
rect 158284 24278 158286 24330
rect 158286 24278 158338 24330
rect 158338 24278 158340 24330
rect 158284 24276 158340 24278
rect 111996 23546 112052 23548
rect 111996 23494 111998 23546
rect 111998 23494 112050 23546
rect 112050 23494 112052 23546
rect 111996 23492 112052 23494
rect 112100 23546 112156 23548
rect 112100 23494 112102 23546
rect 112102 23494 112154 23546
rect 112154 23494 112156 23546
rect 112100 23492 112156 23494
rect 112204 23546 112260 23548
rect 112204 23494 112206 23546
rect 112206 23494 112258 23546
rect 112258 23494 112260 23546
rect 112204 23492 112260 23494
rect 142716 23546 142772 23548
rect 142716 23494 142718 23546
rect 142718 23494 142770 23546
rect 142770 23494 142772 23546
rect 142716 23492 142772 23494
rect 142820 23546 142876 23548
rect 142820 23494 142822 23546
rect 142822 23494 142874 23546
rect 142874 23494 142876 23546
rect 142820 23492 142876 23494
rect 142924 23546 142980 23548
rect 142924 23494 142926 23546
rect 142926 23494 142978 23546
rect 142978 23494 142980 23546
rect 142924 23492 142980 23494
rect 127356 22762 127412 22764
rect 127356 22710 127358 22762
rect 127358 22710 127410 22762
rect 127410 22710 127412 22762
rect 127356 22708 127412 22710
rect 127460 22762 127516 22764
rect 127460 22710 127462 22762
rect 127462 22710 127514 22762
rect 127514 22710 127516 22762
rect 127460 22708 127516 22710
rect 127564 22762 127620 22764
rect 127564 22710 127566 22762
rect 127566 22710 127618 22762
rect 127618 22710 127620 22762
rect 127564 22708 127620 22710
rect 158076 22762 158132 22764
rect 158076 22710 158078 22762
rect 158078 22710 158130 22762
rect 158130 22710 158132 22762
rect 158076 22708 158132 22710
rect 158180 22762 158236 22764
rect 158180 22710 158182 22762
rect 158182 22710 158234 22762
rect 158234 22710 158236 22762
rect 158180 22708 158236 22710
rect 158284 22762 158340 22764
rect 158284 22710 158286 22762
rect 158286 22710 158338 22762
rect 158338 22710 158340 22762
rect 158284 22708 158340 22710
rect 111996 21978 112052 21980
rect 111996 21926 111998 21978
rect 111998 21926 112050 21978
rect 112050 21926 112052 21978
rect 111996 21924 112052 21926
rect 112100 21978 112156 21980
rect 112100 21926 112102 21978
rect 112102 21926 112154 21978
rect 112154 21926 112156 21978
rect 112100 21924 112156 21926
rect 112204 21978 112260 21980
rect 112204 21926 112206 21978
rect 112206 21926 112258 21978
rect 112258 21926 112260 21978
rect 112204 21924 112260 21926
rect 142716 21978 142772 21980
rect 142716 21926 142718 21978
rect 142718 21926 142770 21978
rect 142770 21926 142772 21978
rect 142716 21924 142772 21926
rect 142820 21978 142876 21980
rect 142820 21926 142822 21978
rect 142822 21926 142874 21978
rect 142874 21926 142876 21978
rect 142820 21924 142876 21926
rect 142924 21978 142980 21980
rect 142924 21926 142926 21978
rect 142926 21926 142978 21978
rect 142978 21926 142980 21978
rect 142924 21924 142980 21926
rect 127356 21194 127412 21196
rect 127356 21142 127358 21194
rect 127358 21142 127410 21194
rect 127410 21142 127412 21194
rect 127356 21140 127412 21142
rect 127460 21194 127516 21196
rect 127460 21142 127462 21194
rect 127462 21142 127514 21194
rect 127514 21142 127516 21194
rect 127460 21140 127516 21142
rect 127564 21194 127620 21196
rect 127564 21142 127566 21194
rect 127566 21142 127618 21194
rect 127618 21142 127620 21194
rect 127564 21140 127620 21142
rect 158076 21194 158132 21196
rect 158076 21142 158078 21194
rect 158078 21142 158130 21194
rect 158130 21142 158132 21194
rect 158076 21140 158132 21142
rect 158180 21194 158236 21196
rect 158180 21142 158182 21194
rect 158182 21142 158234 21194
rect 158234 21142 158236 21194
rect 158180 21140 158236 21142
rect 158284 21194 158340 21196
rect 158284 21142 158286 21194
rect 158286 21142 158338 21194
rect 158338 21142 158340 21194
rect 158284 21140 158340 21142
rect 111996 20410 112052 20412
rect 111996 20358 111998 20410
rect 111998 20358 112050 20410
rect 112050 20358 112052 20410
rect 111996 20356 112052 20358
rect 112100 20410 112156 20412
rect 112100 20358 112102 20410
rect 112102 20358 112154 20410
rect 112154 20358 112156 20410
rect 112100 20356 112156 20358
rect 112204 20410 112260 20412
rect 112204 20358 112206 20410
rect 112206 20358 112258 20410
rect 112258 20358 112260 20410
rect 112204 20356 112260 20358
rect 142716 20410 142772 20412
rect 142716 20358 142718 20410
rect 142718 20358 142770 20410
rect 142770 20358 142772 20410
rect 142716 20356 142772 20358
rect 142820 20410 142876 20412
rect 142820 20358 142822 20410
rect 142822 20358 142874 20410
rect 142874 20358 142876 20410
rect 142820 20356 142876 20358
rect 142924 20410 142980 20412
rect 142924 20358 142926 20410
rect 142926 20358 142978 20410
rect 142978 20358 142980 20410
rect 142924 20356 142980 20358
rect 127356 19626 127412 19628
rect 127356 19574 127358 19626
rect 127358 19574 127410 19626
rect 127410 19574 127412 19626
rect 127356 19572 127412 19574
rect 127460 19626 127516 19628
rect 127460 19574 127462 19626
rect 127462 19574 127514 19626
rect 127514 19574 127516 19626
rect 127460 19572 127516 19574
rect 127564 19626 127620 19628
rect 127564 19574 127566 19626
rect 127566 19574 127618 19626
rect 127618 19574 127620 19626
rect 127564 19572 127620 19574
rect 158076 19626 158132 19628
rect 158076 19574 158078 19626
rect 158078 19574 158130 19626
rect 158130 19574 158132 19626
rect 158076 19572 158132 19574
rect 158180 19626 158236 19628
rect 158180 19574 158182 19626
rect 158182 19574 158234 19626
rect 158234 19574 158236 19626
rect 158180 19572 158236 19574
rect 158284 19626 158340 19628
rect 158284 19574 158286 19626
rect 158286 19574 158338 19626
rect 158338 19574 158340 19626
rect 158284 19572 158340 19574
rect 111996 18842 112052 18844
rect 111996 18790 111998 18842
rect 111998 18790 112050 18842
rect 112050 18790 112052 18842
rect 111996 18788 112052 18790
rect 112100 18842 112156 18844
rect 112100 18790 112102 18842
rect 112102 18790 112154 18842
rect 112154 18790 112156 18842
rect 112100 18788 112156 18790
rect 112204 18842 112260 18844
rect 112204 18790 112206 18842
rect 112206 18790 112258 18842
rect 112258 18790 112260 18842
rect 112204 18788 112260 18790
rect 142716 18842 142772 18844
rect 142716 18790 142718 18842
rect 142718 18790 142770 18842
rect 142770 18790 142772 18842
rect 142716 18788 142772 18790
rect 142820 18842 142876 18844
rect 142820 18790 142822 18842
rect 142822 18790 142874 18842
rect 142874 18790 142876 18842
rect 142820 18788 142876 18790
rect 142924 18842 142980 18844
rect 142924 18790 142926 18842
rect 142926 18790 142978 18842
rect 142978 18790 142980 18842
rect 142924 18788 142980 18790
rect 127356 18058 127412 18060
rect 127356 18006 127358 18058
rect 127358 18006 127410 18058
rect 127410 18006 127412 18058
rect 127356 18004 127412 18006
rect 127460 18058 127516 18060
rect 127460 18006 127462 18058
rect 127462 18006 127514 18058
rect 127514 18006 127516 18058
rect 127460 18004 127516 18006
rect 127564 18058 127620 18060
rect 127564 18006 127566 18058
rect 127566 18006 127618 18058
rect 127618 18006 127620 18058
rect 127564 18004 127620 18006
rect 158076 18058 158132 18060
rect 158076 18006 158078 18058
rect 158078 18006 158130 18058
rect 158130 18006 158132 18058
rect 158076 18004 158132 18006
rect 158180 18058 158236 18060
rect 158180 18006 158182 18058
rect 158182 18006 158234 18058
rect 158234 18006 158236 18058
rect 158180 18004 158236 18006
rect 158284 18058 158340 18060
rect 158284 18006 158286 18058
rect 158286 18006 158338 18058
rect 158338 18006 158340 18058
rect 158284 18004 158340 18006
rect 111996 17274 112052 17276
rect 111996 17222 111998 17274
rect 111998 17222 112050 17274
rect 112050 17222 112052 17274
rect 111996 17220 112052 17222
rect 112100 17274 112156 17276
rect 112100 17222 112102 17274
rect 112102 17222 112154 17274
rect 112154 17222 112156 17274
rect 112100 17220 112156 17222
rect 112204 17274 112260 17276
rect 112204 17222 112206 17274
rect 112206 17222 112258 17274
rect 112258 17222 112260 17274
rect 112204 17220 112260 17222
rect 142716 17274 142772 17276
rect 142716 17222 142718 17274
rect 142718 17222 142770 17274
rect 142770 17222 142772 17274
rect 142716 17220 142772 17222
rect 142820 17274 142876 17276
rect 142820 17222 142822 17274
rect 142822 17222 142874 17274
rect 142874 17222 142876 17274
rect 142820 17220 142876 17222
rect 142924 17274 142980 17276
rect 142924 17222 142926 17274
rect 142926 17222 142978 17274
rect 142978 17222 142980 17274
rect 142924 17220 142980 17222
rect 127356 16490 127412 16492
rect 127356 16438 127358 16490
rect 127358 16438 127410 16490
rect 127410 16438 127412 16490
rect 127356 16436 127412 16438
rect 127460 16490 127516 16492
rect 127460 16438 127462 16490
rect 127462 16438 127514 16490
rect 127514 16438 127516 16490
rect 127460 16436 127516 16438
rect 127564 16490 127620 16492
rect 127564 16438 127566 16490
rect 127566 16438 127618 16490
rect 127618 16438 127620 16490
rect 127564 16436 127620 16438
rect 158076 16490 158132 16492
rect 158076 16438 158078 16490
rect 158078 16438 158130 16490
rect 158130 16438 158132 16490
rect 158076 16436 158132 16438
rect 158180 16490 158236 16492
rect 158180 16438 158182 16490
rect 158182 16438 158234 16490
rect 158234 16438 158236 16490
rect 158180 16436 158236 16438
rect 158284 16490 158340 16492
rect 158284 16438 158286 16490
rect 158286 16438 158338 16490
rect 158338 16438 158340 16490
rect 158284 16436 158340 16438
rect 107660 15932 107716 15988
rect 111996 15706 112052 15708
rect 111996 15654 111998 15706
rect 111998 15654 112050 15706
rect 112050 15654 112052 15706
rect 111996 15652 112052 15654
rect 112100 15706 112156 15708
rect 112100 15654 112102 15706
rect 112102 15654 112154 15706
rect 112154 15654 112156 15706
rect 112100 15652 112156 15654
rect 112204 15706 112260 15708
rect 112204 15654 112206 15706
rect 112206 15654 112258 15706
rect 112258 15654 112260 15706
rect 112204 15652 112260 15654
rect 142716 15706 142772 15708
rect 142716 15654 142718 15706
rect 142718 15654 142770 15706
rect 142770 15654 142772 15706
rect 142716 15652 142772 15654
rect 142820 15706 142876 15708
rect 142820 15654 142822 15706
rect 142822 15654 142874 15706
rect 142874 15654 142876 15706
rect 142820 15652 142876 15654
rect 142924 15706 142980 15708
rect 142924 15654 142926 15706
rect 142926 15654 142978 15706
rect 142978 15654 142980 15706
rect 142924 15652 142980 15654
rect 127356 14922 127412 14924
rect 127356 14870 127358 14922
rect 127358 14870 127410 14922
rect 127410 14870 127412 14922
rect 127356 14868 127412 14870
rect 127460 14922 127516 14924
rect 127460 14870 127462 14922
rect 127462 14870 127514 14922
rect 127514 14870 127516 14922
rect 127460 14868 127516 14870
rect 127564 14922 127620 14924
rect 127564 14870 127566 14922
rect 127566 14870 127618 14922
rect 127618 14870 127620 14922
rect 127564 14868 127620 14870
rect 158076 14922 158132 14924
rect 158076 14870 158078 14922
rect 158078 14870 158130 14922
rect 158130 14870 158132 14922
rect 158076 14868 158132 14870
rect 158180 14922 158236 14924
rect 158180 14870 158182 14922
rect 158182 14870 158234 14922
rect 158234 14870 158236 14922
rect 158180 14868 158236 14870
rect 158284 14922 158340 14924
rect 158284 14870 158286 14922
rect 158286 14870 158338 14922
rect 158338 14870 158340 14922
rect 158284 14868 158340 14870
rect 111996 14138 112052 14140
rect 111996 14086 111998 14138
rect 111998 14086 112050 14138
rect 112050 14086 112052 14138
rect 111996 14084 112052 14086
rect 112100 14138 112156 14140
rect 112100 14086 112102 14138
rect 112102 14086 112154 14138
rect 112154 14086 112156 14138
rect 112100 14084 112156 14086
rect 112204 14138 112260 14140
rect 112204 14086 112206 14138
rect 112206 14086 112258 14138
rect 112258 14086 112260 14138
rect 112204 14084 112260 14086
rect 142716 14138 142772 14140
rect 142716 14086 142718 14138
rect 142718 14086 142770 14138
rect 142770 14086 142772 14138
rect 142716 14084 142772 14086
rect 142820 14138 142876 14140
rect 142820 14086 142822 14138
rect 142822 14086 142874 14138
rect 142874 14086 142876 14138
rect 142820 14084 142876 14086
rect 142924 14138 142980 14140
rect 142924 14086 142926 14138
rect 142926 14086 142978 14138
rect 142978 14086 142980 14138
rect 142924 14084 142980 14086
rect 127356 13354 127412 13356
rect 127356 13302 127358 13354
rect 127358 13302 127410 13354
rect 127410 13302 127412 13354
rect 127356 13300 127412 13302
rect 127460 13354 127516 13356
rect 127460 13302 127462 13354
rect 127462 13302 127514 13354
rect 127514 13302 127516 13354
rect 127460 13300 127516 13302
rect 127564 13354 127620 13356
rect 127564 13302 127566 13354
rect 127566 13302 127618 13354
rect 127618 13302 127620 13354
rect 127564 13300 127620 13302
rect 158076 13354 158132 13356
rect 158076 13302 158078 13354
rect 158078 13302 158130 13354
rect 158130 13302 158132 13354
rect 158076 13300 158132 13302
rect 158180 13354 158236 13356
rect 158180 13302 158182 13354
rect 158182 13302 158234 13354
rect 158234 13302 158236 13354
rect 158180 13300 158236 13302
rect 158284 13354 158340 13356
rect 158284 13302 158286 13354
rect 158286 13302 158338 13354
rect 158338 13302 158340 13354
rect 158284 13300 158340 13302
rect 111996 12570 112052 12572
rect 111996 12518 111998 12570
rect 111998 12518 112050 12570
rect 112050 12518 112052 12570
rect 111996 12516 112052 12518
rect 112100 12570 112156 12572
rect 112100 12518 112102 12570
rect 112102 12518 112154 12570
rect 112154 12518 112156 12570
rect 112100 12516 112156 12518
rect 112204 12570 112260 12572
rect 112204 12518 112206 12570
rect 112206 12518 112258 12570
rect 112258 12518 112260 12570
rect 112204 12516 112260 12518
rect 142716 12570 142772 12572
rect 142716 12518 142718 12570
rect 142718 12518 142770 12570
rect 142770 12518 142772 12570
rect 142716 12516 142772 12518
rect 142820 12570 142876 12572
rect 142820 12518 142822 12570
rect 142822 12518 142874 12570
rect 142874 12518 142876 12570
rect 142820 12516 142876 12518
rect 142924 12570 142980 12572
rect 142924 12518 142926 12570
rect 142926 12518 142978 12570
rect 142978 12518 142980 12570
rect 142924 12516 142980 12518
rect 127356 11786 127412 11788
rect 127356 11734 127358 11786
rect 127358 11734 127410 11786
rect 127410 11734 127412 11786
rect 127356 11732 127412 11734
rect 127460 11786 127516 11788
rect 127460 11734 127462 11786
rect 127462 11734 127514 11786
rect 127514 11734 127516 11786
rect 127460 11732 127516 11734
rect 127564 11786 127620 11788
rect 127564 11734 127566 11786
rect 127566 11734 127618 11786
rect 127618 11734 127620 11786
rect 127564 11732 127620 11734
rect 158076 11786 158132 11788
rect 158076 11734 158078 11786
rect 158078 11734 158130 11786
rect 158130 11734 158132 11786
rect 158076 11732 158132 11734
rect 158180 11786 158236 11788
rect 158180 11734 158182 11786
rect 158182 11734 158234 11786
rect 158234 11734 158236 11786
rect 158180 11732 158236 11734
rect 158284 11786 158340 11788
rect 158284 11734 158286 11786
rect 158286 11734 158338 11786
rect 158338 11734 158340 11786
rect 158284 11732 158340 11734
rect 179452 53788 179508 53844
rect 180124 53842 180180 53844
rect 180124 53790 180126 53842
rect 180126 53790 180178 53842
rect 180178 53790 180180 53842
rect 180124 53788 180180 53790
rect 182140 53788 182196 53844
rect 177660 53618 177716 53620
rect 177660 53566 177662 53618
rect 177662 53566 177714 53618
rect 177714 53566 177716 53618
rect 177660 53564 177716 53566
rect 178108 53564 178164 53620
rect 173436 53338 173492 53340
rect 173436 53286 173438 53338
rect 173438 53286 173490 53338
rect 173490 53286 173492 53338
rect 173436 53284 173492 53286
rect 173540 53338 173596 53340
rect 173540 53286 173542 53338
rect 173542 53286 173594 53338
rect 173594 53286 173596 53338
rect 173540 53284 173596 53286
rect 173644 53338 173700 53340
rect 173644 53286 173646 53338
rect 173646 53286 173698 53338
rect 173698 53286 173700 53338
rect 173644 53284 173700 53286
rect 182812 53788 182868 53844
rect 185052 56194 185108 56196
rect 185052 56142 185054 56194
rect 185054 56142 185106 56194
rect 185106 56142 185108 56194
rect 185052 56140 185108 56142
rect 187180 56140 187236 56196
rect 186172 55410 186228 55412
rect 186172 55358 186174 55410
rect 186174 55358 186226 55410
rect 186226 55358 186228 55410
rect 186172 55356 186228 55358
rect 186396 55410 186452 55412
rect 186396 55358 186398 55410
rect 186398 55358 186450 55410
rect 186450 55358 186452 55410
rect 186396 55356 186452 55358
rect 189868 56194 189924 56196
rect 189868 56142 189870 56194
rect 189870 56142 189922 56194
rect 189922 56142 189924 56194
rect 189868 56140 189924 56142
rect 190876 56082 190932 56084
rect 190876 56030 190878 56082
rect 190878 56030 190930 56082
rect 190930 56030 190932 56082
rect 190876 56028 190932 56030
rect 187852 55970 187908 55972
rect 187852 55918 187854 55970
rect 187854 55918 187906 55970
rect 187906 55918 187908 55970
rect 187852 55916 187908 55918
rect 189084 55970 189140 55972
rect 189084 55918 189086 55970
rect 189086 55918 189138 55970
rect 189138 55918 189140 55970
rect 189084 55916 189140 55918
rect 188796 55690 188852 55692
rect 188796 55638 188798 55690
rect 188798 55638 188850 55690
rect 188850 55638 188852 55690
rect 188796 55636 188852 55638
rect 188900 55690 188956 55692
rect 188900 55638 188902 55690
rect 188902 55638 188954 55690
rect 188954 55638 188956 55690
rect 188900 55636 188956 55638
rect 189004 55690 189060 55692
rect 189004 55638 189006 55690
rect 189006 55638 189058 55690
rect 189058 55638 189060 55690
rect 189004 55636 189060 55638
rect 193900 56140 193956 56196
rect 191772 56028 191828 56084
rect 188300 55410 188356 55412
rect 188300 55358 188302 55410
rect 188302 55358 188354 55410
rect 188354 55358 188356 55410
rect 188300 55356 188356 55358
rect 186956 55186 187012 55188
rect 186956 55134 186958 55186
rect 186958 55134 187010 55186
rect 187010 55134 187012 55186
rect 186956 55132 187012 55134
rect 187516 55186 187572 55188
rect 187516 55134 187518 55186
rect 187518 55134 187570 55186
rect 187570 55134 187572 55186
rect 187516 55132 187572 55134
rect 183372 53452 183428 53508
rect 186508 53676 186564 53732
rect 182476 53116 182532 53172
rect 185836 53170 185892 53172
rect 185836 53118 185838 53170
rect 185838 53118 185890 53170
rect 185890 53118 185892 53170
rect 185836 53116 185892 53118
rect 187964 53676 188020 53732
rect 186508 53116 186564 53172
rect 181468 52834 181524 52836
rect 181468 52782 181470 52834
rect 181470 52782 181522 52834
rect 181522 52782 181524 52834
rect 181468 52780 181524 52782
rect 183260 52834 183316 52836
rect 183260 52782 183262 52834
rect 183262 52782 183314 52834
rect 183314 52782 183316 52834
rect 183260 52780 183316 52782
rect 173436 51770 173492 51772
rect 173436 51718 173438 51770
rect 173438 51718 173490 51770
rect 173490 51718 173492 51770
rect 173436 51716 173492 51718
rect 173540 51770 173596 51772
rect 173540 51718 173542 51770
rect 173542 51718 173594 51770
rect 173594 51718 173596 51770
rect 173540 51716 173596 51718
rect 173644 51770 173700 51772
rect 173644 51718 173646 51770
rect 173646 51718 173698 51770
rect 173698 51718 173700 51770
rect 173644 51716 173700 51718
rect 173436 50202 173492 50204
rect 173436 50150 173438 50202
rect 173438 50150 173490 50202
rect 173490 50150 173492 50202
rect 173436 50148 173492 50150
rect 173540 50202 173596 50204
rect 173540 50150 173542 50202
rect 173542 50150 173594 50202
rect 173594 50150 173596 50202
rect 173540 50148 173596 50150
rect 173644 50202 173700 50204
rect 173644 50150 173646 50202
rect 173646 50150 173698 50202
rect 173698 50150 173700 50202
rect 173644 50148 173700 50150
rect 173436 48634 173492 48636
rect 173436 48582 173438 48634
rect 173438 48582 173490 48634
rect 173490 48582 173492 48634
rect 173436 48580 173492 48582
rect 173540 48634 173596 48636
rect 173540 48582 173542 48634
rect 173542 48582 173594 48634
rect 173594 48582 173596 48634
rect 173540 48580 173596 48582
rect 173644 48634 173700 48636
rect 173644 48582 173646 48634
rect 173646 48582 173698 48634
rect 173698 48582 173700 48634
rect 173644 48580 173700 48582
rect 173436 47066 173492 47068
rect 173436 47014 173438 47066
rect 173438 47014 173490 47066
rect 173490 47014 173492 47066
rect 173436 47012 173492 47014
rect 173540 47066 173596 47068
rect 173540 47014 173542 47066
rect 173542 47014 173594 47066
rect 173594 47014 173596 47066
rect 173540 47012 173596 47014
rect 173644 47066 173700 47068
rect 173644 47014 173646 47066
rect 173646 47014 173698 47066
rect 173698 47014 173700 47066
rect 173644 47012 173700 47014
rect 173436 45498 173492 45500
rect 173436 45446 173438 45498
rect 173438 45446 173490 45498
rect 173490 45446 173492 45498
rect 173436 45444 173492 45446
rect 173540 45498 173596 45500
rect 173540 45446 173542 45498
rect 173542 45446 173594 45498
rect 173594 45446 173596 45498
rect 173540 45444 173596 45446
rect 173644 45498 173700 45500
rect 173644 45446 173646 45498
rect 173646 45446 173698 45498
rect 173698 45446 173700 45498
rect 173644 45444 173700 45446
rect 173436 43930 173492 43932
rect 173436 43878 173438 43930
rect 173438 43878 173490 43930
rect 173490 43878 173492 43930
rect 173436 43876 173492 43878
rect 173540 43930 173596 43932
rect 173540 43878 173542 43930
rect 173542 43878 173594 43930
rect 173594 43878 173596 43930
rect 173540 43876 173596 43878
rect 173644 43930 173700 43932
rect 173644 43878 173646 43930
rect 173646 43878 173698 43930
rect 173698 43878 173700 43930
rect 173644 43876 173700 43878
rect 173436 42362 173492 42364
rect 173436 42310 173438 42362
rect 173438 42310 173490 42362
rect 173490 42310 173492 42362
rect 173436 42308 173492 42310
rect 173540 42362 173596 42364
rect 173540 42310 173542 42362
rect 173542 42310 173594 42362
rect 173594 42310 173596 42362
rect 173540 42308 173596 42310
rect 173644 42362 173700 42364
rect 173644 42310 173646 42362
rect 173646 42310 173698 42362
rect 173698 42310 173700 42362
rect 173644 42308 173700 42310
rect 173436 40794 173492 40796
rect 173436 40742 173438 40794
rect 173438 40742 173490 40794
rect 173490 40742 173492 40794
rect 173436 40740 173492 40742
rect 173540 40794 173596 40796
rect 173540 40742 173542 40794
rect 173542 40742 173594 40794
rect 173594 40742 173596 40794
rect 173540 40740 173596 40742
rect 173644 40794 173700 40796
rect 173644 40742 173646 40794
rect 173646 40742 173698 40794
rect 173698 40742 173700 40794
rect 173644 40740 173700 40742
rect 173436 39226 173492 39228
rect 173436 39174 173438 39226
rect 173438 39174 173490 39226
rect 173490 39174 173492 39226
rect 173436 39172 173492 39174
rect 173540 39226 173596 39228
rect 173540 39174 173542 39226
rect 173542 39174 173594 39226
rect 173594 39174 173596 39226
rect 173540 39172 173596 39174
rect 173644 39226 173700 39228
rect 173644 39174 173646 39226
rect 173646 39174 173698 39226
rect 173698 39174 173700 39226
rect 173644 39172 173700 39174
rect 173436 37658 173492 37660
rect 173436 37606 173438 37658
rect 173438 37606 173490 37658
rect 173490 37606 173492 37658
rect 173436 37604 173492 37606
rect 173540 37658 173596 37660
rect 173540 37606 173542 37658
rect 173542 37606 173594 37658
rect 173594 37606 173596 37658
rect 173540 37604 173596 37606
rect 173644 37658 173700 37660
rect 173644 37606 173646 37658
rect 173646 37606 173698 37658
rect 173698 37606 173700 37658
rect 173644 37604 173700 37606
rect 173436 36090 173492 36092
rect 173436 36038 173438 36090
rect 173438 36038 173490 36090
rect 173490 36038 173492 36090
rect 173436 36036 173492 36038
rect 173540 36090 173596 36092
rect 173540 36038 173542 36090
rect 173542 36038 173594 36090
rect 173594 36038 173596 36090
rect 173540 36036 173596 36038
rect 173644 36090 173700 36092
rect 173644 36038 173646 36090
rect 173646 36038 173698 36090
rect 173698 36038 173700 36090
rect 173644 36036 173700 36038
rect 173436 34522 173492 34524
rect 173436 34470 173438 34522
rect 173438 34470 173490 34522
rect 173490 34470 173492 34522
rect 173436 34468 173492 34470
rect 173540 34522 173596 34524
rect 173540 34470 173542 34522
rect 173542 34470 173594 34522
rect 173594 34470 173596 34522
rect 173540 34468 173596 34470
rect 173644 34522 173700 34524
rect 173644 34470 173646 34522
rect 173646 34470 173698 34522
rect 173698 34470 173700 34522
rect 173644 34468 173700 34470
rect 173436 32954 173492 32956
rect 173436 32902 173438 32954
rect 173438 32902 173490 32954
rect 173490 32902 173492 32954
rect 173436 32900 173492 32902
rect 173540 32954 173596 32956
rect 173540 32902 173542 32954
rect 173542 32902 173594 32954
rect 173594 32902 173596 32954
rect 173540 32900 173596 32902
rect 173644 32954 173700 32956
rect 173644 32902 173646 32954
rect 173646 32902 173698 32954
rect 173698 32902 173700 32954
rect 173644 32900 173700 32902
rect 173436 31386 173492 31388
rect 173436 31334 173438 31386
rect 173438 31334 173490 31386
rect 173490 31334 173492 31386
rect 173436 31332 173492 31334
rect 173540 31386 173596 31388
rect 173540 31334 173542 31386
rect 173542 31334 173594 31386
rect 173594 31334 173596 31386
rect 173540 31332 173596 31334
rect 173644 31386 173700 31388
rect 173644 31334 173646 31386
rect 173646 31334 173698 31386
rect 173698 31334 173700 31386
rect 173644 31332 173700 31334
rect 173436 29818 173492 29820
rect 173436 29766 173438 29818
rect 173438 29766 173490 29818
rect 173490 29766 173492 29818
rect 173436 29764 173492 29766
rect 173540 29818 173596 29820
rect 173540 29766 173542 29818
rect 173542 29766 173594 29818
rect 173594 29766 173596 29818
rect 173540 29764 173596 29766
rect 173644 29818 173700 29820
rect 173644 29766 173646 29818
rect 173646 29766 173698 29818
rect 173698 29766 173700 29818
rect 173644 29764 173700 29766
rect 173436 28250 173492 28252
rect 173436 28198 173438 28250
rect 173438 28198 173490 28250
rect 173490 28198 173492 28250
rect 173436 28196 173492 28198
rect 173540 28250 173596 28252
rect 173540 28198 173542 28250
rect 173542 28198 173594 28250
rect 173594 28198 173596 28250
rect 173540 28196 173596 28198
rect 173644 28250 173700 28252
rect 173644 28198 173646 28250
rect 173646 28198 173698 28250
rect 173698 28198 173700 28250
rect 173644 28196 173700 28198
rect 173436 26682 173492 26684
rect 173436 26630 173438 26682
rect 173438 26630 173490 26682
rect 173490 26630 173492 26682
rect 173436 26628 173492 26630
rect 173540 26682 173596 26684
rect 173540 26630 173542 26682
rect 173542 26630 173594 26682
rect 173594 26630 173596 26682
rect 173540 26628 173596 26630
rect 173644 26682 173700 26684
rect 173644 26630 173646 26682
rect 173646 26630 173698 26682
rect 173698 26630 173700 26682
rect 173644 26628 173700 26630
rect 173436 25114 173492 25116
rect 173436 25062 173438 25114
rect 173438 25062 173490 25114
rect 173490 25062 173492 25114
rect 173436 25060 173492 25062
rect 173540 25114 173596 25116
rect 173540 25062 173542 25114
rect 173542 25062 173594 25114
rect 173594 25062 173596 25114
rect 173540 25060 173596 25062
rect 173644 25114 173700 25116
rect 173644 25062 173646 25114
rect 173646 25062 173698 25114
rect 173698 25062 173700 25114
rect 173644 25060 173700 25062
rect 173436 23546 173492 23548
rect 173436 23494 173438 23546
rect 173438 23494 173490 23546
rect 173490 23494 173492 23546
rect 173436 23492 173492 23494
rect 173540 23546 173596 23548
rect 173540 23494 173542 23546
rect 173542 23494 173594 23546
rect 173594 23494 173596 23546
rect 173540 23492 173596 23494
rect 173644 23546 173700 23548
rect 173644 23494 173646 23546
rect 173646 23494 173698 23546
rect 173698 23494 173700 23546
rect 173644 23492 173700 23494
rect 173436 21978 173492 21980
rect 173436 21926 173438 21978
rect 173438 21926 173490 21978
rect 173490 21926 173492 21978
rect 173436 21924 173492 21926
rect 173540 21978 173596 21980
rect 173540 21926 173542 21978
rect 173542 21926 173594 21978
rect 173594 21926 173596 21978
rect 173540 21924 173596 21926
rect 173644 21978 173700 21980
rect 173644 21926 173646 21978
rect 173646 21926 173698 21978
rect 173698 21926 173700 21978
rect 173644 21924 173700 21926
rect 178892 20972 178948 21028
rect 173436 20410 173492 20412
rect 173436 20358 173438 20410
rect 173438 20358 173490 20410
rect 173490 20358 173492 20410
rect 173436 20356 173492 20358
rect 173540 20410 173596 20412
rect 173540 20358 173542 20410
rect 173542 20358 173594 20410
rect 173594 20358 173596 20410
rect 173540 20356 173596 20358
rect 173644 20410 173700 20412
rect 173644 20358 173646 20410
rect 173646 20358 173698 20410
rect 173698 20358 173700 20410
rect 173644 20356 173700 20358
rect 173436 18842 173492 18844
rect 173436 18790 173438 18842
rect 173438 18790 173490 18842
rect 173490 18790 173492 18842
rect 173436 18788 173492 18790
rect 173540 18842 173596 18844
rect 173540 18790 173542 18842
rect 173542 18790 173594 18842
rect 173594 18790 173596 18842
rect 173540 18788 173596 18790
rect 173644 18842 173700 18844
rect 173644 18790 173646 18842
rect 173646 18790 173698 18842
rect 173698 18790 173700 18842
rect 173644 18788 173700 18790
rect 173436 17274 173492 17276
rect 173436 17222 173438 17274
rect 173438 17222 173490 17274
rect 173490 17222 173492 17274
rect 173436 17220 173492 17222
rect 173540 17274 173596 17276
rect 173540 17222 173542 17274
rect 173542 17222 173594 17274
rect 173594 17222 173596 17274
rect 173540 17220 173596 17222
rect 173644 17274 173700 17276
rect 173644 17222 173646 17274
rect 173646 17222 173698 17274
rect 173698 17222 173700 17274
rect 173644 17220 173700 17222
rect 173436 15706 173492 15708
rect 173436 15654 173438 15706
rect 173438 15654 173490 15706
rect 173490 15654 173492 15706
rect 173436 15652 173492 15654
rect 173540 15706 173596 15708
rect 173540 15654 173542 15706
rect 173542 15654 173594 15706
rect 173594 15654 173596 15706
rect 173540 15652 173596 15654
rect 173644 15706 173700 15708
rect 173644 15654 173646 15706
rect 173646 15654 173698 15706
rect 173698 15654 173700 15706
rect 173644 15652 173700 15654
rect 173436 14138 173492 14140
rect 173436 14086 173438 14138
rect 173438 14086 173490 14138
rect 173490 14086 173492 14138
rect 173436 14084 173492 14086
rect 173540 14138 173596 14140
rect 173540 14086 173542 14138
rect 173542 14086 173594 14138
rect 173594 14086 173596 14138
rect 173540 14084 173596 14086
rect 173644 14138 173700 14140
rect 173644 14086 173646 14138
rect 173646 14086 173698 14138
rect 173698 14086 173700 14138
rect 173644 14084 173700 14086
rect 173436 12570 173492 12572
rect 173436 12518 173438 12570
rect 173438 12518 173490 12570
rect 173490 12518 173492 12570
rect 173436 12516 173492 12518
rect 173540 12570 173596 12572
rect 173540 12518 173542 12570
rect 173542 12518 173594 12570
rect 173594 12518 173596 12570
rect 173540 12516 173596 12518
rect 173644 12570 173700 12572
rect 173644 12518 173646 12570
rect 173646 12518 173698 12570
rect 173698 12518 173700 12570
rect 173644 12516 173700 12518
rect 171948 11228 172004 11284
rect 111996 11002 112052 11004
rect 111996 10950 111998 11002
rect 111998 10950 112050 11002
rect 112050 10950 112052 11002
rect 111996 10948 112052 10950
rect 112100 11002 112156 11004
rect 112100 10950 112102 11002
rect 112102 10950 112154 11002
rect 112154 10950 112156 11002
rect 112100 10948 112156 10950
rect 112204 11002 112260 11004
rect 112204 10950 112206 11002
rect 112206 10950 112258 11002
rect 112258 10950 112260 11002
rect 112204 10948 112260 10950
rect 142716 11002 142772 11004
rect 142716 10950 142718 11002
rect 142718 10950 142770 11002
rect 142770 10950 142772 11002
rect 142716 10948 142772 10950
rect 142820 11002 142876 11004
rect 142820 10950 142822 11002
rect 142822 10950 142874 11002
rect 142874 10950 142876 11002
rect 142820 10948 142876 10950
rect 142924 11002 142980 11004
rect 142924 10950 142926 11002
rect 142926 10950 142978 11002
rect 142978 10950 142980 11002
rect 142924 10948 142980 10950
rect 173436 11002 173492 11004
rect 173436 10950 173438 11002
rect 173438 10950 173490 11002
rect 173490 10950 173492 11002
rect 173436 10948 173492 10950
rect 173540 11002 173596 11004
rect 173540 10950 173542 11002
rect 173542 10950 173594 11002
rect 173594 10950 173596 11002
rect 173540 10948 173596 10950
rect 173644 11002 173700 11004
rect 173644 10950 173646 11002
rect 173646 10950 173698 11002
rect 173698 10950 173700 11002
rect 173644 10948 173700 10950
rect 127356 10218 127412 10220
rect 127356 10166 127358 10218
rect 127358 10166 127410 10218
rect 127410 10166 127412 10218
rect 127356 10164 127412 10166
rect 127460 10218 127516 10220
rect 127460 10166 127462 10218
rect 127462 10166 127514 10218
rect 127514 10166 127516 10218
rect 127460 10164 127516 10166
rect 127564 10218 127620 10220
rect 127564 10166 127566 10218
rect 127566 10166 127618 10218
rect 127618 10166 127620 10218
rect 127564 10164 127620 10166
rect 158076 10218 158132 10220
rect 158076 10166 158078 10218
rect 158078 10166 158130 10218
rect 158130 10166 158132 10218
rect 158076 10164 158132 10166
rect 158180 10218 158236 10220
rect 158180 10166 158182 10218
rect 158182 10166 158234 10218
rect 158234 10166 158236 10218
rect 158180 10164 158236 10166
rect 158284 10218 158340 10220
rect 158284 10166 158286 10218
rect 158286 10166 158338 10218
rect 158338 10166 158340 10218
rect 158284 10164 158340 10166
rect 111996 9434 112052 9436
rect 111996 9382 111998 9434
rect 111998 9382 112050 9434
rect 112050 9382 112052 9434
rect 111996 9380 112052 9382
rect 112100 9434 112156 9436
rect 112100 9382 112102 9434
rect 112102 9382 112154 9434
rect 112154 9382 112156 9434
rect 112100 9380 112156 9382
rect 112204 9434 112260 9436
rect 112204 9382 112206 9434
rect 112206 9382 112258 9434
rect 112258 9382 112260 9434
rect 112204 9380 112260 9382
rect 142716 9434 142772 9436
rect 142716 9382 142718 9434
rect 142718 9382 142770 9434
rect 142770 9382 142772 9434
rect 142716 9380 142772 9382
rect 142820 9434 142876 9436
rect 142820 9382 142822 9434
rect 142822 9382 142874 9434
rect 142874 9382 142876 9434
rect 142820 9380 142876 9382
rect 142924 9434 142980 9436
rect 142924 9382 142926 9434
rect 142926 9382 142978 9434
rect 142978 9382 142980 9434
rect 142924 9380 142980 9382
rect 173436 9434 173492 9436
rect 173436 9382 173438 9434
rect 173438 9382 173490 9434
rect 173490 9382 173492 9434
rect 173436 9380 173492 9382
rect 173540 9434 173596 9436
rect 173540 9382 173542 9434
rect 173542 9382 173594 9434
rect 173594 9382 173596 9434
rect 173540 9380 173596 9382
rect 173644 9434 173700 9436
rect 173644 9382 173646 9434
rect 173646 9382 173698 9434
rect 173698 9382 173700 9434
rect 173644 9380 173700 9382
rect 99932 9212 99988 9268
rect 119196 9100 119252 9156
rect 96636 8650 96692 8652
rect 96636 8598 96638 8650
rect 96638 8598 96690 8650
rect 96690 8598 96692 8650
rect 96636 8596 96692 8598
rect 96740 8650 96796 8652
rect 96740 8598 96742 8650
rect 96742 8598 96794 8650
rect 96794 8598 96796 8650
rect 96740 8596 96796 8598
rect 96844 8650 96900 8652
rect 96844 8598 96846 8650
rect 96846 8598 96898 8650
rect 96898 8598 96900 8650
rect 96844 8596 96900 8598
rect 111996 7866 112052 7868
rect 111996 7814 111998 7866
rect 111998 7814 112050 7866
rect 112050 7814 112052 7866
rect 111996 7812 112052 7814
rect 112100 7866 112156 7868
rect 112100 7814 112102 7866
rect 112102 7814 112154 7866
rect 112154 7814 112156 7866
rect 112100 7812 112156 7814
rect 112204 7866 112260 7868
rect 112204 7814 112206 7866
rect 112206 7814 112258 7866
rect 112258 7814 112260 7866
rect 112204 7812 112260 7814
rect 96636 7082 96692 7084
rect 96636 7030 96638 7082
rect 96638 7030 96690 7082
rect 96690 7030 96692 7082
rect 96636 7028 96692 7030
rect 96740 7082 96796 7084
rect 96740 7030 96742 7082
rect 96742 7030 96794 7082
rect 96794 7030 96796 7082
rect 96740 7028 96796 7030
rect 96844 7082 96900 7084
rect 96844 7030 96846 7082
rect 96846 7030 96898 7082
rect 96898 7030 96900 7082
rect 96844 7028 96900 7030
rect 111996 6298 112052 6300
rect 111996 6246 111998 6298
rect 111998 6246 112050 6298
rect 112050 6246 112052 6298
rect 111996 6244 112052 6246
rect 112100 6298 112156 6300
rect 112100 6246 112102 6298
rect 112102 6246 112154 6298
rect 112154 6246 112156 6298
rect 112100 6244 112156 6246
rect 112204 6298 112260 6300
rect 112204 6246 112206 6298
rect 112206 6246 112258 6298
rect 112258 6246 112260 6298
rect 112204 6244 112260 6246
rect 93548 5852 93604 5908
rect 96636 5514 96692 5516
rect 96636 5462 96638 5514
rect 96638 5462 96690 5514
rect 96690 5462 96692 5514
rect 96636 5460 96692 5462
rect 96740 5514 96796 5516
rect 96740 5462 96742 5514
rect 96742 5462 96794 5514
rect 96794 5462 96796 5514
rect 96740 5460 96796 5462
rect 96844 5514 96900 5516
rect 96844 5462 96846 5514
rect 96846 5462 96898 5514
rect 96898 5462 96900 5514
rect 96844 5460 96900 5462
rect 91644 4508 91700 4564
rect 111996 4730 112052 4732
rect 111996 4678 111998 4730
rect 111998 4678 112050 4730
rect 112050 4678 112052 4730
rect 111996 4676 112052 4678
rect 112100 4730 112156 4732
rect 112100 4678 112102 4730
rect 112102 4678 112154 4730
rect 112154 4678 112156 4730
rect 112100 4676 112156 4678
rect 112204 4730 112260 4732
rect 112204 4678 112206 4730
rect 112206 4678 112258 4730
rect 112258 4678 112260 4730
rect 112204 4676 112260 4678
rect 96236 4562 96292 4564
rect 96236 4510 96238 4562
rect 96238 4510 96290 4562
rect 96290 4510 96292 4562
rect 96236 4508 96292 4510
rect 89628 4284 89684 4340
rect 89068 4226 89124 4228
rect 89068 4174 89070 4226
rect 89070 4174 89122 4226
rect 89122 4174 89124 4226
rect 89068 4172 89124 4174
rect 88732 3500 88788 3556
rect 89404 3554 89460 3556
rect 89404 3502 89406 3554
rect 89406 3502 89458 3554
rect 89458 3502 89460 3554
rect 89404 3500 89460 3502
rect 90972 4338 91028 4340
rect 90972 4286 90974 4338
rect 90974 4286 91026 4338
rect 91026 4286 91028 4338
rect 90972 4284 91028 4286
rect 90748 4060 90804 4116
rect 91980 4114 92036 4116
rect 91980 4062 91982 4114
rect 91982 4062 92034 4114
rect 92034 4062 92036 4114
rect 91980 4060 92036 4062
rect 96796 4450 96852 4452
rect 96796 4398 96798 4450
rect 96798 4398 96850 4450
rect 96850 4398 96852 4450
rect 96796 4396 96852 4398
rect 97580 4396 97636 4452
rect 96636 3946 96692 3948
rect 96636 3894 96638 3946
rect 96638 3894 96690 3946
rect 96690 3894 96692 3946
rect 96636 3892 96692 3894
rect 96740 3946 96796 3948
rect 96740 3894 96742 3946
rect 96742 3894 96794 3946
rect 96794 3894 96796 3946
rect 96740 3892 96796 3894
rect 96844 3946 96900 3948
rect 96844 3894 96846 3946
rect 96846 3894 96898 3946
rect 96898 3894 96900 3946
rect 96844 3892 96900 3894
rect 103964 3388 104020 3444
rect 104748 3442 104804 3444
rect 104748 3390 104750 3442
rect 104750 3390 104802 3442
rect 104802 3390 104804 3442
rect 104748 3388 104804 3390
rect 107772 3388 107828 3444
rect 108556 3442 108612 3444
rect 108556 3390 108558 3442
rect 108558 3390 108610 3442
rect 108610 3390 108612 3442
rect 108556 3388 108612 3390
rect 111468 3554 111524 3556
rect 111468 3502 111470 3554
rect 111470 3502 111522 3554
rect 111522 3502 111524 3554
rect 111468 3500 111524 3502
rect 111804 3500 111860 3556
rect 109340 3388 109396 3444
rect 111996 3162 112052 3164
rect 111996 3110 111998 3162
rect 111998 3110 112050 3162
rect 112050 3110 112052 3162
rect 111996 3108 112052 3110
rect 112100 3162 112156 3164
rect 112100 3110 112102 3162
rect 112102 3110 112154 3162
rect 112154 3110 112156 3162
rect 112100 3108 112156 3110
rect 112204 3162 112260 3164
rect 112204 3110 112206 3162
rect 112206 3110 112258 3162
rect 112258 3110 112260 3162
rect 112204 3108 112260 3110
rect 112812 3500 112868 3556
rect 115052 3554 115108 3556
rect 115052 3502 115054 3554
rect 115054 3502 115106 3554
rect 115106 3502 115108 3554
rect 115052 3500 115108 3502
rect 127356 8650 127412 8652
rect 127356 8598 127358 8650
rect 127358 8598 127410 8650
rect 127410 8598 127412 8650
rect 127356 8596 127412 8598
rect 127460 8650 127516 8652
rect 127460 8598 127462 8650
rect 127462 8598 127514 8650
rect 127514 8598 127516 8650
rect 127460 8596 127516 8598
rect 127564 8650 127620 8652
rect 127564 8598 127566 8650
rect 127566 8598 127618 8650
rect 127618 8598 127620 8650
rect 127564 8596 127620 8598
rect 158076 8650 158132 8652
rect 158076 8598 158078 8650
rect 158078 8598 158130 8650
rect 158130 8598 158132 8650
rect 158076 8596 158132 8598
rect 158180 8650 158236 8652
rect 158180 8598 158182 8650
rect 158182 8598 158234 8650
rect 158234 8598 158236 8650
rect 158180 8596 158236 8598
rect 158284 8650 158340 8652
rect 158284 8598 158286 8650
rect 158286 8598 158338 8650
rect 158338 8598 158340 8650
rect 158284 8596 158340 8598
rect 142716 7866 142772 7868
rect 142716 7814 142718 7866
rect 142718 7814 142770 7866
rect 142770 7814 142772 7866
rect 142716 7812 142772 7814
rect 142820 7866 142876 7868
rect 142820 7814 142822 7866
rect 142822 7814 142874 7866
rect 142874 7814 142876 7866
rect 142820 7812 142876 7814
rect 142924 7866 142980 7868
rect 142924 7814 142926 7866
rect 142926 7814 142978 7866
rect 142978 7814 142980 7866
rect 142924 7812 142980 7814
rect 173436 7866 173492 7868
rect 173436 7814 173438 7866
rect 173438 7814 173490 7866
rect 173490 7814 173492 7866
rect 173436 7812 173492 7814
rect 173540 7866 173596 7868
rect 173540 7814 173542 7866
rect 173542 7814 173594 7866
rect 173594 7814 173596 7866
rect 173540 7812 173596 7814
rect 173644 7866 173700 7868
rect 173644 7814 173646 7866
rect 173646 7814 173698 7866
rect 173698 7814 173700 7866
rect 173644 7812 173700 7814
rect 137900 7644 137956 7700
rect 127356 7082 127412 7084
rect 127356 7030 127358 7082
rect 127358 7030 127410 7082
rect 127410 7030 127412 7082
rect 127356 7028 127412 7030
rect 127460 7082 127516 7084
rect 127460 7030 127462 7082
rect 127462 7030 127514 7082
rect 127514 7030 127516 7082
rect 127460 7028 127516 7030
rect 127564 7082 127620 7084
rect 127564 7030 127566 7082
rect 127566 7030 127618 7082
rect 127618 7030 127620 7082
rect 127564 7028 127620 7030
rect 127356 5514 127412 5516
rect 127356 5462 127358 5514
rect 127358 5462 127410 5514
rect 127410 5462 127412 5514
rect 127356 5460 127412 5462
rect 127460 5514 127516 5516
rect 127460 5462 127462 5514
rect 127462 5462 127514 5514
rect 127514 5462 127516 5514
rect 127460 5460 127516 5462
rect 127564 5514 127620 5516
rect 127564 5462 127566 5514
rect 127566 5462 127618 5514
rect 127618 5462 127620 5514
rect 127564 5460 127620 5462
rect 122556 5068 122612 5124
rect 115388 3500 115444 3556
rect 112812 2268 112868 2324
rect 109340 1036 109396 1092
rect 134316 4844 134372 4900
rect 123900 4060 123956 4116
rect 127356 3946 127412 3948
rect 127356 3894 127358 3946
rect 127358 3894 127410 3946
rect 127410 3894 127412 3946
rect 127356 3892 127412 3894
rect 127460 3946 127516 3948
rect 127460 3894 127462 3946
rect 127462 3894 127514 3946
rect 127514 3894 127516 3946
rect 127460 3892 127516 3894
rect 127564 3946 127620 3948
rect 127564 3894 127566 3946
rect 127566 3894 127618 3946
rect 127618 3894 127620 3946
rect 127564 3892 127620 3894
rect 131516 3724 131572 3780
rect 124348 3500 124404 3556
rect 127708 3500 127764 3556
rect 124348 1484 124404 1540
rect 158076 7082 158132 7084
rect 158076 7030 158078 7082
rect 158078 7030 158130 7082
rect 158130 7030 158132 7082
rect 158076 7028 158132 7030
rect 158180 7082 158236 7084
rect 158180 7030 158182 7082
rect 158182 7030 158234 7082
rect 158234 7030 158236 7082
rect 158180 7028 158236 7030
rect 158284 7082 158340 7084
rect 158284 7030 158286 7082
rect 158286 7030 158338 7082
rect 158338 7030 158340 7082
rect 158284 7028 158340 7030
rect 145068 6860 145124 6916
rect 142716 6298 142772 6300
rect 142716 6246 142718 6298
rect 142718 6246 142770 6298
rect 142770 6246 142772 6298
rect 142716 6244 142772 6246
rect 142820 6298 142876 6300
rect 142820 6246 142822 6298
rect 142822 6246 142874 6298
rect 142874 6246 142876 6298
rect 142820 6244 142876 6246
rect 142924 6298 142980 6300
rect 142924 6246 142926 6298
rect 142926 6246 142978 6298
rect 142978 6246 142980 6298
rect 142924 6244 142980 6246
rect 141484 6076 141540 6132
rect 142716 4730 142772 4732
rect 142716 4678 142718 4730
rect 142718 4678 142770 4730
rect 142770 4678 142772 4730
rect 142716 4676 142772 4678
rect 142820 4730 142876 4732
rect 142820 4678 142822 4730
rect 142822 4678 142874 4730
rect 142874 4678 142876 4730
rect 142820 4676 142876 4678
rect 142924 4730 142980 4732
rect 142924 4678 142926 4730
rect 142926 4678 142978 4730
rect 142978 4678 142980 4730
rect 142924 4676 142980 4678
rect 142716 3162 142772 3164
rect 142716 3110 142718 3162
rect 142718 3110 142770 3162
rect 142770 3110 142772 3162
rect 142716 3108 142772 3110
rect 142820 3162 142876 3164
rect 142820 3110 142822 3162
rect 142822 3110 142874 3162
rect 142874 3110 142876 3162
rect 142820 3108 142876 3110
rect 142924 3162 142980 3164
rect 142924 3110 142926 3162
rect 142926 3110 142978 3162
rect 142978 3110 142980 3162
rect 142924 3108 142980 3110
rect 148652 6412 148708 6468
rect 173436 6298 173492 6300
rect 173436 6246 173438 6298
rect 173438 6246 173490 6298
rect 173490 6246 173492 6298
rect 173436 6244 173492 6246
rect 173540 6298 173596 6300
rect 173540 6246 173542 6298
rect 173542 6246 173594 6298
rect 173594 6246 173596 6298
rect 173540 6244 173596 6246
rect 173644 6298 173700 6300
rect 173644 6246 173646 6298
rect 173646 6246 173698 6298
rect 173698 6246 173700 6298
rect 173644 6244 173700 6246
rect 158076 5514 158132 5516
rect 158076 5462 158078 5514
rect 158078 5462 158130 5514
rect 158130 5462 158132 5514
rect 158076 5460 158132 5462
rect 158180 5514 158236 5516
rect 158180 5462 158182 5514
rect 158182 5462 158234 5514
rect 158234 5462 158236 5514
rect 158180 5460 158236 5462
rect 158284 5514 158340 5516
rect 158284 5462 158286 5514
rect 158286 5462 158338 5514
rect 158338 5462 158340 5514
rect 158284 5460 158340 5462
rect 173436 4730 173492 4732
rect 173436 4678 173438 4730
rect 173438 4678 173490 4730
rect 173490 4678 173492 4730
rect 173436 4676 173492 4678
rect 173540 4730 173596 4732
rect 173540 4678 173542 4730
rect 173542 4678 173594 4730
rect 173594 4678 173596 4730
rect 173540 4676 173596 4678
rect 173644 4730 173700 4732
rect 173644 4678 173646 4730
rect 173646 4678 173698 4730
rect 173698 4678 173700 4730
rect 173644 4676 173700 4678
rect 173740 4508 173796 4564
rect 152236 4172 152292 4228
rect 158076 3946 158132 3948
rect 158076 3894 158078 3946
rect 158078 3894 158130 3946
rect 158130 3894 158132 3946
rect 158076 3892 158132 3894
rect 158180 3946 158236 3948
rect 158180 3894 158182 3946
rect 158182 3894 158234 3946
rect 158234 3894 158236 3946
rect 158180 3892 158236 3894
rect 158284 3946 158340 3948
rect 158284 3894 158286 3946
rect 158286 3894 158338 3946
rect 158338 3894 158340 3946
rect 158284 3892 158340 3894
rect 170156 3836 170212 3892
rect 156268 2380 156324 2436
rect 159628 1932 159684 1988
rect 162988 2828 163044 2884
rect 166572 3442 166628 3444
rect 166572 3390 166574 3442
rect 166574 3390 166626 3442
rect 166626 3390 166628 3442
rect 166572 3388 166628 3390
rect 169932 3388 169988 3444
rect 169932 2716 169988 2772
rect 173436 3162 173492 3164
rect 173436 3110 173438 3162
rect 173438 3110 173490 3162
rect 173490 3110 173492 3162
rect 173436 3108 173492 3110
rect 173540 3162 173596 3164
rect 173540 3110 173542 3162
rect 173542 3110 173594 3162
rect 173594 3110 173596 3162
rect 173540 3108 173596 3110
rect 173644 3162 173700 3164
rect 173644 3110 173646 3162
rect 173646 3110 173698 3162
rect 173698 3110 173700 3162
rect 173644 3108 173700 3110
rect 186172 52780 186228 52836
rect 187180 52834 187236 52836
rect 187180 52782 187182 52834
rect 187182 52782 187234 52834
rect 187234 52782 187236 52834
rect 187180 52780 187236 52782
rect 186172 52274 186228 52276
rect 186172 52222 186174 52274
rect 186174 52222 186226 52274
rect 186226 52222 186228 52274
rect 186172 52220 186228 52222
rect 185388 19292 185444 19348
rect 187292 49532 187348 49588
rect 183372 17612 183428 17668
rect 182252 15932 182308 15988
rect 182252 7532 182308 7588
rect 182364 5852 182420 5908
rect 181580 4060 181636 4116
rect 182252 4060 182308 4116
rect 182028 3724 182084 3780
rect 181020 3612 181076 3668
rect 178892 2492 178948 2548
rect 177324 1148 177380 1204
rect 184828 14252 184884 14308
rect 184492 7420 184548 7476
rect 184044 6466 184100 6468
rect 184044 6414 184046 6466
rect 184046 6414 184098 6466
rect 184098 6414 184100 6466
rect 184044 6412 184100 6414
rect 183708 5906 183764 5908
rect 183708 5854 183710 5906
rect 183710 5854 183762 5906
rect 183762 5854 183764 5906
rect 183708 5852 183764 5854
rect 184604 5906 184660 5908
rect 184604 5854 184606 5906
rect 184606 5854 184658 5906
rect 184658 5854 184660 5906
rect 184604 5852 184660 5854
rect 183596 4956 183652 5012
rect 184716 5292 184772 5348
rect 184604 4956 184660 5012
rect 182812 4338 182868 4340
rect 182812 4286 182814 4338
rect 182814 4286 182866 4338
rect 182866 4286 182868 4338
rect 182812 4284 182868 4286
rect 183708 4338 183764 4340
rect 183708 4286 183710 4338
rect 183710 4286 183762 4338
rect 183762 4286 183764 4338
rect 183708 4284 183764 4286
rect 185276 12684 185332 12740
rect 187292 8988 187348 9044
rect 190428 54460 190484 54516
rect 191436 54514 191492 54516
rect 191436 54462 191438 54514
rect 191438 54462 191490 54514
rect 191490 54462 191492 54514
rect 191436 54460 191492 54462
rect 188796 54122 188852 54124
rect 188796 54070 188798 54122
rect 188798 54070 188850 54122
rect 188850 54070 188852 54122
rect 188796 54068 188852 54070
rect 188900 54122 188956 54124
rect 188900 54070 188902 54122
rect 188902 54070 188954 54122
rect 188954 54070 188956 54122
rect 188900 54068 188956 54070
rect 189004 54122 189060 54124
rect 189004 54070 189006 54122
rect 189006 54070 189058 54122
rect 189058 54070 189060 54122
rect 189004 54068 189060 54070
rect 189756 53730 189812 53732
rect 189756 53678 189758 53730
rect 189758 53678 189810 53730
rect 189810 53678 189812 53730
rect 189756 53676 189812 53678
rect 195916 56194 195972 56196
rect 195916 56142 195918 56194
rect 195918 56142 195970 56194
rect 195970 56142 195972 56194
rect 195916 56140 195972 56142
rect 204156 56474 204212 56476
rect 204156 56422 204158 56474
rect 204158 56422 204210 56474
rect 204210 56422 204212 56474
rect 204156 56420 204212 56422
rect 204260 56474 204316 56476
rect 204260 56422 204262 56474
rect 204262 56422 204314 56474
rect 204314 56422 204316 56474
rect 204260 56420 204316 56422
rect 204364 56474 204420 56476
rect 204364 56422 204366 56474
rect 204366 56422 204418 56474
rect 204418 56422 204420 56474
rect 204364 56420 204420 56422
rect 206332 56252 206388 56308
rect 208348 56306 208404 56308
rect 208348 56254 208350 56306
rect 208350 56254 208402 56306
rect 208402 56254 208404 56306
rect 208348 56252 208404 56254
rect 202972 55916 203028 55972
rect 203756 55970 203812 55972
rect 203756 55918 203758 55970
rect 203758 55918 203810 55970
rect 203810 55918 203812 55970
rect 203756 55916 203812 55918
rect 205772 55916 205828 55972
rect 204156 54906 204212 54908
rect 204156 54854 204158 54906
rect 204158 54854 204210 54906
rect 204210 54854 204212 54906
rect 204156 54852 204212 54854
rect 204260 54906 204316 54908
rect 204260 54854 204262 54906
rect 204262 54854 204314 54906
rect 204314 54854 204316 54906
rect 204260 54852 204316 54854
rect 204364 54906 204420 54908
rect 204364 54854 204366 54906
rect 204366 54854 204418 54906
rect 204418 54854 204420 54906
rect 204364 54852 204420 54854
rect 194572 54514 194628 54516
rect 194572 54462 194574 54514
rect 194574 54462 194626 54514
rect 194626 54462 194628 54514
rect 194572 54460 194628 54462
rect 193228 53842 193284 53844
rect 193228 53790 193230 53842
rect 193230 53790 193282 53842
rect 193282 53790 193284 53842
rect 193228 53788 193284 53790
rect 195804 53788 195860 53844
rect 190428 53730 190484 53732
rect 190428 53678 190430 53730
rect 190430 53678 190482 53730
rect 190482 53678 190484 53730
rect 190428 53676 190484 53678
rect 189420 53506 189476 53508
rect 189420 53454 189422 53506
rect 189422 53454 189474 53506
rect 189474 53454 189476 53506
rect 189420 53452 189476 53454
rect 191100 53452 191156 53508
rect 188796 52554 188852 52556
rect 188796 52502 188798 52554
rect 188798 52502 188850 52554
rect 188850 52502 188852 52554
rect 188796 52500 188852 52502
rect 188900 52554 188956 52556
rect 188900 52502 188902 52554
rect 188902 52502 188954 52554
rect 188954 52502 188956 52554
rect 188900 52500 188956 52502
rect 189004 52554 189060 52556
rect 189004 52502 189006 52554
rect 189006 52502 189058 52554
rect 189058 52502 189060 52554
rect 189004 52500 189060 52502
rect 189308 52108 189364 52164
rect 190652 52108 190708 52164
rect 188796 50986 188852 50988
rect 188796 50934 188798 50986
rect 188798 50934 188850 50986
rect 188850 50934 188852 50986
rect 188796 50932 188852 50934
rect 188900 50986 188956 50988
rect 188900 50934 188902 50986
rect 188902 50934 188954 50986
rect 188954 50934 188956 50986
rect 188900 50932 188956 50934
rect 189004 50986 189060 50988
rect 189004 50934 189006 50986
rect 189006 50934 189058 50986
rect 189058 50934 189060 50986
rect 189004 50932 189060 50934
rect 188796 49418 188852 49420
rect 188796 49366 188798 49418
rect 188798 49366 188850 49418
rect 188850 49366 188852 49418
rect 188796 49364 188852 49366
rect 188900 49418 188956 49420
rect 188900 49366 188902 49418
rect 188902 49366 188954 49418
rect 188954 49366 188956 49418
rect 188900 49364 188956 49366
rect 189004 49418 189060 49420
rect 189004 49366 189006 49418
rect 189006 49366 189058 49418
rect 189058 49366 189060 49418
rect 189004 49364 189060 49366
rect 188796 47850 188852 47852
rect 188796 47798 188798 47850
rect 188798 47798 188850 47850
rect 188850 47798 188852 47850
rect 188796 47796 188852 47798
rect 188900 47850 188956 47852
rect 188900 47798 188902 47850
rect 188902 47798 188954 47850
rect 188954 47798 188956 47850
rect 188900 47796 188956 47798
rect 189004 47850 189060 47852
rect 189004 47798 189006 47850
rect 189006 47798 189058 47850
rect 189058 47798 189060 47850
rect 189004 47796 189060 47798
rect 188796 46282 188852 46284
rect 188796 46230 188798 46282
rect 188798 46230 188850 46282
rect 188850 46230 188852 46282
rect 188796 46228 188852 46230
rect 188900 46282 188956 46284
rect 188900 46230 188902 46282
rect 188902 46230 188954 46282
rect 188954 46230 188956 46282
rect 188900 46228 188956 46230
rect 189004 46282 189060 46284
rect 189004 46230 189006 46282
rect 189006 46230 189058 46282
rect 189058 46230 189060 46282
rect 189004 46228 189060 46230
rect 188796 44714 188852 44716
rect 188796 44662 188798 44714
rect 188798 44662 188850 44714
rect 188850 44662 188852 44714
rect 188796 44660 188852 44662
rect 188900 44714 188956 44716
rect 188900 44662 188902 44714
rect 188902 44662 188954 44714
rect 188954 44662 188956 44714
rect 188900 44660 188956 44662
rect 189004 44714 189060 44716
rect 189004 44662 189006 44714
rect 189006 44662 189058 44714
rect 189058 44662 189060 44714
rect 189004 44660 189060 44662
rect 188796 43146 188852 43148
rect 188796 43094 188798 43146
rect 188798 43094 188850 43146
rect 188850 43094 188852 43146
rect 188796 43092 188852 43094
rect 188900 43146 188956 43148
rect 188900 43094 188902 43146
rect 188902 43094 188954 43146
rect 188954 43094 188956 43146
rect 188900 43092 188956 43094
rect 189004 43146 189060 43148
rect 189004 43094 189006 43146
rect 189006 43094 189058 43146
rect 189058 43094 189060 43146
rect 189004 43092 189060 43094
rect 188796 41578 188852 41580
rect 188796 41526 188798 41578
rect 188798 41526 188850 41578
rect 188850 41526 188852 41578
rect 188796 41524 188852 41526
rect 188900 41578 188956 41580
rect 188900 41526 188902 41578
rect 188902 41526 188954 41578
rect 188954 41526 188956 41578
rect 188900 41524 188956 41526
rect 189004 41578 189060 41580
rect 189004 41526 189006 41578
rect 189006 41526 189058 41578
rect 189058 41526 189060 41578
rect 189004 41524 189060 41526
rect 188796 40010 188852 40012
rect 188796 39958 188798 40010
rect 188798 39958 188850 40010
rect 188850 39958 188852 40010
rect 188796 39956 188852 39958
rect 188900 40010 188956 40012
rect 188900 39958 188902 40010
rect 188902 39958 188954 40010
rect 188954 39958 188956 40010
rect 188900 39956 188956 39958
rect 189004 40010 189060 40012
rect 189004 39958 189006 40010
rect 189006 39958 189058 40010
rect 189058 39958 189060 40010
rect 189004 39956 189060 39958
rect 188796 38442 188852 38444
rect 188796 38390 188798 38442
rect 188798 38390 188850 38442
rect 188850 38390 188852 38442
rect 188796 38388 188852 38390
rect 188900 38442 188956 38444
rect 188900 38390 188902 38442
rect 188902 38390 188954 38442
rect 188954 38390 188956 38442
rect 188900 38388 188956 38390
rect 189004 38442 189060 38444
rect 189004 38390 189006 38442
rect 189006 38390 189058 38442
rect 189058 38390 189060 38442
rect 189004 38388 189060 38390
rect 188796 36874 188852 36876
rect 188796 36822 188798 36874
rect 188798 36822 188850 36874
rect 188850 36822 188852 36874
rect 188796 36820 188852 36822
rect 188900 36874 188956 36876
rect 188900 36822 188902 36874
rect 188902 36822 188954 36874
rect 188954 36822 188956 36874
rect 188900 36820 188956 36822
rect 189004 36874 189060 36876
rect 189004 36822 189006 36874
rect 189006 36822 189058 36874
rect 189058 36822 189060 36874
rect 189004 36820 189060 36822
rect 188796 35306 188852 35308
rect 188796 35254 188798 35306
rect 188798 35254 188850 35306
rect 188850 35254 188852 35306
rect 188796 35252 188852 35254
rect 188900 35306 188956 35308
rect 188900 35254 188902 35306
rect 188902 35254 188954 35306
rect 188954 35254 188956 35306
rect 188900 35252 188956 35254
rect 189004 35306 189060 35308
rect 189004 35254 189006 35306
rect 189006 35254 189058 35306
rect 189058 35254 189060 35306
rect 189004 35252 189060 35254
rect 188796 33738 188852 33740
rect 188796 33686 188798 33738
rect 188798 33686 188850 33738
rect 188850 33686 188852 33738
rect 188796 33684 188852 33686
rect 188900 33738 188956 33740
rect 188900 33686 188902 33738
rect 188902 33686 188954 33738
rect 188954 33686 188956 33738
rect 188900 33684 188956 33686
rect 189004 33738 189060 33740
rect 189004 33686 189006 33738
rect 189006 33686 189058 33738
rect 189058 33686 189060 33738
rect 189004 33684 189060 33686
rect 188796 32170 188852 32172
rect 188796 32118 188798 32170
rect 188798 32118 188850 32170
rect 188850 32118 188852 32170
rect 188796 32116 188852 32118
rect 188900 32170 188956 32172
rect 188900 32118 188902 32170
rect 188902 32118 188954 32170
rect 188954 32118 188956 32170
rect 188900 32116 188956 32118
rect 189004 32170 189060 32172
rect 189004 32118 189006 32170
rect 189006 32118 189058 32170
rect 189058 32118 189060 32170
rect 189004 32116 189060 32118
rect 188796 30602 188852 30604
rect 188796 30550 188798 30602
rect 188798 30550 188850 30602
rect 188850 30550 188852 30602
rect 188796 30548 188852 30550
rect 188900 30602 188956 30604
rect 188900 30550 188902 30602
rect 188902 30550 188954 30602
rect 188954 30550 188956 30602
rect 188900 30548 188956 30550
rect 189004 30602 189060 30604
rect 189004 30550 189006 30602
rect 189006 30550 189058 30602
rect 189058 30550 189060 30602
rect 189004 30548 189060 30550
rect 188796 29034 188852 29036
rect 188796 28982 188798 29034
rect 188798 28982 188850 29034
rect 188850 28982 188852 29034
rect 188796 28980 188852 28982
rect 188900 29034 188956 29036
rect 188900 28982 188902 29034
rect 188902 28982 188954 29034
rect 188954 28982 188956 29034
rect 188900 28980 188956 28982
rect 189004 29034 189060 29036
rect 189004 28982 189006 29034
rect 189006 28982 189058 29034
rect 189058 28982 189060 29034
rect 189004 28980 189060 28982
rect 188796 27466 188852 27468
rect 188796 27414 188798 27466
rect 188798 27414 188850 27466
rect 188850 27414 188852 27466
rect 188796 27412 188852 27414
rect 188900 27466 188956 27468
rect 188900 27414 188902 27466
rect 188902 27414 188954 27466
rect 188954 27414 188956 27466
rect 188900 27412 188956 27414
rect 189004 27466 189060 27468
rect 189004 27414 189006 27466
rect 189006 27414 189058 27466
rect 189058 27414 189060 27466
rect 189004 27412 189060 27414
rect 188796 25898 188852 25900
rect 188796 25846 188798 25898
rect 188798 25846 188850 25898
rect 188850 25846 188852 25898
rect 188796 25844 188852 25846
rect 188900 25898 188956 25900
rect 188900 25846 188902 25898
rect 188902 25846 188954 25898
rect 188954 25846 188956 25898
rect 188900 25844 188956 25846
rect 189004 25898 189060 25900
rect 189004 25846 189006 25898
rect 189006 25846 189058 25898
rect 189058 25846 189060 25898
rect 189004 25844 189060 25846
rect 188796 24330 188852 24332
rect 188796 24278 188798 24330
rect 188798 24278 188850 24330
rect 188850 24278 188852 24330
rect 188796 24276 188852 24278
rect 188900 24330 188956 24332
rect 188900 24278 188902 24330
rect 188902 24278 188954 24330
rect 188954 24278 188956 24330
rect 188900 24276 188956 24278
rect 189004 24330 189060 24332
rect 189004 24278 189006 24330
rect 189006 24278 189058 24330
rect 189058 24278 189060 24330
rect 189004 24276 189060 24278
rect 188796 22762 188852 22764
rect 188796 22710 188798 22762
rect 188798 22710 188850 22762
rect 188850 22710 188852 22762
rect 188796 22708 188852 22710
rect 188900 22762 188956 22764
rect 188900 22710 188902 22762
rect 188902 22710 188954 22762
rect 188954 22710 188956 22762
rect 188900 22708 188956 22710
rect 189004 22762 189060 22764
rect 189004 22710 189006 22762
rect 189006 22710 189058 22762
rect 189058 22710 189060 22762
rect 189004 22708 189060 22710
rect 188796 21194 188852 21196
rect 188796 21142 188798 21194
rect 188798 21142 188850 21194
rect 188850 21142 188852 21194
rect 188796 21140 188852 21142
rect 188900 21194 188956 21196
rect 188900 21142 188902 21194
rect 188902 21142 188954 21194
rect 188954 21142 188956 21194
rect 188900 21140 188956 21142
rect 189004 21194 189060 21196
rect 189004 21142 189006 21194
rect 189006 21142 189058 21194
rect 189058 21142 189060 21194
rect 189004 21140 189060 21142
rect 188796 19626 188852 19628
rect 188796 19574 188798 19626
rect 188798 19574 188850 19626
rect 188850 19574 188852 19626
rect 188796 19572 188852 19574
rect 188900 19626 188956 19628
rect 188900 19574 188902 19626
rect 188902 19574 188954 19626
rect 188954 19574 188956 19626
rect 188900 19572 188956 19574
rect 189004 19626 189060 19628
rect 189004 19574 189006 19626
rect 189006 19574 189058 19626
rect 189058 19574 189060 19626
rect 189004 19572 189060 19574
rect 188796 18058 188852 18060
rect 188796 18006 188798 18058
rect 188798 18006 188850 18058
rect 188850 18006 188852 18058
rect 188796 18004 188852 18006
rect 188900 18058 188956 18060
rect 188900 18006 188902 18058
rect 188902 18006 188954 18058
rect 188954 18006 188956 18058
rect 188900 18004 188956 18006
rect 189004 18058 189060 18060
rect 189004 18006 189006 18058
rect 189006 18006 189058 18058
rect 189058 18006 189060 18058
rect 189004 18004 189060 18006
rect 188796 16490 188852 16492
rect 188796 16438 188798 16490
rect 188798 16438 188850 16490
rect 188850 16438 188852 16490
rect 188796 16436 188852 16438
rect 188900 16490 188956 16492
rect 188900 16438 188902 16490
rect 188902 16438 188954 16490
rect 188954 16438 188956 16490
rect 188900 16436 188956 16438
rect 189004 16490 189060 16492
rect 189004 16438 189006 16490
rect 189006 16438 189058 16490
rect 189058 16438 189060 16490
rect 189004 16436 189060 16438
rect 188796 14922 188852 14924
rect 188796 14870 188798 14922
rect 188798 14870 188850 14922
rect 188850 14870 188852 14922
rect 188796 14868 188852 14870
rect 188900 14922 188956 14924
rect 188900 14870 188902 14922
rect 188902 14870 188954 14922
rect 188954 14870 188956 14922
rect 188900 14868 188956 14870
rect 189004 14922 189060 14924
rect 189004 14870 189006 14922
rect 189006 14870 189058 14922
rect 189058 14870 189060 14922
rect 189004 14868 189060 14870
rect 188796 13354 188852 13356
rect 188796 13302 188798 13354
rect 188798 13302 188850 13354
rect 188850 13302 188852 13354
rect 188796 13300 188852 13302
rect 188900 13354 188956 13356
rect 188900 13302 188902 13354
rect 188902 13302 188954 13354
rect 188954 13302 188956 13354
rect 188900 13300 188956 13302
rect 189004 13354 189060 13356
rect 189004 13302 189006 13354
rect 189006 13302 189058 13354
rect 189058 13302 189060 13354
rect 189004 13300 189060 13302
rect 188796 11786 188852 11788
rect 188796 11734 188798 11786
rect 188798 11734 188850 11786
rect 188850 11734 188852 11786
rect 188796 11732 188852 11734
rect 188900 11786 188956 11788
rect 188900 11734 188902 11786
rect 188902 11734 188954 11786
rect 188954 11734 188956 11786
rect 188900 11732 188956 11734
rect 189004 11786 189060 11788
rect 189004 11734 189006 11786
rect 189006 11734 189058 11786
rect 189058 11734 189060 11786
rect 189004 11732 189060 11734
rect 188796 10218 188852 10220
rect 188796 10166 188798 10218
rect 188798 10166 188850 10218
rect 188850 10166 188852 10218
rect 188796 10164 188852 10166
rect 188900 10218 188956 10220
rect 188900 10166 188902 10218
rect 188902 10166 188954 10218
rect 188954 10166 188956 10218
rect 188900 10164 188956 10166
rect 189004 10218 189060 10220
rect 189004 10166 189006 10218
rect 189006 10166 189058 10218
rect 189058 10166 189060 10218
rect 190652 10220 190708 10276
rect 191324 17612 191380 17668
rect 189004 10164 189060 10166
rect 188796 8650 188852 8652
rect 188796 8598 188798 8650
rect 188798 8598 188850 8650
rect 188850 8598 188852 8650
rect 188796 8596 188852 8598
rect 188900 8650 188956 8652
rect 188900 8598 188902 8650
rect 188902 8598 188954 8650
rect 188954 8598 188956 8650
rect 188900 8596 188956 8598
rect 189004 8650 189060 8652
rect 189004 8598 189006 8650
rect 189006 8598 189058 8650
rect 189058 8598 189060 8650
rect 189004 8596 189060 8598
rect 188636 8258 188692 8260
rect 188636 8206 188638 8258
rect 188638 8206 188690 8258
rect 188690 8206 188692 8258
rect 188636 8204 188692 8206
rect 189084 8258 189140 8260
rect 189084 8206 189086 8258
rect 189086 8206 189138 8258
rect 189138 8206 189140 8258
rect 189084 8204 189140 8206
rect 187628 7644 187684 7700
rect 185388 7586 185444 7588
rect 185388 7534 185390 7586
rect 185390 7534 185442 7586
rect 185442 7534 185444 7586
rect 185388 7532 185444 7534
rect 185612 7474 185668 7476
rect 185612 7422 185614 7474
rect 185614 7422 185666 7474
rect 185666 7422 185668 7474
rect 185612 7420 185668 7422
rect 186284 7420 186340 7476
rect 187516 7420 187572 7476
rect 186732 6860 186788 6916
rect 185388 5404 185444 5460
rect 185948 5234 186004 5236
rect 185948 5182 185950 5234
rect 185950 5182 186002 5234
rect 186002 5182 186004 5234
rect 185948 5180 186004 5182
rect 186732 5906 186788 5908
rect 186732 5854 186734 5906
rect 186734 5854 186786 5906
rect 186786 5854 186788 5906
rect 186732 5852 186788 5854
rect 186172 5068 186228 5124
rect 186396 5628 186452 5684
rect 187068 5404 187124 5460
rect 187516 6300 187572 6356
rect 187516 5964 187572 6020
rect 187404 5292 187460 5348
rect 186620 5010 186676 5012
rect 186620 4958 186622 5010
rect 186622 4958 186674 5010
rect 186674 4958 186676 5010
rect 186620 4956 186676 4958
rect 186172 4844 186228 4900
rect 183932 3724 183988 3780
rect 182812 3554 182868 3556
rect 182812 3502 182814 3554
rect 182814 3502 182866 3554
rect 182866 3502 182868 3554
rect 182812 3500 182868 3502
rect 186284 4172 186340 4228
rect 185948 3554 186004 3556
rect 185948 3502 185950 3554
rect 185950 3502 186002 3554
rect 186002 3502 186004 3554
rect 185948 3500 186004 3502
rect 184828 3330 184884 3332
rect 184828 3278 184830 3330
rect 184830 3278 184882 3330
rect 184882 3278 184884 3330
rect 184828 3276 184884 3278
rect 186732 3500 186788 3556
rect 186284 2604 186340 2660
rect 186844 2268 186900 2324
rect 187404 4898 187460 4900
rect 187404 4846 187406 4898
rect 187406 4846 187458 4898
rect 187458 4846 187460 4898
rect 187404 4844 187460 4846
rect 187852 7980 187908 8036
rect 188636 7644 188692 7700
rect 188076 7586 188132 7588
rect 188076 7534 188078 7586
rect 188078 7534 188130 7586
rect 188130 7534 188132 7586
rect 188076 7532 188132 7534
rect 189308 7644 189364 7700
rect 188300 7196 188356 7252
rect 188796 7082 188852 7084
rect 188796 7030 188798 7082
rect 188798 7030 188850 7082
rect 188850 7030 188852 7082
rect 188796 7028 188852 7030
rect 188900 7082 188956 7084
rect 188900 7030 188902 7082
rect 188902 7030 188954 7082
rect 188954 7030 188956 7082
rect 188900 7028 188956 7030
rect 189004 7082 189060 7084
rect 189004 7030 189006 7082
rect 189006 7030 189058 7082
rect 189058 7030 189060 7082
rect 189004 7028 189060 7030
rect 187964 6018 188020 6020
rect 187964 5966 187966 6018
rect 187966 5966 188018 6018
rect 188018 5966 188020 6018
rect 187964 5964 188020 5966
rect 187628 4956 187684 5012
rect 187964 4450 188020 4452
rect 187964 4398 187966 4450
rect 187966 4398 188018 4450
rect 188018 4398 188020 4450
rect 187964 4396 188020 4398
rect 187516 3724 187572 3780
rect 187068 2268 187124 2324
rect 187852 3442 187908 3444
rect 187852 3390 187854 3442
rect 187854 3390 187906 3442
rect 187906 3390 187908 3442
rect 187852 3388 187908 3390
rect 191100 8540 191156 8596
rect 189756 8370 189812 8372
rect 189756 8318 189758 8370
rect 189758 8318 189810 8370
rect 189810 8318 189812 8370
rect 189756 8316 189812 8318
rect 190764 8258 190820 8260
rect 190764 8206 190766 8258
rect 190766 8206 190818 8258
rect 190818 8206 190820 8258
rect 190764 8204 190820 8206
rect 190428 8034 190484 8036
rect 190428 7982 190430 8034
rect 190430 7982 190482 8034
rect 190482 7982 190484 8034
rect 190428 7980 190484 7982
rect 193228 15932 193284 15988
rect 192556 11116 192612 11172
rect 192668 9042 192724 9044
rect 192668 8990 192670 9042
rect 192670 8990 192722 9042
rect 192722 8990 192724 9042
rect 192668 8988 192724 8990
rect 191324 7644 191380 7700
rect 191100 7586 191156 7588
rect 191100 7534 191102 7586
rect 191102 7534 191154 7586
rect 191154 7534 191156 7586
rect 191100 7532 191156 7534
rect 190652 7474 190708 7476
rect 190652 7422 190654 7474
rect 190654 7422 190706 7474
rect 190706 7422 190708 7474
rect 190652 7420 190708 7422
rect 189868 7250 189924 7252
rect 189868 7198 189870 7250
rect 189870 7198 189922 7250
rect 189922 7198 189924 7250
rect 189868 7196 189924 7198
rect 190876 6748 190932 6804
rect 190316 6412 190372 6468
rect 189420 6300 189476 6356
rect 189196 5740 189252 5796
rect 188860 5628 188916 5684
rect 188796 5514 188852 5516
rect 188796 5462 188798 5514
rect 188798 5462 188850 5514
rect 188850 5462 188852 5514
rect 188796 5460 188852 5462
rect 188900 5514 188956 5516
rect 188900 5462 188902 5514
rect 188902 5462 188954 5514
rect 188954 5462 188956 5514
rect 188900 5460 188956 5462
rect 189004 5514 189060 5516
rect 189004 5462 189006 5514
rect 189006 5462 189058 5514
rect 189058 5462 189060 5514
rect 189004 5460 189060 5462
rect 188300 4396 188356 4452
rect 190428 5794 190484 5796
rect 190428 5742 190430 5794
rect 190430 5742 190482 5794
rect 190482 5742 190484 5794
rect 190428 5740 190484 5742
rect 190652 5628 190708 5684
rect 190316 5292 190372 5348
rect 189420 4620 189476 4676
rect 189868 5068 189924 5124
rect 190652 5180 190708 5236
rect 190316 4732 190372 4788
rect 188860 4396 188916 4452
rect 188796 3946 188852 3948
rect 188796 3894 188798 3946
rect 188798 3894 188850 3946
rect 188850 3894 188852 3946
rect 188796 3892 188852 3894
rect 188900 3946 188956 3948
rect 188900 3894 188902 3946
rect 188902 3894 188954 3946
rect 188954 3894 188956 3946
rect 188900 3892 188956 3894
rect 189004 3946 189060 3948
rect 189004 3894 189006 3946
rect 189006 3894 189058 3946
rect 189058 3894 189060 3946
rect 189004 3892 189060 3894
rect 189868 3612 189924 3668
rect 188524 3388 188580 3444
rect 190540 4450 190596 4452
rect 190540 4398 190542 4450
rect 190542 4398 190594 4450
rect 190594 4398 190596 4450
rect 190540 4396 190596 4398
rect 190988 6690 191044 6692
rect 190988 6638 190990 6690
rect 190990 6638 191042 6690
rect 191042 6638 191044 6690
rect 190988 6636 191044 6638
rect 192892 6748 192948 6804
rect 191660 6076 191716 6132
rect 191772 6018 191828 6020
rect 191772 5966 191774 6018
rect 191774 5966 191826 6018
rect 191826 5966 191828 6018
rect 191772 5964 191828 5966
rect 191100 5906 191156 5908
rect 191100 5854 191102 5906
rect 191102 5854 191154 5906
rect 191154 5854 191156 5906
rect 191100 5852 191156 5854
rect 192332 5740 192388 5796
rect 191660 5180 191716 5236
rect 190988 5122 191044 5124
rect 190988 5070 190990 5122
rect 190990 5070 191042 5122
rect 191042 5070 191044 5122
rect 190988 5068 191044 5070
rect 192332 5180 192388 5236
rect 192668 6524 192724 6580
rect 192780 6466 192836 6468
rect 192780 6414 192782 6466
rect 192782 6414 192834 6466
rect 192834 6414 192836 6466
rect 192780 6412 192836 6414
rect 192892 5964 192948 6020
rect 192668 5404 192724 5460
rect 195020 11116 195076 11172
rect 193564 9212 193620 9268
rect 193228 6690 193284 6692
rect 193228 6638 193230 6690
rect 193230 6638 193282 6690
rect 193282 6638 193284 6690
rect 193228 6636 193284 6638
rect 193340 7756 193396 7812
rect 193116 6412 193172 6468
rect 193900 7756 193956 7812
rect 193676 5180 193732 5236
rect 191660 4172 191716 4228
rect 192780 4060 192836 4116
rect 186732 2156 186788 2212
rect 193452 4338 193508 4340
rect 193452 4286 193454 4338
rect 193454 4286 193506 4338
rect 193506 4286 193508 4338
rect 193452 4284 193508 4286
rect 204156 53338 204212 53340
rect 204156 53286 204158 53338
rect 204158 53286 204210 53338
rect 204210 53286 204212 53338
rect 204156 53284 204212 53286
rect 204260 53338 204316 53340
rect 204260 53286 204262 53338
rect 204262 53286 204314 53338
rect 204314 53286 204316 53338
rect 204260 53284 204316 53286
rect 204364 53338 204420 53340
rect 204364 53286 204366 53338
rect 204366 53286 204418 53338
rect 204418 53286 204420 53338
rect 204364 53284 204420 53286
rect 204156 51770 204212 51772
rect 204156 51718 204158 51770
rect 204158 51718 204210 51770
rect 204210 51718 204212 51770
rect 204156 51716 204212 51718
rect 204260 51770 204316 51772
rect 204260 51718 204262 51770
rect 204262 51718 204314 51770
rect 204314 51718 204316 51770
rect 204260 51716 204316 51718
rect 204364 51770 204420 51772
rect 204364 51718 204366 51770
rect 204366 51718 204418 51770
rect 204418 51718 204420 51770
rect 204364 51716 204420 51718
rect 204156 50202 204212 50204
rect 204156 50150 204158 50202
rect 204158 50150 204210 50202
rect 204210 50150 204212 50202
rect 204156 50148 204212 50150
rect 204260 50202 204316 50204
rect 204260 50150 204262 50202
rect 204262 50150 204314 50202
rect 204314 50150 204316 50202
rect 204260 50148 204316 50150
rect 204364 50202 204420 50204
rect 204364 50150 204366 50202
rect 204366 50150 204418 50202
rect 204418 50150 204420 50202
rect 204364 50148 204420 50150
rect 204156 48634 204212 48636
rect 204156 48582 204158 48634
rect 204158 48582 204210 48634
rect 204210 48582 204212 48634
rect 204156 48580 204212 48582
rect 204260 48634 204316 48636
rect 204260 48582 204262 48634
rect 204262 48582 204314 48634
rect 204314 48582 204316 48634
rect 204260 48580 204316 48582
rect 204364 48634 204420 48636
rect 204364 48582 204366 48634
rect 204366 48582 204418 48634
rect 204418 48582 204420 48634
rect 204364 48580 204420 48582
rect 204156 47066 204212 47068
rect 204156 47014 204158 47066
rect 204158 47014 204210 47066
rect 204210 47014 204212 47066
rect 204156 47012 204212 47014
rect 204260 47066 204316 47068
rect 204260 47014 204262 47066
rect 204262 47014 204314 47066
rect 204314 47014 204316 47066
rect 204260 47012 204316 47014
rect 204364 47066 204420 47068
rect 204364 47014 204366 47066
rect 204366 47014 204418 47066
rect 204418 47014 204420 47066
rect 204364 47012 204420 47014
rect 204156 45498 204212 45500
rect 204156 45446 204158 45498
rect 204158 45446 204210 45498
rect 204210 45446 204212 45498
rect 204156 45444 204212 45446
rect 204260 45498 204316 45500
rect 204260 45446 204262 45498
rect 204262 45446 204314 45498
rect 204314 45446 204316 45498
rect 204260 45444 204316 45446
rect 204364 45498 204420 45500
rect 204364 45446 204366 45498
rect 204366 45446 204418 45498
rect 204418 45446 204420 45498
rect 204364 45444 204420 45446
rect 204156 43930 204212 43932
rect 204156 43878 204158 43930
rect 204158 43878 204210 43930
rect 204210 43878 204212 43930
rect 204156 43876 204212 43878
rect 204260 43930 204316 43932
rect 204260 43878 204262 43930
rect 204262 43878 204314 43930
rect 204314 43878 204316 43930
rect 204260 43876 204316 43878
rect 204364 43930 204420 43932
rect 204364 43878 204366 43930
rect 204366 43878 204418 43930
rect 204418 43878 204420 43930
rect 204364 43876 204420 43878
rect 204156 42362 204212 42364
rect 204156 42310 204158 42362
rect 204158 42310 204210 42362
rect 204210 42310 204212 42362
rect 204156 42308 204212 42310
rect 204260 42362 204316 42364
rect 204260 42310 204262 42362
rect 204262 42310 204314 42362
rect 204314 42310 204316 42362
rect 204260 42308 204316 42310
rect 204364 42362 204420 42364
rect 204364 42310 204366 42362
rect 204366 42310 204418 42362
rect 204418 42310 204420 42362
rect 204364 42308 204420 42310
rect 204156 40794 204212 40796
rect 204156 40742 204158 40794
rect 204158 40742 204210 40794
rect 204210 40742 204212 40794
rect 204156 40740 204212 40742
rect 204260 40794 204316 40796
rect 204260 40742 204262 40794
rect 204262 40742 204314 40794
rect 204314 40742 204316 40794
rect 204260 40740 204316 40742
rect 204364 40794 204420 40796
rect 204364 40742 204366 40794
rect 204366 40742 204418 40794
rect 204418 40742 204420 40794
rect 204364 40740 204420 40742
rect 204156 39226 204212 39228
rect 204156 39174 204158 39226
rect 204158 39174 204210 39226
rect 204210 39174 204212 39226
rect 204156 39172 204212 39174
rect 204260 39226 204316 39228
rect 204260 39174 204262 39226
rect 204262 39174 204314 39226
rect 204314 39174 204316 39226
rect 204260 39172 204316 39174
rect 204364 39226 204420 39228
rect 204364 39174 204366 39226
rect 204366 39174 204418 39226
rect 204418 39174 204420 39226
rect 204364 39172 204420 39174
rect 204156 37658 204212 37660
rect 204156 37606 204158 37658
rect 204158 37606 204210 37658
rect 204210 37606 204212 37658
rect 204156 37604 204212 37606
rect 204260 37658 204316 37660
rect 204260 37606 204262 37658
rect 204262 37606 204314 37658
rect 204314 37606 204316 37658
rect 204260 37604 204316 37606
rect 204364 37658 204420 37660
rect 204364 37606 204366 37658
rect 204366 37606 204418 37658
rect 204418 37606 204420 37658
rect 204364 37604 204420 37606
rect 204156 36090 204212 36092
rect 204156 36038 204158 36090
rect 204158 36038 204210 36090
rect 204210 36038 204212 36090
rect 204156 36036 204212 36038
rect 204260 36090 204316 36092
rect 204260 36038 204262 36090
rect 204262 36038 204314 36090
rect 204314 36038 204316 36090
rect 204260 36036 204316 36038
rect 204364 36090 204420 36092
rect 204364 36038 204366 36090
rect 204366 36038 204418 36090
rect 204418 36038 204420 36090
rect 204364 36036 204420 36038
rect 204156 34522 204212 34524
rect 204156 34470 204158 34522
rect 204158 34470 204210 34522
rect 204210 34470 204212 34522
rect 204156 34468 204212 34470
rect 204260 34522 204316 34524
rect 204260 34470 204262 34522
rect 204262 34470 204314 34522
rect 204314 34470 204316 34522
rect 204260 34468 204316 34470
rect 204364 34522 204420 34524
rect 204364 34470 204366 34522
rect 204366 34470 204418 34522
rect 204418 34470 204420 34522
rect 204364 34468 204420 34470
rect 204156 32954 204212 32956
rect 204156 32902 204158 32954
rect 204158 32902 204210 32954
rect 204210 32902 204212 32954
rect 204156 32900 204212 32902
rect 204260 32954 204316 32956
rect 204260 32902 204262 32954
rect 204262 32902 204314 32954
rect 204314 32902 204316 32954
rect 204260 32900 204316 32902
rect 204364 32954 204420 32956
rect 204364 32902 204366 32954
rect 204366 32902 204418 32954
rect 204418 32902 204420 32954
rect 204364 32900 204420 32902
rect 204156 31386 204212 31388
rect 204156 31334 204158 31386
rect 204158 31334 204210 31386
rect 204210 31334 204212 31386
rect 204156 31332 204212 31334
rect 204260 31386 204316 31388
rect 204260 31334 204262 31386
rect 204262 31334 204314 31386
rect 204314 31334 204316 31386
rect 204260 31332 204316 31334
rect 204364 31386 204420 31388
rect 204364 31334 204366 31386
rect 204366 31334 204418 31386
rect 204418 31334 204420 31386
rect 204364 31332 204420 31334
rect 205772 30268 205828 30324
rect 204156 29818 204212 29820
rect 204156 29766 204158 29818
rect 204158 29766 204210 29818
rect 204210 29766 204212 29818
rect 204156 29764 204212 29766
rect 204260 29818 204316 29820
rect 204260 29766 204262 29818
rect 204262 29766 204314 29818
rect 204314 29766 204316 29818
rect 204260 29764 204316 29766
rect 204364 29818 204420 29820
rect 204364 29766 204366 29818
rect 204366 29766 204418 29818
rect 204418 29766 204420 29818
rect 204364 29764 204420 29766
rect 204156 28250 204212 28252
rect 204156 28198 204158 28250
rect 204158 28198 204210 28250
rect 204210 28198 204212 28250
rect 204156 28196 204212 28198
rect 204260 28250 204316 28252
rect 204260 28198 204262 28250
rect 204262 28198 204314 28250
rect 204314 28198 204316 28250
rect 204260 28196 204316 28198
rect 204364 28250 204420 28252
rect 204364 28198 204366 28250
rect 204366 28198 204418 28250
rect 204418 28198 204420 28250
rect 204364 28196 204420 28198
rect 202300 27692 202356 27748
rect 198492 19292 198548 19348
rect 196700 14252 196756 14308
rect 195804 10108 195860 10164
rect 196140 10332 196196 10388
rect 195468 9884 195524 9940
rect 195356 7644 195412 7700
rect 195244 7532 195300 7588
rect 195020 5404 195076 5460
rect 194348 5068 194404 5124
rect 194572 5180 194628 5236
rect 195132 5068 195188 5124
rect 195244 6300 195300 6356
rect 195356 6076 195412 6132
rect 195244 5180 195300 5236
rect 194796 4844 194852 4900
rect 196028 9772 196084 9828
rect 196252 9996 196308 10052
rect 196028 6412 196084 6468
rect 196028 5906 196084 5908
rect 196028 5854 196030 5906
rect 196030 5854 196082 5906
rect 196082 5854 196084 5906
rect 196028 5852 196084 5854
rect 195468 5292 195524 5348
rect 196140 4898 196196 4900
rect 196140 4846 196142 4898
rect 196142 4846 196194 4898
rect 196194 4846 196196 4898
rect 196140 4844 196196 4846
rect 195804 4060 195860 4116
rect 195356 3554 195412 3556
rect 195356 3502 195358 3554
rect 195358 3502 195410 3554
rect 195410 3502 195412 3554
rect 195356 3500 195412 3502
rect 194684 3388 194740 3444
rect 193340 2492 193396 2548
rect 193004 1372 193060 1428
rect 195916 3442 195972 3444
rect 195916 3390 195918 3442
rect 195918 3390 195970 3442
rect 195970 3390 195972 3442
rect 195916 3388 195972 3390
rect 196364 4620 196420 4676
rect 197596 9212 197652 9268
rect 199164 10220 199220 10276
rect 199724 10108 199780 10164
rect 199724 9548 199780 9604
rect 198828 8316 198884 8372
rect 199052 8764 199108 8820
rect 200956 9602 201012 9604
rect 200956 9550 200958 9602
rect 200958 9550 201010 9602
rect 201010 9550 201012 9602
rect 200956 9548 201012 9550
rect 204156 26682 204212 26684
rect 204156 26630 204158 26682
rect 204158 26630 204210 26682
rect 204210 26630 204212 26682
rect 204156 26628 204212 26630
rect 204260 26682 204316 26684
rect 204260 26630 204262 26682
rect 204262 26630 204314 26682
rect 204314 26630 204316 26682
rect 204260 26628 204316 26630
rect 204364 26682 204420 26684
rect 204364 26630 204366 26682
rect 204366 26630 204418 26682
rect 204418 26630 204420 26682
rect 204364 26628 204420 26630
rect 204156 25114 204212 25116
rect 204156 25062 204158 25114
rect 204158 25062 204210 25114
rect 204210 25062 204212 25114
rect 204156 25060 204212 25062
rect 204260 25114 204316 25116
rect 204260 25062 204262 25114
rect 204262 25062 204314 25114
rect 204314 25062 204316 25114
rect 204260 25060 204316 25062
rect 204364 25114 204420 25116
rect 204364 25062 204366 25114
rect 204366 25062 204418 25114
rect 204418 25062 204420 25114
rect 204364 25060 204420 25062
rect 204156 23546 204212 23548
rect 204156 23494 204158 23546
rect 204158 23494 204210 23546
rect 204210 23494 204212 23546
rect 204156 23492 204212 23494
rect 204260 23546 204316 23548
rect 204260 23494 204262 23546
rect 204262 23494 204314 23546
rect 204314 23494 204316 23546
rect 204260 23492 204316 23494
rect 204364 23546 204420 23548
rect 204364 23494 204366 23546
rect 204366 23494 204418 23546
rect 204418 23494 204420 23546
rect 204364 23492 204420 23494
rect 204156 21978 204212 21980
rect 204156 21926 204158 21978
rect 204158 21926 204210 21978
rect 204210 21926 204212 21978
rect 204156 21924 204212 21926
rect 204260 21978 204316 21980
rect 204260 21926 204262 21978
rect 204262 21926 204314 21978
rect 204314 21926 204316 21978
rect 204260 21924 204316 21926
rect 204364 21978 204420 21980
rect 204364 21926 204366 21978
rect 204366 21926 204418 21978
rect 204418 21926 204420 21978
rect 204364 21924 204420 21926
rect 204156 20410 204212 20412
rect 204156 20358 204158 20410
rect 204158 20358 204210 20410
rect 204210 20358 204212 20410
rect 204156 20356 204212 20358
rect 204260 20410 204316 20412
rect 204260 20358 204262 20410
rect 204262 20358 204314 20410
rect 204314 20358 204316 20410
rect 204260 20356 204316 20358
rect 204364 20410 204420 20412
rect 204364 20358 204366 20410
rect 204366 20358 204418 20410
rect 204418 20358 204420 20410
rect 204364 20356 204420 20358
rect 204156 18842 204212 18844
rect 204156 18790 204158 18842
rect 204158 18790 204210 18842
rect 204210 18790 204212 18842
rect 204156 18788 204212 18790
rect 204260 18842 204316 18844
rect 204260 18790 204262 18842
rect 204262 18790 204314 18842
rect 204314 18790 204316 18842
rect 204260 18788 204316 18790
rect 204364 18842 204420 18844
rect 204364 18790 204366 18842
rect 204366 18790 204418 18842
rect 204418 18790 204420 18842
rect 204364 18788 204420 18790
rect 209132 55804 209188 55860
rect 206892 17612 206948 17668
rect 207900 20972 207956 21028
rect 204156 17274 204212 17276
rect 204156 17222 204158 17274
rect 204158 17222 204210 17274
rect 204210 17222 204212 17274
rect 204156 17220 204212 17222
rect 204260 17274 204316 17276
rect 204260 17222 204262 17274
rect 204262 17222 204314 17274
rect 204314 17222 204316 17274
rect 204260 17220 204316 17222
rect 204364 17274 204420 17276
rect 204364 17222 204366 17274
rect 204366 17222 204418 17274
rect 204418 17222 204420 17274
rect 204364 17220 204420 17222
rect 204156 15706 204212 15708
rect 204156 15654 204158 15706
rect 204158 15654 204210 15706
rect 204210 15654 204212 15706
rect 204156 15652 204212 15654
rect 204260 15706 204316 15708
rect 204260 15654 204262 15706
rect 204262 15654 204314 15706
rect 204314 15654 204316 15706
rect 204260 15652 204316 15654
rect 204364 15706 204420 15708
rect 204364 15654 204366 15706
rect 204366 15654 204418 15706
rect 204418 15654 204420 15706
rect 204364 15652 204420 15654
rect 204156 14138 204212 14140
rect 204156 14086 204158 14138
rect 204158 14086 204210 14138
rect 204210 14086 204212 14138
rect 204156 14084 204212 14086
rect 204260 14138 204316 14140
rect 204260 14086 204262 14138
rect 204262 14086 204314 14138
rect 204314 14086 204316 14138
rect 204260 14084 204316 14086
rect 204364 14138 204420 14140
rect 204364 14086 204366 14138
rect 204366 14086 204418 14138
rect 204418 14086 204420 14138
rect 204364 14084 204420 14086
rect 203644 12684 203700 12740
rect 202300 9266 202356 9268
rect 202300 9214 202302 9266
rect 202302 9214 202354 9266
rect 202354 9214 202356 9266
rect 202300 9212 202356 9214
rect 203084 9548 203140 9604
rect 204156 12570 204212 12572
rect 204156 12518 204158 12570
rect 204158 12518 204210 12570
rect 204210 12518 204212 12570
rect 204156 12516 204212 12518
rect 204260 12570 204316 12572
rect 204260 12518 204262 12570
rect 204262 12518 204314 12570
rect 204314 12518 204316 12570
rect 204260 12516 204316 12518
rect 204364 12570 204420 12572
rect 204364 12518 204366 12570
rect 204366 12518 204418 12570
rect 204418 12518 204420 12570
rect 204364 12516 204420 12518
rect 204156 11002 204212 11004
rect 204156 10950 204158 11002
rect 204158 10950 204210 11002
rect 204210 10950 204212 11002
rect 204156 10948 204212 10950
rect 204260 11002 204316 11004
rect 204260 10950 204262 11002
rect 204262 10950 204314 11002
rect 204314 10950 204316 11002
rect 204260 10948 204316 10950
rect 204364 11002 204420 11004
rect 204364 10950 204366 11002
rect 204366 10950 204418 11002
rect 204418 10950 204420 11002
rect 204364 10948 204420 10950
rect 204156 9434 204212 9436
rect 204156 9382 204158 9434
rect 204158 9382 204210 9434
rect 204210 9382 204212 9434
rect 204156 9380 204212 9382
rect 204260 9434 204316 9436
rect 204260 9382 204262 9434
rect 204262 9382 204314 9434
rect 204314 9382 204316 9434
rect 204260 9380 204316 9382
rect 204364 9434 204420 9436
rect 204364 9382 204366 9434
rect 204366 9382 204418 9434
rect 204418 9382 204420 9434
rect 204364 9380 204420 9382
rect 201292 8988 201348 9044
rect 199500 8764 199556 8820
rect 199612 8370 199668 8372
rect 199612 8318 199614 8370
rect 199614 8318 199666 8370
rect 199666 8318 199668 8370
rect 199612 8316 199668 8318
rect 200060 8146 200116 8148
rect 200060 8094 200062 8146
rect 200062 8094 200114 8146
rect 200114 8094 200116 8146
rect 200060 8092 200116 8094
rect 199724 7980 199780 8036
rect 199276 7420 199332 7476
rect 199388 7644 199444 7700
rect 198492 7308 198548 7364
rect 196812 5180 196868 5236
rect 197708 6130 197764 6132
rect 197708 6078 197710 6130
rect 197710 6078 197762 6130
rect 197762 6078 197764 6130
rect 197708 6076 197764 6078
rect 197596 5010 197652 5012
rect 197596 4958 197598 5010
rect 197598 4958 197650 5010
rect 197650 4958 197652 5010
rect 197596 4956 197652 4958
rect 197708 5068 197764 5124
rect 197148 4562 197204 4564
rect 197148 4510 197150 4562
rect 197150 4510 197202 4562
rect 197202 4510 197204 4562
rect 197148 4508 197204 4510
rect 199612 7196 199668 7252
rect 197932 4508 197988 4564
rect 198156 5628 198212 5684
rect 198156 4620 198212 4676
rect 196700 4396 196756 4452
rect 197708 4338 197764 4340
rect 197708 4286 197710 4338
rect 197710 4286 197762 4338
rect 197762 4286 197764 4338
rect 197708 4284 197764 4286
rect 197148 3442 197204 3444
rect 197148 3390 197150 3442
rect 197150 3390 197202 3442
rect 197202 3390 197204 3442
rect 197148 3388 197204 3390
rect 197596 3442 197652 3444
rect 197596 3390 197598 3442
rect 197598 3390 197650 3442
rect 197650 3390 197652 3442
rect 197596 3388 197652 3390
rect 199164 4956 199220 5012
rect 200844 8092 200900 8148
rect 200396 7474 200452 7476
rect 200396 7422 200398 7474
rect 200398 7422 200450 7474
rect 200450 7422 200452 7474
rect 200396 7420 200452 7422
rect 200956 7980 201012 8036
rect 200172 7250 200228 7252
rect 200172 7198 200174 7250
rect 200174 7198 200226 7250
rect 200226 7198 200228 7250
rect 200172 7196 200228 7198
rect 199836 6636 199892 6692
rect 199724 5964 199780 6020
rect 200620 5906 200676 5908
rect 200620 5854 200622 5906
rect 200622 5854 200674 5906
rect 200674 5854 200676 5906
rect 200620 5852 200676 5854
rect 199724 5740 199780 5796
rect 201180 6860 201236 6916
rect 200956 5404 201012 5460
rect 200844 5292 200900 5348
rect 199500 4508 199556 4564
rect 200620 4508 200676 4564
rect 199052 3612 199108 3668
rect 198716 3388 198772 3444
rect 198716 2828 198772 2884
rect 198716 2492 198772 2548
rect 200396 3442 200452 3444
rect 200396 3390 200398 3442
rect 200398 3390 200450 3442
rect 200450 3390 200452 3442
rect 200396 3388 200452 3390
rect 201068 5180 201124 5236
rect 203644 8988 203700 9044
rect 201852 8316 201908 8372
rect 203868 8764 203924 8820
rect 202972 8316 203028 8372
rect 202188 8146 202244 8148
rect 202188 8094 202190 8146
rect 202190 8094 202242 8146
rect 202242 8094 202244 8146
rect 202188 8092 202244 8094
rect 202412 8092 202468 8148
rect 202412 7420 202468 7476
rect 202972 7474 203028 7476
rect 202972 7422 202974 7474
rect 202974 7422 203026 7474
rect 203026 7422 203028 7474
rect 202972 7420 203028 7422
rect 202860 7308 202916 7364
rect 201628 6690 201684 6692
rect 201628 6638 201630 6690
rect 201630 6638 201682 6690
rect 201682 6638 201684 6690
rect 201628 6636 201684 6638
rect 203420 7980 203476 8036
rect 202860 6524 202916 6580
rect 202972 6636 203028 6692
rect 203084 6412 203140 6468
rect 203532 6130 203588 6132
rect 203532 6078 203534 6130
rect 203534 6078 203586 6130
rect 203586 6078 203588 6130
rect 203532 6076 203588 6078
rect 202972 5628 203028 5684
rect 201852 5180 201908 5236
rect 201740 5122 201796 5124
rect 201740 5070 201742 5122
rect 201742 5070 201794 5122
rect 201794 5070 201796 5122
rect 201740 5068 201796 5070
rect 201180 4172 201236 4228
rect 201292 3948 201348 4004
rect 200844 2716 200900 2772
rect 201292 3612 201348 3668
rect 201740 4396 201796 4452
rect 197596 2044 197652 2100
rect 195804 1596 195860 1652
rect 202972 5292 203028 5348
rect 202076 4396 202132 4452
rect 201852 3836 201908 3892
rect 201292 1260 201348 1316
rect 203980 8428 204036 8484
rect 205212 8316 205268 8372
rect 204156 7866 204212 7868
rect 204156 7814 204158 7866
rect 204158 7814 204210 7866
rect 204210 7814 204212 7866
rect 204156 7812 204212 7814
rect 204260 7866 204316 7868
rect 204260 7814 204262 7866
rect 204262 7814 204314 7866
rect 204314 7814 204316 7866
rect 204260 7812 204316 7814
rect 204364 7866 204420 7868
rect 204364 7814 204366 7866
rect 204366 7814 204418 7866
rect 204418 7814 204420 7866
rect 204364 7812 204420 7814
rect 204876 7980 204932 8036
rect 204652 7420 204708 7476
rect 204876 7362 204932 7364
rect 204876 7310 204878 7362
rect 204878 7310 204930 7362
rect 204930 7310 204932 7362
rect 204876 7308 204932 7310
rect 204988 6860 205044 6916
rect 204428 6636 204484 6692
rect 204652 6690 204708 6692
rect 204652 6638 204654 6690
rect 204654 6638 204706 6690
rect 204706 6638 204708 6690
rect 204652 6636 204708 6638
rect 204156 6298 204212 6300
rect 204156 6246 204158 6298
rect 204158 6246 204210 6298
rect 204210 6246 204212 6298
rect 204156 6244 204212 6246
rect 204260 6298 204316 6300
rect 204260 6246 204262 6298
rect 204262 6246 204314 6298
rect 204314 6246 204316 6298
rect 204260 6244 204316 6246
rect 204364 6298 204420 6300
rect 204364 6246 204366 6298
rect 204366 6246 204418 6298
rect 204418 6246 204420 6298
rect 204540 6300 204596 6356
rect 204364 6244 204420 6246
rect 203980 5794 204036 5796
rect 203980 5742 203982 5794
rect 203982 5742 204034 5794
rect 204034 5742 204036 5794
rect 203980 5740 204036 5742
rect 203868 5516 203924 5572
rect 203084 5068 203140 5124
rect 202972 4450 203028 4452
rect 202972 4398 202974 4450
rect 202974 4398 203026 4450
rect 203026 4398 203028 4450
rect 202972 4396 203028 4398
rect 202412 3554 202468 3556
rect 202412 3502 202414 3554
rect 202414 3502 202466 3554
rect 202466 3502 202468 3554
rect 202412 3500 202468 3502
rect 202748 3388 202804 3444
rect 203532 3554 203588 3556
rect 203532 3502 203534 3554
rect 203534 3502 203586 3554
rect 203586 3502 203588 3554
rect 203532 3500 203588 3502
rect 203980 5404 204036 5460
rect 204540 6076 204596 6132
rect 204764 6300 204820 6356
rect 205100 6578 205156 6580
rect 205100 6526 205102 6578
rect 205102 6526 205154 6578
rect 205154 6526 205156 6578
rect 205100 6524 205156 6526
rect 204652 5964 204708 6020
rect 204876 5852 204932 5908
rect 204092 4844 204148 4900
rect 204156 4730 204212 4732
rect 204156 4678 204158 4730
rect 204158 4678 204210 4730
rect 204210 4678 204212 4730
rect 204156 4676 204212 4678
rect 204260 4730 204316 4732
rect 204260 4678 204262 4730
rect 204262 4678 204314 4730
rect 204314 4678 204316 4730
rect 204260 4676 204316 4678
rect 204364 4730 204420 4732
rect 204364 4678 204366 4730
rect 204366 4678 204418 4730
rect 204418 4678 204420 4730
rect 204364 4676 204420 4678
rect 204540 4396 204596 4452
rect 204652 4844 204708 4900
rect 204540 4114 204596 4116
rect 204540 4062 204542 4114
rect 204542 4062 204594 4114
rect 204594 4062 204596 4114
rect 204540 4060 204596 4062
rect 204204 3724 204260 3780
rect 204988 5794 205044 5796
rect 204988 5742 204990 5794
rect 204990 5742 205042 5794
rect 205042 5742 205044 5794
rect 204988 5740 205044 5742
rect 205548 6076 205604 6132
rect 205212 5516 205268 5572
rect 205548 5740 205604 5796
rect 204156 3162 204212 3164
rect 204156 3110 204158 3162
rect 204158 3110 204210 3162
rect 204210 3110 204212 3162
rect 204156 3108 204212 3110
rect 204260 3162 204316 3164
rect 204260 3110 204262 3162
rect 204262 3110 204314 3162
rect 204314 3110 204316 3162
rect 204260 3108 204316 3110
rect 204364 3162 204420 3164
rect 204364 3110 204366 3162
rect 204366 3110 204418 3162
rect 204418 3110 204420 3162
rect 204364 3108 204420 3110
rect 205100 4396 205156 4452
rect 205324 4284 205380 4340
rect 205548 4338 205604 4340
rect 205548 4286 205550 4338
rect 205550 4286 205602 4338
rect 205602 4286 205604 4338
rect 205548 4284 205604 4286
rect 206332 8930 206388 8932
rect 206332 8878 206334 8930
rect 206334 8878 206386 8930
rect 206386 8878 206388 8930
rect 206332 8876 206388 8878
rect 207676 8876 207732 8932
rect 205884 8316 205940 8372
rect 205772 7980 205828 8036
rect 205996 8034 206052 8036
rect 205996 7982 205998 8034
rect 205998 7982 206050 8034
rect 206050 7982 206052 8034
rect 205996 7980 206052 7982
rect 206892 7756 206948 7812
rect 207340 8092 207396 8148
rect 206108 6972 206164 7028
rect 205772 5906 205828 5908
rect 205772 5854 205774 5906
rect 205774 5854 205826 5906
rect 205826 5854 205828 5906
rect 205772 5852 205828 5854
rect 205772 5516 205828 5572
rect 205660 3836 205716 3892
rect 206220 5628 206276 5684
rect 205996 5404 206052 5460
rect 207452 6690 207508 6692
rect 207452 6638 207454 6690
rect 207454 6638 207506 6690
rect 207506 6638 207508 6690
rect 207452 6636 207508 6638
rect 207004 6300 207060 6356
rect 208236 12796 208292 12852
rect 208124 8316 208180 8372
rect 207900 6466 207956 6468
rect 207900 6414 207902 6466
rect 207902 6414 207954 6466
rect 207954 6414 207956 6466
rect 207900 6412 207956 6414
rect 207452 5964 207508 6020
rect 206556 5906 206612 5908
rect 206556 5854 206558 5906
rect 206558 5854 206610 5906
rect 206610 5854 206612 5906
rect 206556 5852 206612 5854
rect 206332 5068 206388 5124
rect 205660 3666 205716 3668
rect 205660 3614 205662 3666
rect 205662 3614 205714 3666
rect 205714 3614 205716 3666
rect 205660 3612 205716 3614
rect 204764 2940 204820 2996
rect 204876 3442 204932 3444
rect 204876 3390 204878 3442
rect 204878 3390 204930 3442
rect 204930 3390 204932 3442
rect 204876 3388 204932 3390
rect 203196 2828 203252 2884
rect 203084 2716 203140 2772
rect 205660 3388 205716 3444
rect 204876 1932 204932 1988
rect 205996 5010 206052 5012
rect 205996 4958 205998 5010
rect 205998 4958 206050 5010
rect 206050 4958 206052 5010
rect 205996 4956 206052 4958
rect 206444 5740 206500 5796
rect 206556 5234 206612 5236
rect 206556 5182 206558 5234
rect 206558 5182 206610 5234
rect 206610 5182 206612 5234
rect 206556 5180 206612 5182
rect 206220 4898 206276 4900
rect 206220 4846 206222 4898
rect 206222 4846 206274 4898
rect 206274 4846 206276 4898
rect 206220 4844 206276 4846
rect 207340 5346 207396 5348
rect 207340 5294 207342 5346
rect 207342 5294 207394 5346
rect 207394 5294 207396 5346
rect 207340 5292 207396 5294
rect 207340 5068 207396 5124
rect 207228 5010 207284 5012
rect 207228 4958 207230 5010
rect 207230 4958 207282 5010
rect 207282 4958 207284 5010
rect 207228 4956 207284 4958
rect 207004 4898 207060 4900
rect 207004 4846 207006 4898
rect 207006 4846 207058 4898
rect 207058 4846 207060 4898
rect 207004 4844 207060 4846
rect 206220 4284 206276 4340
rect 205884 4172 205940 4228
rect 205772 2380 205828 2436
rect 206108 3836 206164 3892
rect 206668 3724 206724 3780
rect 205996 1148 206052 1204
rect 207564 5628 207620 5684
rect 210028 30268 210084 30324
rect 209916 9100 209972 9156
rect 209132 8876 209188 8932
rect 209468 8204 209524 8260
rect 209804 7756 209860 7812
rect 211932 11676 211988 11732
rect 210700 9660 210756 9716
rect 210700 9100 210756 9156
rect 210140 8204 210196 8260
rect 210364 8204 210420 8260
rect 211036 9714 211092 9716
rect 211036 9662 211038 9714
rect 211038 9662 211090 9714
rect 211090 9662 211092 9714
rect 211036 9660 211092 9662
rect 211260 9154 211316 9156
rect 211260 9102 211262 9154
rect 211262 9102 211314 9154
rect 211314 9102 211316 9154
rect 211260 9100 211316 9102
rect 209468 7420 209524 7476
rect 208012 4508 208068 4564
rect 207564 3388 207620 3444
rect 208124 3948 208180 4004
rect 208236 4732 208292 4788
rect 208348 4284 208404 4340
rect 209468 7084 209524 7140
rect 209468 5852 209524 5908
rect 210588 6748 210644 6804
rect 208796 5516 208852 5572
rect 209468 5122 209524 5124
rect 209468 5070 209470 5122
rect 209470 5070 209522 5122
rect 209522 5070 209524 5122
rect 209468 5068 209524 5070
rect 208908 4844 208964 4900
rect 209020 4284 209076 4340
rect 208460 3388 208516 3444
rect 209916 5068 209972 5124
rect 210364 5906 210420 5908
rect 210364 5854 210366 5906
rect 210366 5854 210418 5906
rect 210418 5854 210420 5906
rect 210364 5852 210420 5854
rect 211148 8258 211204 8260
rect 211148 8206 211150 8258
rect 211150 8206 211202 8258
rect 211202 8206 211204 8258
rect 211148 8204 211204 8206
rect 211708 9100 211764 9156
rect 212492 9548 212548 9604
rect 211372 8146 211428 8148
rect 211372 8094 211374 8146
rect 211374 8094 211426 8146
rect 211426 8094 211428 8146
rect 211372 8092 211428 8094
rect 211260 7980 211316 8036
rect 211932 8034 211988 8036
rect 211932 7982 211934 8034
rect 211934 7982 211986 8034
rect 211986 7982 211988 8034
rect 211932 7980 211988 7982
rect 212156 8316 212212 8372
rect 212156 7868 212212 7924
rect 211596 7586 211652 7588
rect 211596 7534 211598 7586
rect 211598 7534 211650 7586
rect 211650 7534 211652 7586
rect 211596 7532 211652 7534
rect 210924 7474 210980 7476
rect 210924 7422 210926 7474
rect 210926 7422 210978 7474
rect 210978 7422 210980 7474
rect 210924 7420 210980 7422
rect 211260 5906 211316 5908
rect 211260 5854 211262 5906
rect 211262 5854 211314 5906
rect 211314 5854 211316 5906
rect 211260 5852 211316 5854
rect 209804 4396 209860 4452
rect 210252 4844 210308 4900
rect 210028 4338 210084 4340
rect 210028 4286 210030 4338
rect 210030 4286 210082 4338
rect 210082 4286 210084 4338
rect 210028 4284 210084 4286
rect 209132 3388 209188 3444
rect 210028 3388 210084 3444
rect 208012 3164 208068 3220
rect 207340 2604 207396 2660
rect 206892 1036 206948 1092
rect 210700 5516 210756 5572
rect 211036 4732 211092 4788
rect 210812 4450 210868 4452
rect 210812 4398 210814 4450
rect 210814 4398 210866 4450
rect 210866 4398 210868 4450
rect 210812 4396 210868 4398
rect 211148 4284 211204 4340
rect 210588 3554 210644 3556
rect 210588 3502 210590 3554
rect 210590 3502 210642 3554
rect 210642 3502 210644 3554
rect 210588 3500 210644 3502
rect 211596 5404 211652 5460
rect 212380 8258 212436 8260
rect 212380 8206 212382 8258
rect 212382 8206 212434 8258
rect 212434 8206 212436 8258
rect 212380 8204 212436 8206
rect 219516 55690 219572 55692
rect 219516 55638 219518 55690
rect 219518 55638 219570 55690
rect 219570 55638 219572 55690
rect 219516 55636 219572 55638
rect 219620 55690 219676 55692
rect 219620 55638 219622 55690
rect 219622 55638 219674 55690
rect 219674 55638 219676 55690
rect 219620 55636 219676 55638
rect 219724 55690 219780 55692
rect 219724 55638 219726 55690
rect 219726 55638 219778 55690
rect 219778 55638 219780 55690
rect 219724 55636 219780 55638
rect 220668 54572 220724 54628
rect 219516 54122 219572 54124
rect 219516 54070 219518 54122
rect 219518 54070 219570 54122
rect 219570 54070 219572 54122
rect 219516 54068 219572 54070
rect 219620 54122 219676 54124
rect 219620 54070 219622 54122
rect 219622 54070 219674 54122
rect 219674 54070 219676 54122
rect 219620 54068 219676 54070
rect 219724 54122 219780 54124
rect 219724 54070 219726 54122
rect 219726 54070 219778 54122
rect 219778 54070 219780 54122
rect 219724 54068 219780 54070
rect 219516 52554 219572 52556
rect 219516 52502 219518 52554
rect 219518 52502 219570 52554
rect 219570 52502 219572 52554
rect 219516 52500 219572 52502
rect 219620 52554 219676 52556
rect 219620 52502 219622 52554
rect 219622 52502 219674 52554
rect 219674 52502 219676 52554
rect 219620 52500 219676 52502
rect 219724 52554 219780 52556
rect 219724 52502 219726 52554
rect 219726 52502 219778 52554
rect 219778 52502 219780 52554
rect 219724 52500 219780 52502
rect 219516 50986 219572 50988
rect 219516 50934 219518 50986
rect 219518 50934 219570 50986
rect 219570 50934 219572 50986
rect 219516 50932 219572 50934
rect 219620 50986 219676 50988
rect 219620 50934 219622 50986
rect 219622 50934 219674 50986
rect 219674 50934 219676 50986
rect 219620 50932 219676 50934
rect 219724 50986 219780 50988
rect 219724 50934 219726 50986
rect 219726 50934 219778 50986
rect 219778 50934 219780 50986
rect 219724 50932 219780 50934
rect 219516 49418 219572 49420
rect 219516 49366 219518 49418
rect 219518 49366 219570 49418
rect 219570 49366 219572 49418
rect 219516 49364 219572 49366
rect 219620 49418 219676 49420
rect 219620 49366 219622 49418
rect 219622 49366 219674 49418
rect 219674 49366 219676 49418
rect 219620 49364 219676 49366
rect 219724 49418 219780 49420
rect 219724 49366 219726 49418
rect 219726 49366 219778 49418
rect 219778 49366 219780 49418
rect 219724 49364 219780 49366
rect 219516 47850 219572 47852
rect 219516 47798 219518 47850
rect 219518 47798 219570 47850
rect 219570 47798 219572 47850
rect 219516 47796 219572 47798
rect 219620 47850 219676 47852
rect 219620 47798 219622 47850
rect 219622 47798 219674 47850
rect 219674 47798 219676 47850
rect 219620 47796 219676 47798
rect 219724 47850 219780 47852
rect 219724 47798 219726 47850
rect 219726 47798 219778 47850
rect 219778 47798 219780 47850
rect 219724 47796 219780 47798
rect 219516 46282 219572 46284
rect 219516 46230 219518 46282
rect 219518 46230 219570 46282
rect 219570 46230 219572 46282
rect 219516 46228 219572 46230
rect 219620 46282 219676 46284
rect 219620 46230 219622 46282
rect 219622 46230 219674 46282
rect 219674 46230 219676 46282
rect 219620 46228 219676 46230
rect 219724 46282 219780 46284
rect 219724 46230 219726 46282
rect 219726 46230 219778 46282
rect 219778 46230 219780 46282
rect 219724 46228 219780 46230
rect 219516 44714 219572 44716
rect 219516 44662 219518 44714
rect 219518 44662 219570 44714
rect 219570 44662 219572 44714
rect 219516 44660 219572 44662
rect 219620 44714 219676 44716
rect 219620 44662 219622 44714
rect 219622 44662 219674 44714
rect 219674 44662 219676 44714
rect 219620 44660 219676 44662
rect 219724 44714 219780 44716
rect 219724 44662 219726 44714
rect 219726 44662 219778 44714
rect 219778 44662 219780 44714
rect 219724 44660 219780 44662
rect 219516 43146 219572 43148
rect 219516 43094 219518 43146
rect 219518 43094 219570 43146
rect 219570 43094 219572 43146
rect 219516 43092 219572 43094
rect 219620 43146 219676 43148
rect 219620 43094 219622 43146
rect 219622 43094 219674 43146
rect 219674 43094 219676 43146
rect 219620 43092 219676 43094
rect 219724 43146 219780 43148
rect 219724 43094 219726 43146
rect 219726 43094 219778 43146
rect 219778 43094 219780 43146
rect 219724 43092 219780 43094
rect 219516 41578 219572 41580
rect 219516 41526 219518 41578
rect 219518 41526 219570 41578
rect 219570 41526 219572 41578
rect 219516 41524 219572 41526
rect 219620 41578 219676 41580
rect 219620 41526 219622 41578
rect 219622 41526 219674 41578
rect 219674 41526 219676 41578
rect 219620 41524 219676 41526
rect 219724 41578 219780 41580
rect 219724 41526 219726 41578
rect 219726 41526 219778 41578
rect 219778 41526 219780 41578
rect 219724 41524 219780 41526
rect 219516 40010 219572 40012
rect 219516 39958 219518 40010
rect 219518 39958 219570 40010
rect 219570 39958 219572 40010
rect 219516 39956 219572 39958
rect 219620 40010 219676 40012
rect 219620 39958 219622 40010
rect 219622 39958 219674 40010
rect 219674 39958 219676 40010
rect 219620 39956 219676 39958
rect 219724 40010 219780 40012
rect 219724 39958 219726 40010
rect 219726 39958 219778 40010
rect 219778 39958 219780 40010
rect 219724 39956 219780 39958
rect 219516 38442 219572 38444
rect 219516 38390 219518 38442
rect 219518 38390 219570 38442
rect 219570 38390 219572 38442
rect 219516 38388 219572 38390
rect 219620 38442 219676 38444
rect 219620 38390 219622 38442
rect 219622 38390 219674 38442
rect 219674 38390 219676 38442
rect 219620 38388 219676 38390
rect 219724 38442 219780 38444
rect 219724 38390 219726 38442
rect 219726 38390 219778 38442
rect 219778 38390 219780 38442
rect 219724 38388 219780 38390
rect 219516 36874 219572 36876
rect 219516 36822 219518 36874
rect 219518 36822 219570 36874
rect 219570 36822 219572 36874
rect 219516 36820 219572 36822
rect 219620 36874 219676 36876
rect 219620 36822 219622 36874
rect 219622 36822 219674 36874
rect 219674 36822 219676 36874
rect 219620 36820 219676 36822
rect 219724 36874 219780 36876
rect 219724 36822 219726 36874
rect 219726 36822 219778 36874
rect 219778 36822 219780 36874
rect 219724 36820 219780 36822
rect 219516 35306 219572 35308
rect 219516 35254 219518 35306
rect 219518 35254 219570 35306
rect 219570 35254 219572 35306
rect 219516 35252 219572 35254
rect 219620 35306 219676 35308
rect 219620 35254 219622 35306
rect 219622 35254 219674 35306
rect 219674 35254 219676 35306
rect 219620 35252 219676 35254
rect 219724 35306 219780 35308
rect 219724 35254 219726 35306
rect 219726 35254 219778 35306
rect 219778 35254 219780 35306
rect 219724 35252 219780 35254
rect 219516 33738 219572 33740
rect 219516 33686 219518 33738
rect 219518 33686 219570 33738
rect 219570 33686 219572 33738
rect 219516 33684 219572 33686
rect 219620 33738 219676 33740
rect 219620 33686 219622 33738
rect 219622 33686 219674 33738
rect 219674 33686 219676 33738
rect 219620 33684 219676 33686
rect 219724 33738 219780 33740
rect 219724 33686 219726 33738
rect 219726 33686 219778 33738
rect 219778 33686 219780 33738
rect 219724 33684 219780 33686
rect 219516 32170 219572 32172
rect 219516 32118 219518 32170
rect 219518 32118 219570 32170
rect 219570 32118 219572 32170
rect 219516 32116 219572 32118
rect 219620 32170 219676 32172
rect 219620 32118 219622 32170
rect 219622 32118 219674 32170
rect 219674 32118 219676 32170
rect 219620 32116 219676 32118
rect 219724 32170 219780 32172
rect 219724 32118 219726 32170
rect 219726 32118 219778 32170
rect 219778 32118 219780 32170
rect 219724 32116 219780 32118
rect 219516 30602 219572 30604
rect 219516 30550 219518 30602
rect 219518 30550 219570 30602
rect 219570 30550 219572 30602
rect 219516 30548 219572 30550
rect 219620 30602 219676 30604
rect 219620 30550 219622 30602
rect 219622 30550 219674 30602
rect 219674 30550 219676 30602
rect 219620 30548 219676 30550
rect 219724 30602 219780 30604
rect 219724 30550 219726 30602
rect 219726 30550 219778 30602
rect 219778 30550 219780 30602
rect 219724 30548 219780 30550
rect 219516 29034 219572 29036
rect 219516 28982 219518 29034
rect 219518 28982 219570 29034
rect 219570 28982 219572 29034
rect 219516 28980 219572 28982
rect 219620 29034 219676 29036
rect 219620 28982 219622 29034
rect 219622 28982 219674 29034
rect 219674 28982 219676 29034
rect 219620 28980 219676 28982
rect 219724 29034 219780 29036
rect 219724 28982 219726 29034
rect 219726 28982 219778 29034
rect 219778 28982 219780 29034
rect 219724 28980 219780 28982
rect 219516 27466 219572 27468
rect 219516 27414 219518 27466
rect 219518 27414 219570 27466
rect 219570 27414 219572 27466
rect 219516 27412 219572 27414
rect 219620 27466 219676 27468
rect 219620 27414 219622 27466
rect 219622 27414 219674 27466
rect 219674 27414 219676 27466
rect 219620 27412 219676 27414
rect 219724 27466 219780 27468
rect 219724 27414 219726 27466
rect 219726 27414 219778 27466
rect 219778 27414 219780 27466
rect 219724 27412 219780 27414
rect 219516 25898 219572 25900
rect 219516 25846 219518 25898
rect 219518 25846 219570 25898
rect 219570 25846 219572 25898
rect 219516 25844 219572 25846
rect 219620 25898 219676 25900
rect 219620 25846 219622 25898
rect 219622 25846 219674 25898
rect 219674 25846 219676 25898
rect 219620 25844 219676 25846
rect 219724 25898 219780 25900
rect 219724 25846 219726 25898
rect 219726 25846 219778 25898
rect 219778 25846 219780 25898
rect 219724 25844 219780 25846
rect 219516 24330 219572 24332
rect 219516 24278 219518 24330
rect 219518 24278 219570 24330
rect 219570 24278 219572 24330
rect 219516 24276 219572 24278
rect 219620 24330 219676 24332
rect 219620 24278 219622 24330
rect 219622 24278 219674 24330
rect 219674 24278 219676 24330
rect 219620 24276 219676 24278
rect 219724 24330 219780 24332
rect 219724 24278 219726 24330
rect 219726 24278 219778 24330
rect 219778 24278 219780 24330
rect 219724 24276 219780 24278
rect 219516 22762 219572 22764
rect 219516 22710 219518 22762
rect 219518 22710 219570 22762
rect 219570 22710 219572 22762
rect 219516 22708 219572 22710
rect 219620 22762 219676 22764
rect 219620 22710 219622 22762
rect 219622 22710 219674 22762
rect 219674 22710 219676 22762
rect 219620 22708 219676 22710
rect 219724 22762 219780 22764
rect 219724 22710 219726 22762
rect 219726 22710 219778 22762
rect 219778 22710 219780 22762
rect 219724 22708 219780 22710
rect 219516 21194 219572 21196
rect 219516 21142 219518 21194
rect 219518 21142 219570 21194
rect 219570 21142 219572 21194
rect 219516 21140 219572 21142
rect 219620 21194 219676 21196
rect 219620 21142 219622 21194
rect 219622 21142 219674 21194
rect 219674 21142 219676 21194
rect 219620 21140 219676 21142
rect 219724 21194 219780 21196
rect 219724 21142 219726 21194
rect 219726 21142 219778 21194
rect 219778 21142 219780 21194
rect 219724 21140 219780 21142
rect 219516 19626 219572 19628
rect 219516 19574 219518 19626
rect 219518 19574 219570 19626
rect 219570 19574 219572 19626
rect 219516 19572 219572 19574
rect 219620 19626 219676 19628
rect 219620 19574 219622 19626
rect 219622 19574 219674 19626
rect 219674 19574 219676 19626
rect 219620 19572 219676 19574
rect 219724 19626 219780 19628
rect 219724 19574 219726 19626
rect 219726 19574 219778 19626
rect 219778 19574 219780 19626
rect 219724 19572 219780 19574
rect 219516 18058 219572 18060
rect 219516 18006 219518 18058
rect 219518 18006 219570 18058
rect 219570 18006 219572 18058
rect 219516 18004 219572 18006
rect 219620 18058 219676 18060
rect 219620 18006 219622 18058
rect 219622 18006 219674 18058
rect 219674 18006 219676 18058
rect 219620 18004 219676 18006
rect 219724 18058 219780 18060
rect 219724 18006 219726 18058
rect 219726 18006 219778 18058
rect 219778 18006 219780 18058
rect 219724 18004 219780 18006
rect 219516 16490 219572 16492
rect 219516 16438 219518 16490
rect 219518 16438 219570 16490
rect 219570 16438 219572 16490
rect 219516 16436 219572 16438
rect 219620 16490 219676 16492
rect 219620 16438 219622 16490
rect 219622 16438 219674 16490
rect 219674 16438 219676 16490
rect 219620 16436 219676 16438
rect 219724 16490 219780 16492
rect 219724 16438 219726 16490
rect 219726 16438 219778 16490
rect 219778 16438 219780 16490
rect 219724 16436 219780 16438
rect 219516 14922 219572 14924
rect 219516 14870 219518 14922
rect 219518 14870 219570 14922
rect 219570 14870 219572 14922
rect 219516 14868 219572 14870
rect 219620 14922 219676 14924
rect 219620 14870 219622 14922
rect 219622 14870 219674 14922
rect 219674 14870 219676 14922
rect 219620 14868 219676 14870
rect 219724 14922 219780 14924
rect 219724 14870 219726 14922
rect 219726 14870 219778 14922
rect 219778 14870 219780 14922
rect 219724 14868 219780 14870
rect 219516 13354 219572 13356
rect 219516 13302 219518 13354
rect 219518 13302 219570 13354
rect 219570 13302 219572 13354
rect 219516 13300 219572 13302
rect 219620 13354 219676 13356
rect 219620 13302 219622 13354
rect 219622 13302 219674 13354
rect 219674 13302 219676 13354
rect 219620 13300 219676 13302
rect 219724 13354 219780 13356
rect 219724 13302 219726 13354
rect 219726 13302 219778 13354
rect 219778 13302 219780 13354
rect 219724 13300 219780 13302
rect 217308 11788 217364 11844
rect 217420 12908 217476 12964
rect 213612 10332 213668 10388
rect 213388 9100 213444 9156
rect 219516 11786 219572 11788
rect 219516 11734 219518 11786
rect 219518 11734 219570 11786
rect 219570 11734 219572 11786
rect 219516 11732 219572 11734
rect 219620 11786 219676 11788
rect 219620 11734 219622 11786
rect 219622 11734 219674 11786
rect 219674 11734 219676 11786
rect 219620 11732 219676 11734
rect 219724 11786 219780 11788
rect 219724 11734 219726 11786
rect 219726 11734 219778 11786
rect 219778 11734 219780 11786
rect 219724 11732 219780 11734
rect 219516 10218 219572 10220
rect 219516 10166 219518 10218
rect 219518 10166 219570 10218
rect 219570 10166 219572 10218
rect 219516 10164 219572 10166
rect 219620 10218 219676 10220
rect 219620 10166 219622 10218
rect 219622 10166 219674 10218
rect 219674 10166 219676 10218
rect 219620 10164 219676 10166
rect 219724 10218 219780 10220
rect 219724 10166 219726 10218
rect 219726 10166 219778 10218
rect 219778 10166 219780 10218
rect 219724 10164 219780 10166
rect 216748 9548 216804 9604
rect 220556 9996 220612 10052
rect 218316 9772 218372 9828
rect 217532 9548 217588 9604
rect 213836 9042 213892 9044
rect 213836 8990 213838 9042
rect 213838 8990 213890 9042
rect 213890 8990 213892 9042
rect 213836 8988 213892 8990
rect 216524 9042 216580 9044
rect 216524 8990 216526 9042
rect 216526 8990 216578 9042
rect 216578 8990 216580 9042
rect 216524 8988 216580 8990
rect 215740 8540 215796 8596
rect 213388 8258 213444 8260
rect 213388 8206 213390 8258
rect 213390 8206 213442 8258
rect 213442 8206 213444 8258
rect 213388 8204 213444 8206
rect 212828 8146 212884 8148
rect 212828 8094 212830 8146
rect 212830 8094 212882 8146
rect 212882 8094 212884 8146
rect 212828 8092 212884 8094
rect 212716 7980 212772 8036
rect 214060 7532 214116 7588
rect 214732 7532 214788 7588
rect 214508 7308 214564 7364
rect 213836 6860 213892 6916
rect 214620 6860 214676 6916
rect 213612 6466 213668 6468
rect 213612 6414 213614 6466
rect 213614 6414 213666 6466
rect 213666 6414 213668 6466
rect 213612 6412 213668 6414
rect 211596 4396 211652 4452
rect 211372 3442 211428 3444
rect 211372 3390 211374 3442
rect 211374 3390 211426 3442
rect 211426 3390 211428 3442
rect 211372 3388 211428 3390
rect 212380 4508 212436 4564
rect 212492 4732 212548 4788
rect 211932 4396 211988 4452
rect 212044 3554 212100 3556
rect 212044 3502 212046 3554
rect 212046 3502 212098 3554
rect 212098 3502 212100 3554
rect 212044 3500 212100 3502
rect 216972 8316 217028 8372
rect 216972 7756 217028 7812
rect 217308 8428 217364 8484
rect 216412 7474 216468 7476
rect 216412 7422 216414 7474
rect 216414 7422 216466 7474
rect 216466 7422 216468 7474
rect 216412 7420 216468 7422
rect 214732 5180 214788 5236
rect 213612 4956 213668 5012
rect 214508 4620 214564 4676
rect 215292 5852 215348 5908
rect 215852 5794 215908 5796
rect 215852 5742 215854 5794
rect 215854 5742 215906 5794
rect 215906 5742 215908 5794
rect 215852 5740 215908 5742
rect 216412 5740 216468 5796
rect 216748 6972 216804 7028
rect 217196 7308 217252 7364
rect 217196 6748 217252 6804
rect 215964 5292 216020 5348
rect 215628 5180 215684 5236
rect 215180 4956 215236 5012
rect 215292 4620 215348 4676
rect 215404 4562 215460 4564
rect 215404 4510 215406 4562
rect 215406 4510 215458 4562
rect 215458 4510 215460 4562
rect 215404 4508 215460 4510
rect 216188 5122 216244 5124
rect 216188 5070 216190 5122
rect 216190 5070 216242 5122
rect 216242 5070 216244 5122
rect 216188 5068 216244 5070
rect 216076 5010 216132 5012
rect 216076 4958 216078 5010
rect 216078 4958 216130 5010
rect 216130 4958 216132 5010
rect 216076 4956 216132 4958
rect 216300 4898 216356 4900
rect 216300 4846 216302 4898
rect 216302 4846 216354 4898
rect 216354 4846 216356 4898
rect 216300 4844 216356 4846
rect 215964 4562 216020 4564
rect 215964 4510 215966 4562
rect 215966 4510 216018 4562
rect 216018 4510 216020 4562
rect 215964 4508 216020 4510
rect 217084 5794 217140 5796
rect 217084 5742 217086 5794
rect 217086 5742 217138 5794
rect 217138 5742 217140 5794
rect 217084 5740 217140 5742
rect 217756 9212 217812 9268
rect 217756 8146 217812 8148
rect 217756 8094 217758 8146
rect 217758 8094 217810 8146
rect 217810 8094 217812 8146
rect 217756 8092 217812 8094
rect 217756 7420 217812 7476
rect 217644 6466 217700 6468
rect 217644 6414 217646 6466
rect 217646 6414 217698 6466
rect 217698 6414 217700 6466
rect 217644 6412 217700 6414
rect 217868 6076 217924 6132
rect 216636 4956 216692 5012
rect 217756 5068 217812 5124
rect 216860 4844 216916 4900
rect 216748 4450 216804 4452
rect 216748 4398 216750 4450
rect 216750 4398 216802 4450
rect 216802 4398 216804 4450
rect 216748 4396 216804 4398
rect 216524 4338 216580 4340
rect 216524 4286 216526 4338
rect 216526 4286 216578 4338
rect 216578 4286 216580 4338
rect 216524 4284 216580 4286
rect 212828 3724 212884 3780
rect 212268 3500 212324 3556
rect 211820 2268 211876 2324
rect 212828 3442 212884 3444
rect 212828 3390 212830 3442
rect 212830 3390 212882 3442
rect 212882 3390 212884 3442
rect 212828 3388 212884 3390
rect 217084 4956 217140 5012
rect 217308 4562 217364 4564
rect 217308 4510 217310 4562
rect 217310 4510 217362 4562
rect 217362 4510 217364 4562
rect 217308 4508 217364 4510
rect 218204 8316 218260 8372
rect 218092 8092 218148 8148
rect 218204 6748 218260 6804
rect 218428 9660 218484 9716
rect 219548 9660 219604 9716
rect 219100 9266 219156 9268
rect 219100 9214 219102 9266
rect 219102 9214 219154 9266
rect 219154 9214 219156 9266
rect 219100 9212 219156 9214
rect 219996 9212 220052 9268
rect 218764 9042 218820 9044
rect 218764 8990 218766 9042
rect 218766 8990 218818 9042
rect 218818 8990 218820 9042
rect 218764 8988 218820 8990
rect 219516 8650 219572 8652
rect 219516 8598 219518 8650
rect 219518 8598 219570 8650
rect 219570 8598 219572 8650
rect 219516 8596 219572 8598
rect 219620 8650 219676 8652
rect 219620 8598 219622 8650
rect 219622 8598 219674 8650
rect 219674 8598 219676 8650
rect 219620 8596 219676 8598
rect 219724 8650 219780 8652
rect 219724 8598 219726 8650
rect 219726 8598 219778 8650
rect 219778 8598 219780 8650
rect 219724 8596 219780 8598
rect 220332 9100 220388 9156
rect 221788 11228 221844 11284
rect 225932 53900 225988 53956
rect 222684 10332 222740 10388
rect 224252 53788 224308 53844
rect 221788 9660 221844 9716
rect 221228 9212 221284 9268
rect 221900 9212 221956 9268
rect 222348 9266 222404 9268
rect 222348 9214 222350 9266
rect 222350 9214 222402 9266
rect 222402 9214 222404 9266
rect 222348 9212 222404 9214
rect 224252 9212 224308 9268
rect 220220 8092 220276 8148
rect 220220 7868 220276 7924
rect 220780 7756 220836 7812
rect 220668 7644 220724 7700
rect 219516 7082 219572 7084
rect 219516 7030 219518 7082
rect 219518 7030 219570 7082
rect 219570 7030 219572 7082
rect 219516 7028 219572 7030
rect 219620 7082 219676 7084
rect 219620 7030 219622 7082
rect 219622 7030 219674 7082
rect 219674 7030 219676 7082
rect 219620 7028 219676 7030
rect 219724 7082 219780 7084
rect 219724 7030 219726 7082
rect 219726 7030 219778 7082
rect 219778 7030 219780 7082
rect 219724 7028 219780 7030
rect 218540 5180 218596 5236
rect 218876 6412 218932 6468
rect 219100 6076 219156 6132
rect 218988 5122 219044 5124
rect 218988 5070 218990 5122
rect 218990 5070 219042 5122
rect 219042 5070 219044 5122
rect 218988 5068 219044 5070
rect 217532 4450 217588 4452
rect 217532 4398 217534 4450
rect 217534 4398 217586 4450
rect 217586 4398 217588 4450
rect 217532 4396 217588 4398
rect 217980 4338 218036 4340
rect 217980 4286 217982 4338
rect 217982 4286 218034 4338
rect 218034 4286 218036 4338
rect 217980 4284 218036 4286
rect 219516 5514 219572 5516
rect 219516 5462 219518 5514
rect 219518 5462 219570 5514
rect 219570 5462 219572 5514
rect 219516 5460 219572 5462
rect 219620 5514 219676 5516
rect 219620 5462 219622 5514
rect 219622 5462 219674 5514
rect 219674 5462 219676 5514
rect 219620 5460 219676 5462
rect 219724 5514 219780 5516
rect 219724 5462 219726 5514
rect 219726 5462 219778 5514
rect 219778 5462 219780 5514
rect 219724 5460 219780 5462
rect 221004 8146 221060 8148
rect 221004 8094 221006 8146
rect 221006 8094 221058 8146
rect 221058 8094 221060 8146
rect 221004 8092 221060 8094
rect 221228 7868 221284 7924
rect 219100 4172 219156 4228
rect 216860 3724 216916 3780
rect 210476 2156 210532 2212
rect 210364 1484 210420 1540
rect 216412 3330 216468 3332
rect 216412 3278 216414 3330
rect 216414 3278 216466 3330
rect 216466 3278 216468 3330
rect 216412 3276 216468 3278
rect 219548 4396 219604 4452
rect 219324 4226 219380 4228
rect 219324 4174 219326 4226
rect 219326 4174 219378 4226
rect 219378 4174 219380 4226
rect 219324 4172 219380 4174
rect 219548 4060 219604 4116
rect 219516 3946 219572 3948
rect 219516 3894 219518 3946
rect 219518 3894 219570 3946
rect 219570 3894 219572 3946
rect 219516 3892 219572 3894
rect 219620 3946 219676 3948
rect 219620 3894 219622 3946
rect 219622 3894 219674 3946
rect 219674 3894 219676 3946
rect 219620 3892 219676 3894
rect 219724 3946 219780 3948
rect 219724 3894 219726 3946
rect 219726 3894 219778 3946
rect 219778 3894 219780 3946
rect 219724 3892 219780 3894
rect 220108 4732 220164 4788
rect 220108 4172 220164 4228
rect 220668 4844 220724 4900
rect 220556 4732 220612 4788
rect 220332 4172 220388 4228
rect 219100 2716 219156 2772
rect 220220 3948 220276 4004
rect 220668 4450 220724 4452
rect 220668 4398 220670 4450
rect 220670 4398 220722 4450
rect 220722 4398 220724 4450
rect 220668 4396 220724 4398
rect 220780 4284 220836 4340
rect 221452 8316 221508 8372
rect 221564 8092 221620 8148
rect 221676 7868 221732 7924
rect 222012 8370 222068 8372
rect 222012 8318 222014 8370
rect 222014 8318 222066 8370
rect 222066 8318 222068 8370
rect 222012 8316 222068 8318
rect 234876 56474 234932 56476
rect 234876 56422 234878 56474
rect 234878 56422 234930 56474
rect 234930 56422 234932 56474
rect 234876 56420 234932 56422
rect 234980 56474 235036 56476
rect 234980 56422 234982 56474
rect 234982 56422 235034 56474
rect 235034 56422 235036 56474
rect 234980 56420 235036 56422
rect 235084 56474 235140 56476
rect 235084 56422 235086 56474
rect 235086 56422 235138 56474
rect 235138 56422 235140 56474
rect 235084 56420 235140 56422
rect 233548 56306 233604 56308
rect 233548 56254 233550 56306
rect 233550 56254 233602 56306
rect 233602 56254 233604 56306
rect 233548 56252 233604 56254
rect 234220 56252 234276 56308
rect 265596 56474 265652 56476
rect 265596 56422 265598 56474
rect 265598 56422 265650 56474
rect 265650 56422 265652 56474
rect 265596 56420 265652 56422
rect 265700 56474 265756 56476
rect 265700 56422 265702 56474
rect 265702 56422 265754 56474
rect 265754 56422 265756 56474
rect 265700 56420 265756 56422
rect 265804 56474 265860 56476
rect 265804 56422 265806 56474
rect 265806 56422 265858 56474
rect 265858 56422 265860 56474
rect 265804 56420 265860 56422
rect 260092 56028 260148 56084
rect 260764 56082 260820 56084
rect 260764 56030 260766 56082
rect 260766 56030 260818 56082
rect 260818 56030 260820 56082
rect 260764 56028 260820 56030
rect 271516 56028 271572 56084
rect 272188 56082 272244 56084
rect 272188 56030 272190 56082
rect 272190 56030 272242 56082
rect 272242 56030 272244 56082
rect 272188 56028 272244 56030
rect 296316 56474 296372 56476
rect 296316 56422 296318 56474
rect 296318 56422 296370 56474
rect 296370 56422 296372 56474
rect 296316 56420 296372 56422
rect 296420 56474 296476 56476
rect 296420 56422 296422 56474
rect 296422 56422 296474 56474
rect 296474 56422 296476 56474
rect 296420 56420 296476 56422
rect 296524 56474 296580 56476
rect 296524 56422 296526 56474
rect 296526 56422 296578 56474
rect 296578 56422 296580 56474
rect 296524 56420 296580 56422
rect 281596 56028 281652 56084
rect 282716 56082 282772 56084
rect 282716 56030 282718 56082
rect 282718 56030 282770 56082
rect 282770 56030 282772 56082
rect 282716 56028 282772 56030
rect 283612 56082 283668 56084
rect 283612 56030 283614 56082
rect 283614 56030 283666 56082
rect 283666 56030 283668 56082
rect 283612 56028 283668 56030
rect 234876 54906 234932 54908
rect 234876 54854 234878 54906
rect 234878 54854 234930 54906
rect 234930 54854 234932 54906
rect 234876 54852 234932 54854
rect 234980 54906 235036 54908
rect 234980 54854 234982 54906
rect 234982 54854 235034 54906
rect 235034 54854 235036 54906
rect 234980 54852 235036 54854
rect 235084 54906 235140 54908
rect 235084 54854 235086 54906
rect 235086 54854 235138 54906
rect 235138 54854 235140 54906
rect 235084 54852 235140 54854
rect 239260 54572 239316 54628
rect 233996 53900 234052 53956
rect 228060 53788 228116 53844
rect 234876 53338 234932 53340
rect 234876 53286 234878 53338
rect 234878 53286 234930 53338
rect 234930 53286 234932 53338
rect 234876 53284 234932 53286
rect 234980 53338 235036 53340
rect 234980 53286 234982 53338
rect 234982 53286 235034 53338
rect 235034 53286 235036 53338
rect 234980 53284 235036 53286
rect 235084 53338 235140 53340
rect 235084 53286 235086 53338
rect 235086 53286 235138 53338
rect 235138 53286 235140 53338
rect 235084 53284 235140 53286
rect 234876 51770 234932 51772
rect 234876 51718 234878 51770
rect 234878 51718 234930 51770
rect 234930 51718 234932 51770
rect 234876 51716 234932 51718
rect 234980 51770 235036 51772
rect 234980 51718 234982 51770
rect 234982 51718 235034 51770
rect 235034 51718 235036 51770
rect 234980 51716 235036 51718
rect 235084 51770 235140 51772
rect 235084 51718 235086 51770
rect 235086 51718 235138 51770
rect 235138 51718 235140 51770
rect 235084 51716 235140 51718
rect 234876 50202 234932 50204
rect 234876 50150 234878 50202
rect 234878 50150 234930 50202
rect 234930 50150 234932 50202
rect 234876 50148 234932 50150
rect 234980 50202 235036 50204
rect 234980 50150 234982 50202
rect 234982 50150 235034 50202
rect 235034 50150 235036 50202
rect 234980 50148 235036 50150
rect 235084 50202 235140 50204
rect 235084 50150 235086 50202
rect 235086 50150 235138 50202
rect 235138 50150 235140 50202
rect 235084 50148 235140 50150
rect 234876 48634 234932 48636
rect 234876 48582 234878 48634
rect 234878 48582 234930 48634
rect 234930 48582 234932 48634
rect 234876 48580 234932 48582
rect 234980 48634 235036 48636
rect 234980 48582 234982 48634
rect 234982 48582 235034 48634
rect 235034 48582 235036 48634
rect 234980 48580 235036 48582
rect 235084 48634 235140 48636
rect 235084 48582 235086 48634
rect 235086 48582 235138 48634
rect 235138 48582 235140 48634
rect 235084 48580 235140 48582
rect 234876 47066 234932 47068
rect 234876 47014 234878 47066
rect 234878 47014 234930 47066
rect 234930 47014 234932 47066
rect 234876 47012 234932 47014
rect 234980 47066 235036 47068
rect 234980 47014 234982 47066
rect 234982 47014 235034 47066
rect 235034 47014 235036 47066
rect 234980 47012 235036 47014
rect 235084 47066 235140 47068
rect 235084 47014 235086 47066
rect 235086 47014 235138 47066
rect 235138 47014 235140 47066
rect 235084 47012 235140 47014
rect 234876 45498 234932 45500
rect 234876 45446 234878 45498
rect 234878 45446 234930 45498
rect 234930 45446 234932 45498
rect 234876 45444 234932 45446
rect 234980 45498 235036 45500
rect 234980 45446 234982 45498
rect 234982 45446 235034 45498
rect 235034 45446 235036 45498
rect 234980 45444 235036 45446
rect 235084 45498 235140 45500
rect 235084 45446 235086 45498
rect 235086 45446 235138 45498
rect 235138 45446 235140 45498
rect 235084 45444 235140 45446
rect 234876 43930 234932 43932
rect 234876 43878 234878 43930
rect 234878 43878 234930 43930
rect 234930 43878 234932 43930
rect 234876 43876 234932 43878
rect 234980 43930 235036 43932
rect 234980 43878 234982 43930
rect 234982 43878 235034 43930
rect 235034 43878 235036 43930
rect 234980 43876 235036 43878
rect 235084 43930 235140 43932
rect 235084 43878 235086 43930
rect 235086 43878 235138 43930
rect 235138 43878 235140 43930
rect 235084 43876 235140 43878
rect 234876 42362 234932 42364
rect 234876 42310 234878 42362
rect 234878 42310 234930 42362
rect 234930 42310 234932 42362
rect 234876 42308 234932 42310
rect 234980 42362 235036 42364
rect 234980 42310 234982 42362
rect 234982 42310 235034 42362
rect 235034 42310 235036 42362
rect 234980 42308 235036 42310
rect 235084 42362 235140 42364
rect 235084 42310 235086 42362
rect 235086 42310 235138 42362
rect 235138 42310 235140 42362
rect 235084 42308 235140 42310
rect 234876 40794 234932 40796
rect 234876 40742 234878 40794
rect 234878 40742 234930 40794
rect 234930 40742 234932 40794
rect 234876 40740 234932 40742
rect 234980 40794 235036 40796
rect 234980 40742 234982 40794
rect 234982 40742 235034 40794
rect 235034 40742 235036 40794
rect 234980 40740 235036 40742
rect 235084 40794 235140 40796
rect 235084 40742 235086 40794
rect 235086 40742 235138 40794
rect 235138 40742 235140 40794
rect 235084 40740 235140 40742
rect 234876 39226 234932 39228
rect 234876 39174 234878 39226
rect 234878 39174 234930 39226
rect 234930 39174 234932 39226
rect 234876 39172 234932 39174
rect 234980 39226 235036 39228
rect 234980 39174 234982 39226
rect 234982 39174 235034 39226
rect 235034 39174 235036 39226
rect 234980 39172 235036 39174
rect 235084 39226 235140 39228
rect 235084 39174 235086 39226
rect 235086 39174 235138 39226
rect 235138 39174 235140 39226
rect 235084 39172 235140 39174
rect 234876 37658 234932 37660
rect 234876 37606 234878 37658
rect 234878 37606 234930 37658
rect 234930 37606 234932 37658
rect 234876 37604 234932 37606
rect 234980 37658 235036 37660
rect 234980 37606 234982 37658
rect 234982 37606 235034 37658
rect 235034 37606 235036 37658
rect 234980 37604 235036 37606
rect 235084 37658 235140 37660
rect 235084 37606 235086 37658
rect 235086 37606 235138 37658
rect 235138 37606 235140 37658
rect 235084 37604 235140 37606
rect 234876 36090 234932 36092
rect 234876 36038 234878 36090
rect 234878 36038 234930 36090
rect 234930 36038 234932 36090
rect 234876 36036 234932 36038
rect 234980 36090 235036 36092
rect 234980 36038 234982 36090
rect 234982 36038 235034 36090
rect 235034 36038 235036 36090
rect 234980 36036 235036 36038
rect 235084 36090 235140 36092
rect 235084 36038 235086 36090
rect 235086 36038 235138 36090
rect 235138 36038 235140 36090
rect 235084 36036 235140 36038
rect 234876 34522 234932 34524
rect 234876 34470 234878 34522
rect 234878 34470 234930 34522
rect 234930 34470 234932 34522
rect 234876 34468 234932 34470
rect 234980 34522 235036 34524
rect 234980 34470 234982 34522
rect 234982 34470 235034 34522
rect 235034 34470 235036 34522
rect 234980 34468 235036 34470
rect 235084 34522 235140 34524
rect 235084 34470 235086 34522
rect 235086 34470 235138 34522
rect 235138 34470 235140 34522
rect 235084 34468 235140 34470
rect 234876 32954 234932 32956
rect 234876 32902 234878 32954
rect 234878 32902 234930 32954
rect 234930 32902 234932 32954
rect 234876 32900 234932 32902
rect 234980 32954 235036 32956
rect 234980 32902 234982 32954
rect 234982 32902 235034 32954
rect 235034 32902 235036 32954
rect 234980 32900 235036 32902
rect 235084 32954 235140 32956
rect 235084 32902 235086 32954
rect 235086 32902 235138 32954
rect 235138 32902 235140 32954
rect 235084 32900 235140 32902
rect 234876 31386 234932 31388
rect 234876 31334 234878 31386
rect 234878 31334 234930 31386
rect 234930 31334 234932 31386
rect 234876 31332 234932 31334
rect 234980 31386 235036 31388
rect 234980 31334 234982 31386
rect 234982 31334 235034 31386
rect 235034 31334 235036 31386
rect 234980 31332 235036 31334
rect 235084 31386 235140 31388
rect 235084 31334 235086 31386
rect 235086 31334 235138 31386
rect 235138 31334 235140 31386
rect 235084 31332 235140 31334
rect 234876 29818 234932 29820
rect 234876 29766 234878 29818
rect 234878 29766 234930 29818
rect 234930 29766 234932 29818
rect 234876 29764 234932 29766
rect 234980 29818 235036 29820
rect 234980 29766 234982 29818
rect 234982 29766 235034 29818
rect 235034 29766 235036 29818
rect 234980 29764 235036 29766
rect 235084 29818 235140 29820
rect 235084 29766 235086 29818
rect 235086 29766 235138 29818
rect 235138 29766 235140 29818
rect 235084 29764 235140 29766
rect 234876 28250 234932 28252
rect 234876 28198 234878 28250
rect 234878 28198 234930 28250
rect 234930 28198 234932 28250
rect 234876 28196 234932 28198
rect 234980 28250 235036 28252
rect 234980 28198 234982 28250
rect 234982 28198 235034 28250
rect 235034 28198 235036 28250
rect 234980 28196 235036 28198
rect 235084 28250 235140 28252
rect 235084 28198 235086 28250
rect 235086 28198 235138 28250
rect 235138 28198 235140 28250
rect 235084 28196 235140 28198
rect 234876 26682 234932 26684
rect 234876 26630 234878 26682
rect 234878 26630 234930 26682
rect 234930 26630 234932 26682
rect 234876 26628 234932 26630
rect 234980 26682 235036 26684
rect 234980 26630 234982 26682
rect 234982 26630 235034 26682
rect 235034 26630 235036 26682
rect 234980 26628 235036 26630
rect 235084 26682 235140 26684
rect 235084 26630 235086 26682
rect 235086 26630 235138 26682
rect 235138 26630 235140 26682
rect 235084 26628 235140 26630
rect 234876 25114 234932 25116
rect 234876 25062 234878 25114
rect 234878 25062 234930 25114
rect 234930 25062 234932 25114
rect 234876 25060 234932 25062
rect 234980 25114 235036 25116
rect 234980 25062 234982 25114
rect 234982 25062 235034 25114
rect 235034 25062 235036 25114
rect 234980 25060 235036 25062
rect 235084 25114 235140 25116
rect 235084 25062 235086 25114
rect 235086 25062 235138 25114
rect 235138 25062 235140 25114
rect 235084 25060 235140 25062
rect 234876 23546 234932 23548
rect 234876 23494 234878 23546
rect 234878 23494 234930 23546
rect 234930 23494 234932 23546
rect 234876 23492 234932 23494
rect 234980 23546 235036 23548
rect 234980 23494 234982 23546
rect 234982 23494 235034 23546
rect 235034 23494 235036 23546
rect 234980 23492 235036 23494
rect 235084 23546 235140 23548
rect 235084 23494 235086 23546
rect 235086 23494 235138 23546
rect 235138 23494 235140 23546
rect 235084 23492 235140 23494
rect 234876 21978 234932 21980
rect 234876 21926 234878 21978
rect 234878 21926 234930 21978
rect 234930 21926 234932 21978
rect 234876 21924 234932 21926
rect 234980 21978 235036 21980
rect 234980 21926 234982 21978
rect 234982 21926 235034 21978
rect 235034 21926 235036 21978
rect 234980 21924 235036 21926
rect 235084 21978 235140 21980
rect 235084 21926 235086 21978
rect 235086 21926 235138 21978
rect 235138 21926 235140 21978
rect 235084 21924 235140 21926
rect 234876 20410 234932 20412
rect 234876 20358 234878 20410
rect 234878 20358 234930 20410
rect 234930 20358 234932 20410
rect 234876 20356 234932 20358
rect 234980 20410 235036 20412
rect 234980 20358 234982 20410
rect 234982 20358 235034 20410
rect 235034 20358 235036 20410
rect 234980 20356 235036 20358
rect 235084 20410 235140 20412
rect 235084 20358 235086 20410
rect 235086 20358 235138 20410
rect 235138 20358 235140 20410
rect 235084 20356 235140 20358
rect 234876 18842 234932 18844
rect 234876 18790 234878 18842
rect 234878 18790 234930 18842
rect 234930 18790 234932 18842
rect 234876 18788 234932 18790
rect 234980 18842 235036 18844
rect 234980 18790 234982 18842
rect 234982 18790 235034 18842
rect 235034 18790 235036 18842
rect 234980 18788 235036 18790
rect 235084 18842 235140 18844
rect 235084 18790 235086 18842
rect 235086 18790 235138 18842
rect 235138 18790 235140 18842
rect 235084 18788 235140 18790
rect 234876 17274 234932 17276
rect 234876 17222 234878 17274
rect 234878 17222 234930 17274
rect 234930 17222 234932 17274
rect 234876 17220 234932 17222
rect 234980 17274 235036 17276
rect 234980 17222 234982 17274
rect 234982 17222 235034 17274
rect 235034 17222 235036 17274
rect 234980 17220 235036 17222
rect 235084 17274 235140 17276
rect 235084 17222 235086 17274
rect 235086 17222 235138 17274
rect 235138 17222 235140 17274
rect 235084 17220 235140 17222
rect 234876 15706 234932 15708
rect 234876 15654 234878 15706
rect 234878 15654 234930 15706
rect 234930 15654 234932 15706
rect 234876 15652 234932 15654
rect 234980 15706 235036 15708
rect 234980 15654 234982 15706
rect 234982 15654 235034 15706
rect 235034 15654 235036 15706
rect 234980 15652 235036 15654
rect 235084 15706 235140 15708
rect 235084 15654 235086 15706
rect 235086 15654 235138 15706
rect 235138 15654 235140 15706
rect 235084 15652 235140 15654
rect 234876 14138 234932 14140
rect 234876 14086 234878 14138
rect 234878 14086 234930 14138
rect 234930 14086 234932 14138
rect 234876 14084 234932 14086
rect 234980 14138 235036 14140
rect 234980 14086 234982 14138
rect 234982 14086 235034 14138
rect 235034 14086 235036 14138
rect 234980 14084 235036 14086
rect 235084 14138 235140 14140
rect 235084 14086 235086 14138
rect 235086 14086 235138 14138
rect 235138 14086 235140 14138
rect 235084 14084 235140 14086
rect 234876 12570 234932 12572
rect 234876 12518 234878 12570
rect 234878 12518 234930 12570
rect 234930 12518 234932 12570
rect 234876 12516 234932 12518
rect 234980 12570 235036 12572
rect 234980 12518 234982 12570
rect 234982 12518 235034 12570
rect 235034 12518 235036 12570
rect 234980 12516 235036 12518
rect 235084 12570 235140 12572
rect 235084 12518 235086 12570
rect 235086 12518 235138 12570
rect 235138 12518 235140 12570
rect 235084 12516 235140 12518
rect 250236 55690 250292 55692
rect 250236 55638 250238 55690
rect 250238 55638 250290 55690
rect 250290 55638 250292 55690
rect 250236 55636 250292 55638
rect 250340 55690 250396 55692
rect 250340 55638 250342 55690
rect 250342 55638 250394 55690
rect 250394 55638 250396 55690
rect 250340 55636 250396 55638
rect 250444 55690 250500 55692
rect 250444 55638 250446 55690
rect 250446 55638 250498 55690
rect 250498 55638 250500 55690
rect 250444 55636 250500 55638
rect 250236 54122 250292 54124
rect 250236 54070 250238 54122
rect 250238 54070 250290 54122
rect 250290 54070 250292 54122
rect 250236 54068 250292 54070
rect 250340 54122 250396 54124
rect 250340 54070 250342 54122
rect 250342 54070 250394 54122
rect 250394 54070 250396 54122
rect 250340 54068 250396 54070
rect 250444 54122 250500 54124
rect 250444 54070 250446 54122
rect 250446 54070 250498 54122
rect 250498 54070 250500 54122
rect 250444 54068 250500 54070
rect 250236 52554 250292 52556
rect 250236 52502 250238 52554
rect 250238 52502 250290 52554
rect 250290 52502 250292 52554
rect 250236 52500 250292 52502
rect 250340 52554 250396 52556
rect 250340 52502 250342 52554
rect 250342 52502 250394 52554
rect 250394 52502 250396 52554
rect 250340 52500 250396 52502
rect 250444 52554 250500 52556
rect 250444 52502 250446 52554
rect 250446 52502 250498 52554
rect 250498 52502 250500 52554
rect 250444 52500 250500 52502
rect 250236 50986 250292 50988
rect 250236 50934 250238 50986
rect 250238 50934 250290 50986
rect 250290 50934 250292 50986
rect 250236 50932 250292 50934
rect 250340 50986 250396 50988
rect 250340 50934 250342 50986
rect 250342 50934 250394 50986
rect 250394 50934 250396 50986
rect 250340 50932 250396 50934
rect 250444 50986 250500 50988
rect 250444 50934 250446 50986
rect 250446 50934 250498 50986
rect 250498 50934 250500 50986
rect 250444 50932 250500 50934
rect 250236 49418 250292 49420
rect 250236 49366 250238 49418
rect 250238 49366 250290 49418
rect 250290 49366 250292 49418
rect 250236 49364 250292 49366
rect 250340 49418 250396 49420
rect 250340 49366 250342 49418
rect 250342 49366 250394 49418
rect 250394 49366 250396 49418
rect 250340 49364 250396 49366
rect 250444 49418 250500 49420
rect 250444 49366 250446 49418
rect 250446 49366 250498 49418
rect 250498 49366 250500 49418
rect 250444 49364 250500 49366
rect 250236 47850 250292 47852
rect 250236 47798 250238 47850
rect 250238 47798 250290 47850
rect 250290 47798 250292 47850
rect 250236 47796 250292 47798
rect 250340 47850 250396 47852
rect 250340 47798 250342 47850
rect 250342 47798 250394 47850
rect 250394 47798 250396 47850
rect 250340 47796 250396 47798
rect 250444 47850 250500 47852
rect 250444 47798 250446 47850
rect 250446 47798 250498 47850
rect 250498 47798 250500 47850
rect 250444 47796 250500 47798
rect 250236 46282 250292 46284
rect 250236 46230 250238 46282
rect 250238 46230 250290 46282
rect 250290 46230 250292 46282
rect 250236 46228 250292 46230
rect 250340 46282 250396 46284
rect 250340 46230 250342 46282
rect 250342 46230 250394 46282
rect 250394 46230 250396 46282
rect 250340 46228 250396 46230
rect 250444 46282 250500 46284
rect 250444 46230 250446 46282
rect 250446 46230 250498 46282
rect 250498 46230 250500 46282
rect 250444 46228 250500 46230
rect 250236 44714 250292 44716
rect 250236 44662 250238 44714
rect 250238 44662 250290 44714
rect 250290 44662 250292 44714
rect 250236 44660 250292 44662
rect 250340 44714 250396 44716
rect 250340 44662 250342 44714
rect 250342 44662 250394 44714
rect 250394 44662 250396 44714
rect 250340 44660 250396 44662
rect 250444 44714 250500 44716
rect 250444 44662 250446 44714
rect 250446 44662 250498 44714
rect 250498 44662 250500 44714
rect 250444 44660 250500 44662
rect 250236 43146 250292 43148
rect 250236 43094 250238 43146
rect 250238 43094 250290 43146
rect 250290 43094 250292 43146
rect 250236 43092 250292 43094
rect 250340 43146 250396 43148
rect 250340 43094 250342 43146
rect 250342 43094 250394 43146
rect 250394 43094 250396 43146
rect 250340 43092 250396 43094
rect 250444 43146 250500 43148
rect 250444 43094 250446 43146
rect 250446 43094 250498 43146
rect 250498 43094 250500 43146
rect 250444 43092 250500 43094
rect 250236 41578 250292 41580
rect 250236 41526 250238 41578
rect 250238 41526 250290 41578
rect 250290 41526 250292 41578
rect 250236 41524 250292 41526
rect 250340 41578 250396 41580
rect 250340 41526 250342 41578
rect 250342 41526 250394 41578
rect 250394 41526 250396 41578
rect 250340 41524 250396 41526
rect 250444 41578 250500 41580
rect 250444 41526 250446 41578
rect 250446 41526 250498 41578
rect 250498 41526 250500 41578
rect 250444 41524 250500 41526
rect 250236 40010 250292 40012
rect 250236 39958 250238 40010
rect 250238 39958 250290 40010
rect 250290 39958 250292 40010
rect 250236 39956 250292 39958
rect 250340 40010 250396 40012
rect 250340 39958 250342 40010
rect 250342 39958 250394 40010
rect 250394 39958 250396 40010
rect 250340 39956 250396 39958
rect 250444 40010 250500 40012
rect 250444 39958 250446 40010
rect 250446 39958 250498 40010
rect 250498 39958 250500 40010
rect 250444 39956 250500 39958
rect 250236 38442 250292 38444
rect 250236 38390 250238 38442
rect 250238 38390 250290 38442
rect 250290 38390 250292 38442
rect 250236 38388 250292 38390
rect 250340 38442 250396 38444
rect 250340 38390 250342 38442
rect 250342 38390 250394 38442
rect 250394 38390 250396 38442
rect 250340 38388 250396 38390
rect 250444 38442 250500 38444
rect 250444 38390 250446 38442
rect 250446 38390 250498 38442
rect 250498 38390 250500 38442
rect 250444 38388 250500 38390
rect 250236 36874 250292 36876
rect 250236 36822 250238 36874
rect 250238 36822 250290 36874
rect 250290 36822 250292 36874
rect 250236 36820 250292 36822
rect 250340 36874 250396 36876
rect 250340 36822 250342 36874
rect 250342 36822 250394 36874
rect 250394 36822 250396 36874
rect 250340 36820 250396 36822
rect 250444 36874 250500 36876
rect 250444 36822 250446 36874
rect 250446 36822 250498 36874
rect 250498 36822 250500 36874
rect 250444 36820 250500 36822
rect 250236 35306 250292 35308
rect 250236 35254 250238 35306
rect 250238 35254 250290 35306
rect 250290 35254 250292 35306
rect 250236 35252 250292 35254
rect 250340 35306 250396 35308
rect 250340 35254 250342 35306
rect 250342 35254 250394 35306
rect 250394 35254 250396 35306
rect 250340 35252 250396 35254
rect 250444 35306 250500 35308
rect 250444 35254 250446 35306
rect 250446 35254 250498 35306
rect 250498 35254 250500 35306
rect 250444 35252 250500 35254
rect 250236 33738 250292 33740
rect 250236 33686 250238 33738
rect 250238 33686 250290 33738
rect 250290 33686 250292 33738
rect 250236 33684 250292 33686
rect 250340 33738 250396 33740
rect 250340 33686 250342 33738
rect 250342 33686 250394 33738
rect 250394 33686 250396 33738
rect 250340 33684 250396 33686
rect 250444 33738 250500 33740
rect 250444 33686 250446 33738
rect 250446 33686 250498 33738
rect 250498 33686 250500 33738
rect 250444 33684 250500 33686
rect 250236 32170 250292 32172
rect 250236 32118 250238 32170
rect 250238 32118 250290 32170
rect 250290 32118 250292 32170
rect 250236 32116 250292 32118
rect 250340 32170 250396 32172
rect 250340 32118 250342 32170
rect 250342 32118 250394 32170
rect 250394 32118 250396 32170
rect 250340 32116 250396 32118
rect 250444 32170 250500 32172
rect 250444 32118 250446 32170
rect 250446 32118 250498 32170
rect 250498 32118 250500 32170
rect 250444 32116 250500 32118
rect 250236 30602 250292 30604
rect 250236 30550 250238 30602
rect 250238 30550 250290 30602
rect 250290 30550 250292 30602
rect 250236 30548 250292 30550
rect 250340 30602 250396 30604
rect 250340 30550 250342 30602
rect 250342 30550 250394 30602
rect 250394 30550 250396 30602
rect 250340 30548 250396 30550
rect 250444 30602 250500 30604
rect 250444 30550 250446 30602
rect 250446 30550 250498 30602
rect 250498 30550 250500 30602
rect 250444 30548 250500 30550
rect 250236 29034 250292 29036
rect 250236 28982 250238 29034
rect 250238 28982 250290 29034
rect 250290 28982 250292 29034
rect 250236 28980 250292 28982
rect 250340 29034 250396 29036
rect 250340 28982 250342 29034
rect 250342 28982 250394 29034
rect 250394 28982 250396 29034
rect 250340 28980 250396 28982
rect 250444 29034 250500 29036
rect 250444 28982 250446 29034
rect 250446 28982 250498 29034
rect 250498 28982 250500 29034
rect 250444 28980 250500 28982
rect 250236 27466 250292 27468
rect 250236 27414 250238 27466
rect 250238 27414 250290 27466
rect 250290 27414 250292 27466
rect 250236 27412 250292 27414
rect 250340 27466 250396 27468
rect 250340 27414 250342 27466
rect 250342 27414 250394 27466
rect 250394 27414 250396 27466
rect 250340 27412 250396 27414
rect 250444 27466 250500 27468
rect 250444 27414 250446 27466
rect 250446 27414 250498 27466
rect 250498 27414 250500 27466
rect 250444 27412 250500 27414
rect 250236 25898 250292 25900
rect 250236 25846 250238 25898
rect 250238 25846 250290 25898
rect 250290 25846 250292 25898
rect 250236 25844 250292 25846
rect 250340 25898 250396 25900
rect 250340 25846 250342 25898
rect 250342 25846 250394 25898
rect 250394 25846 250396 25898
rect 250340 25844 250396 25846
rect 250444 25898 250500 25900
rect 250444 25846 250446 25898
rect 250446 25846 250498 25898
rect 250498 25846 250500 25898
rect 250444 25844 250500 25846
rect 250236 24330 250292 24332
rect 250236 24278 250238 24330
rect 250238 24278 250290 24330
rect 250290 24278 250292 24330
rect 250236 24276 250292 24278
rect 250340 24330 250396 24332
rect 250340 24278 250342 24330
rect 250342 24278 250394 24330
rect 250394 24278 250396 24330
rect 250340 24276 250396 24278
rect 250444 24330 250500 24332
rect 250444 24278 250446 24330
rect 250446 24278 250498 24330
rect 250498 24278 250500 24330
rect 250444 24276 250500 24278
rect 250236 22762 250292 22764
rect 250236 22710 250238 22762
rect 250238 22710 250290 22762
rect 250290 22710 250292 22762
rect 250236 22708 250292 22710
rect 250340 22762 250396 22764
rect 250340 22710 250342 22762
rect 250342 22710 250394 22762
rect 250394 22710 250396 22762
rect 250340 22708 250396 22710
rect 250444 22762 250500 22764
rect 250444 22710 250446 22762
rect 250446 22710 250498 22762
rect 250498 22710 250500 22762
rect 250444 22708 250500 22710
rect 250236 21194 250292 21196
rect 250236 21142 250238 21194
rect 250238 21142 250290 21194
rect 250290 21142 250292 21194
rect 250236 21140 250292 21142
rect 250340 21194 250396 21196
rect 250340 21142 250342 21194
rect 250342 21142 250394 21194
rect 250394 21142 250396 21194
rect 250340 21140 250396 21142
rect 250444 21194 250500 21196
rect 250444 21142 250446 21194
rect 250446 21142 250498 21194
rect 250498 21142 250500 21194
rect 250444 21140 250500 21142
rect 250236 19626 250292 19628
rect 250236 19574 250238 19626
rect 250238 19574 250290 19626
rect 250290 19574 250292 19626
rect 250236 19572 250292 19574
rect 250340 19626 250396 19628
rect 250340 19574 250342 19626
rect 250342 19574 250394 19626
rect 250394 19574 250396 19626
rect 250340 19572 250396 19574
rect 250444 19626 250500 19628
rect 250444 19574 250446 19626
rect 250446 19574 250498 19626
rect 250498 19574 250500 19626
rect 250444 19572 250500 19574
rect 250236 18058 250292 18060
rect 250236 18006 250238 18058
rect 250238 18006 250290 18058
rect 250290 18006 250292 18058
rect 250236 18004 250292 18006
rect 250340 18058 250396 18060
rect 250340 18006 250342 18058
rect 250342 18006 250394 18058
rect 250394 18006 250396 18058
rect 250340 18004 250396 18006
rect 250444 18058 250500 18060
rect 250444 18006 250446 18058
rect 250446 18006 250498 18058
rect 250498 18006 250500 18058
rect 250444 18004 250500 18006
rect 250236 16490 250292 16492
rect 250236 16438 250238 16490
rect 250238 16438 250290 16490
rect 250290 16438 250292 16490
rect 250236 16436 250292 16438
rect 250340 16490 250396 16492
rect 250340 16438 250342 16490
rect 250342 16438 250394 16490
rect 250394 16438 250396 16490
rect 250340 16436 250396 16438
rect 250444 16490 250500 16492
rect 250444 16438 250446 16490
rect 250446 16438 250498 16490
rect 250498 16438 250500 16490
rect 250444 16436 250500 16438
rect 250236 14922 250292 14924
rect 250236 14870 250238 14922
rect 250238 14870 250290 14922
rect 250290 14870 250292 14922
rect 250236 14868 250292 14870
rect 250340 14922 250396 14924
rect 250340 14870 250342 14922
rect 250342 14870 250394 14922
rect 250394 14870 250396 14922
rect 250340 14868 250396 14870
rect 250444 14922 250500 14924
rect 250444 14870 250446 14922
rect 250446 14870 250498 14922
rect 250498 14870 250500 14922
rect 250444 14868 250500 14870
rect 256060 14252 256116 14308
rect 250236 13354 250292 13356
rect 250236 13302 250238 13354
rect 250238 13302 250290 13354
rect 250290 13302 250292 13354
rect 250236 13300 250292 13302
rect 250340 13354 250396 13356
rect 250340 13302 250342 13354
rect 250342 13302 250394 13354
rect 250394 13302 250396 13354
rect 250340 13300 250396 13302
rect 250444 13354 250500 13356
rect 250444 13302 250446 13354
rect 250446 13302 250498 13354
rect 250498 13302 250500 13354
rect 250444 13300 250500 13302
rect 250124 12908 250180 12964
rect 250236 11786 250292 11788
rect 250236 11734 250238 11786
rect 250238 11734 250290 11786
rect 250290 11734 250292 11786
rect 250236 11732 250292 11734
rect 250340 11786 250396 11788
rect 250340 11734 250342 11786
rect 250342 11734 250394 11786
rect 250394 11734 250396 11786
rect 250340 11732 250396 11734
rect 250444 11786 250500 11788
rect 250444 11734 250446 11786
rect 250446 11734 250498 11786
rect 250498 11734 250500 11786
rect 250444 11732 250500 11734
rect 244748 11228 244804 11284
rect 264572 55916 264628 55972
rect 266364 55970 266420 55972
rect 266364 55918 266366 55970
rect 266366 55918 266418 55970
rect 266418 55918 266420 55970
rect 266364 55916 266420 55918
rect 265596 54906 265652 54908
rect 265596 54854 265598 54906
rect 265598 54854 265650 54906
rect 265650 54854 265652 54906
rect 265596 54852 265652 54854
rect 265700 54906 265756 54908
rect 265700 54854 265702 54906
rect 265702 54854 265754 54906
rect 265754 54854 265756 54906
rect 265700 54852 265756 54854
rect 265804 54906 265860 54908
rect 265804 54854 265806 54906
rect 265806 54854 265858 54906
rect 265858 54854 265860 54906
rect 265804 54852 265860 54854
rect 265596 53338 265652 53340
rect 265596 53286 265598 53338
rect 265598 53286 265650 53338
rect 265650 53286 265652 53338
rect 265596 53284 265652 53286
rect 265700 53338 265756 53340
rect 265700 53286 265702 53338
rect 265702 53286 265754 53338
rect 265754 53286 265756 53338
rect 265700 53284 265756 53286
rect 265804 53338 265860 53340
rect 265804 53286 265806 53338
rect 265806 53286 265858 53338
rect 265858 53286 265860 53338
rect 265804 53284 265860 53286
rect 265596 51770 265652 51772
rect 265596 51718 265598 51770
rect 265598 51718 265650 51770
rect 265650 51718 265652 51770
rect 265596 51716 265652 51718
rect 265700 51770 265756 51772
rect 265700 51718 265702 51770
rect 265702 51718 265754 51770
rect 265754 51718 265756 51770
rect 265700 51716 265756 51718
rect 265804 51770 265860 51772
rect 265804 51718 265806 51770
rect 265806 51718 265858 51770
rect 265858 51718 265860 51770
rect 265804 51716 265860 51718
rect 265596 50202 265652 50204
rect 265596 50150 265598 50202
rect 265598 50150 265650 50202
rect 265650 50150 265652 50202
rect 265596 50148 265652 50150
rect 265700 50202 265756 50204
rect 265700 50150 265702 50202
rect 265702 50150 265754 50202
rect 265754 50150 265756 50202
rect 265700 50148 265756 50150
rect 265804 50202 265860 50204
rect 265804 50150 265806 50202
rect 265806 50150 265858 50202
rect 265858 50150 265860 50202
rect 265804 50148 265860 50150
rect 265596 48634 265652 48636
rect 265596 48582 265598 48634
rect 265598 48582 265650 48634
rect 265650 48582 265652 48634
rect 265596 48580 265652 48582
rect 265700 48634 265756 48636
rect 265700 48582 265702 48634
rect 265702 48582 265754 48634
rect 265754 48582 265756 48634
rect 265700 48580 265756 48582
rect 265804 48634 265860 48636
rect 265804 48582 265806 48634
rect 265806 48582 265858 48634
rect 265858 48582 265860 48634
rect 265804 48580 265860 48582
rect 265596 47066 265652 47068
rect 265596 47014 265598 47066
rect 265598 47014 265650 47066
rect 265650 47014 265652 47066
rect 265596 47012 265652 47014
rect 265700 47066 265756 47068
rect 265700 47014 265702 47066
rect 265702 47014 265754 47066
rect 265754 47014 265756 47066
rect 265700 47012 265756 47014
rect 265804 47066 265860 47068
rect 265804 47014 265806 47066
rect 265806 47014 265858 47066
rect 265858 47014 265860 47066
rect 265804 47012 265860 47014
rect 265596 45498 265652 45500
rect 265596 45446 265598 45498
rect 265598 45446 265650 45498
rect 265650 45446 265652 45498
rect 265596 45444 265652 45446
rect 265700 45498 265756 45500
rect 265700 45446 265702 45498
rect 265702 45446 265754 45498
rect 265754 45446 265756 45498
rect 265700 45444 265756 45446
rect 265804 45498 265860 45500
rect 265804 45446 265806 45498
rect 265806 45446 265858 45498
rect 265858 45446 265860 45498
rect 265804 45444 265860 45446
rect 265596 43930 265652 43932
rect 265596 43878 265598 43930
rect 265598 43878 265650 43930
rect 265650 43878 265652 43930
rect 265596 43876 265652 43878
rect 265700 43930 265756 43932
rect 265700 43878 265702 43930
rect 265702 43878 265754 43930
rect 265754 43878 265756 43930
rect 265700 43876 265756 43878
rect 265804 43930 265860 43932
rect 265804 43878 265806 43930
rect 265806 43878 265858 43930
rect 265858 43878 265860 43930
rect 265804 43876 265860 43878
rect 265596 42362 265652 42364
rect 265596 42310 265598 42362
rect 265598 42310 265650 42362
rect 265650 42310 265652 42362
rect 265596 42308 265652 42310
rect 265700 42362 265756 42364
rect 265700 42310 265702 42362
rect 265702 42310 265754 42362
rect 265754 42310 265756 42362
rect 265700 42308 265756 42310
rect 265804 42362 265860 42364
rect 265804 42310 265806 42362
rect 265806 42310 265858 42362
rect 265858 42310 265860 42362
rect 265804 42308 265860 42310
rect 265596 40794 265652 40796
rect 265596 40742 265598 40794
rect 265598 40742 265650 40794
rect 265650 40742 265652 40794
rect 265596 40740 265652 40742
rect 265700 40794 265756 40796
rect 265700 40742 265702 40794
rect 265702 40742 265754 40794
rect 265754 40742 265756 40794
rect 265700 40740 265756 40742
rect 265804 40794 265860 40796
rect 265804 40742 265806 40794
rect 265806 40742 265858 40794
rect 265858 40742 265860 40794
rect 265804 40740 265860 40742
rect 265596 39226 265652 39228
rect 265596 39174 265598 39226
rect 265598 39174 265650 39226
rect 265650 39174 265652 39226
rect 265596 39172 265652 39174
rect 265700 39226 265756 39228
rect 265700 39174 265702 39226
rect 265702 39174 265754 39226
rect 265754 39174 265756 39226
rect 265700 39172 265756 39174
rect 265804 39226 265860 39228
rect 265804 39174 265806 39226
rect 265806 39174 265858 39226
rect 265858 39174 265860 39226
rect 265804 39172 265860 39174
rect 265596 37658 265652 37660
rect 265596 37606 265598 37658
rect 265598 37606 265650 37658
rect 265650 37606 265652 37658
rect 265596 37604 265652 37606
rect 265700 37658 265756 37660
rect 265700 37606 265702 37658
rect 265702 37606 265754 37658
rect 265754 37606 265756 37658
rect 265700 37604 265756 37606
rect 265804 37658 265860 37660
rect 265804 37606 265806 37658
rect 265806 37606 265858 37658
rect 265858 37606 265860 37658
rect 265804 37604 265860 37606
rect 265596 36090 265652 36092
rect 265596 36038 265598 36090
rect 265598 36038 265650 36090
rect 265650 36038 265652 36090
rect 265596 36036 265652 36038
rect 265700 36090 265756 36092
rect 265700 36038 265702 36090
rect 265702 36038 265754 36090
rect 265754 36038 265756 36090
rect 265700 36036 265756 36038
rect 265804 36090 265860 36092
rect 265804 36038 265806 36090
rect 265806 36038 265858 36090
rect 265858 36038 265860 36090
rect 265804 36036 265860 36038
rect 265596 34522 265652 34524
rect 265596 34470 265598 34522
rect 265598 34470 265650 34522
rect 265650 34470 265652 34522
rect 265596 34468 265652 34470
rect 265700 34522 265756 34524
rect 265700 34470 265702 34522
rect 265702 34470 265754 34522
rect 265754 34470 265756 34522
rect 265700 34468 265756 34470
rect 265804 34522 265860 34524
rect 265804 34470 265806 34522
rect 265806 34470 265858 34522
rect 265858 34470 265860 34522
rect 265804 34468 265860 34470
rect 265596 32954 265652 32956
rect 265596 32902 265598 32954
rect 265598 32902 265650 32954
rect 265650 32902 265652 32954
rect 265596 32900 265652 32902
rect 265700 32954 265756 32956
rect 265700 32902 265702 32954
rect 265702 32902 265754 32954
rect 265754 32902 265756 32954
rect 265700 32900 265756 32902
rect 265804 32954 265860 32956
rect 265804 32902 265806 32954
rect 265806 32902 265858 32954
rect 265858 32902 265860 32954
rect 265804 32900 265860 32902
rect 265596 31386 265652 31388
rect 265596 31334 265598 31386
rect 265598 31334 265650 31386
rect 265650 31334 265652 31386
rect 265596 31332 265652 31334
rect 265700 31386 265756 31388
rect 265700 31334 265702 31386
rect 265702 31334 265754 31386
rect 265754 31334 265756 31386
rect 265700 31332 265756 31334
rect 265804 31386 265860 31388
rect 265804 31334 265806 31386
rect 265806 31334 265858 31386
rect 265858 31334 265860 31386
rect 265804 31332 265860 31334
rect 265596 29818 265652 29820
rect 265596 29766 265598 29818
rect 265598 29766 265650 29818
rect 265650 29766 265652 29818
rect 265596 29764 265652 29766
rect 265700 29818 265756 29820
rect 265700 29766 265702 29818
rect 265702 29766 265754 29818
rect 265754 29766 265756 29818
rect 265700 29764 265756 29766
rect 265804 29818 265860 29820
rect 265804 29766 265806 29818
rect 265806 29766 265858 29818
rect 265858 29766 265860 29818
rect 265804 29764 265860 29766
rect 265596 28250 265652 28252
rect 265596 28198 265598 28250
rect 265598 28198 265650 28250
rect 265650 28198 265652 28250
rect 265596 28196 265652 28198
rect 265700 28250 265756 28252
rect 265700 28198 265702 28250
rect 265702 28198 265754 28250
rect 265754 28198 265756 28250
rect 265700 28196 265756 28198
rect 265804 28250 265860 28252
rect 265804 28198 265806 28250
rect 265806 28198 265858 28250
rect 265858 28198 265860 28250
rect 265804 28196 265860 28198
rect 265596 26682 265652 26684
rect 265596 26630 265598 26682
rect 265598 26630 265650 26682
rect 265650 26630 265652 26682
rect 265596 26628 265652 26630
rect 265700 26682 265756 26684
rect 265700 26630 265702 26682
rect 265702 26630 265754 26682
rect 265754 26630 265756 26682
rect 265700 26628 265756 26630
rect 265804 26682 265860 26684
rect 265804 26630 265806 26682
rect 265806 26630 265858 26682
rect 265858 26630 265860 26682
rect 265804 26628 265860 26630
rect 265596 25114 265652 25116
rect 265596 25062 265598 25114
rect 265598 25062 265650 25114
rect 265650 25062 265652 25114
rect 265596 25060 265652 25062
rect 265700 25114 265756 25116
rect 265700 25062 265702 25114
rect 265702 25062 265754 25114
rect 265754 25062 265756 25114
rect 265700 25060 265756 25062
rect 265804 25114 265860 25116
rect 265804 25062 265806 25114
rect 265806 25062 265858 25114
rect 265858 25062 265860 25114
rect 265804 25060 265860 25062
rect 265596 23546 265652 23548
rect 265596 23494 265598 23546
rect 265598 23494 265650 23546
rect 265650 23494 265652 23546
rect 265596 23492 265652 23494
rect 265700 23546 265756 23548
rect 265700 23494 265702 23546
rect 265702 23494 265754 23546
rect 265754 23494 265756 23546
rect 265700 23492 265756 23494
rect 265804 23546 265860 23548
rect 265804 23494 265806 23546
rect 265806 23494 265858 23546
rect 265858 23494 265860 23546
rect 265804 23492 265860 23494
rect 265596 21978 265652 21980
rect 265596 21926 265598 21978
rect 265598 21926 265650 21978
rect 265650 21926 265652 21978
rect 265596 21924 265652 21926
rect 265700 21978 265756 21980
rect 265700 21926 265702 21978
rect 265702 21926 265754 21978
rect 265754 21926 265756 21978
rect 265700 21924 265756 21926
rect 265804 21978 265860 21980
rect 265804 21926 265806 21978
rect 265806 21926 265858 21978
rect 265858 21926 265860 21978
rect 265804 21924 265860 21926
rect 265596 20410 265652 20412
rect 265596 20358 265598 20410
rect 265598 20358 265650 20410
rect 265650 20358 265652 20410
rect 265596 20356 265652 20358
rect 265700 20410 265756 20412
rect 265700 20358 265702 20410
rect 265702 20358 265754 20410
rect 265754 20358 265756 20410
rect 265700 20356 265756 20358
rect 265804 20410 265860 20412
rect 265804 20358 265806 20410
rect 265806 20358 265858 20410
rect 265858 20358 265860 20410
rect 265804 20356 265860 20358
rect 265596 18842 265652 18844
rect 265596 18790 265598 18842
rect 265598 18790 265650 18842
rect 265650 18790 265652 18842
rect 265596 18788 265652 18790
rect 265700 18842 265756 18844
rect 265700 18790 265702 18842
rect 265702 18790 265754 18842
rect 265754 18790 265756 18842
rect 265700 18788 265756 18790
rect 265804 18842 265860 18844
rect 265804 18790 265806 18842
rect 265806 18790 265858 18842
rect 265858 18790 265860 18842
rect 265804 18788 265860 18790
rect 265596 17274 265652 17276
rect 265596 17222 265598 17274
rect 265598 17222 265650 17274
rect 265650 17222 265652 17274
rect 265596 17220 265652 17222
rect 265700 17274 265756 17276
rect 265700 17222 265702 17274
rect 265702 17222 265754 17274
rect 265754 17222 265756 17274
rect 265700 17220 265756 17222
rect 265804 17274 265860 17276
rect 265804 17222 265806 17274
rect 265806 17222 265858 17274
rect 265858 17222 265860 17274
rect 265804 17220 265860 17222
rect 264572 15932 264628 15988
rect 265596 15706 265652 15708
rect 265596 15654 265598 15706
rect 265598 15654 265650 15706
rect 265650 15654 265652 15706
rect 265596 15652 265652 15654
rect 265700 15706 265756 15708
rect 265700 15654 265702 15706
rect 265702 15654 265754 15706
rect 265754 15654 265756 15706
rect 265700 15652 265756 15654
rect 265804 15706 265860 15708
rect 265804 15654 265806 15706
rect 265806 15654 265858 15706
rect 265858 15654 265860 15706
rect 265804 15652 265860 15654
rect 265596 14138 265652 14140
rect 265596 14086 265598 14138
rect 265598 14086 265650 14138
rect 265650 14086 265652 14138
rect 265596 14084 265652 14086
rect 265700 14138 265756 14140
rect 265700 14086 265702 14138
rect 265702 14086 265754 14138
rect 265754 14086 265756 14138
rect 265700 14084 265756 14086
rect 265804 14138 265860 14140
rect 265804 14086 265806 14138
rect 265806 14086 265858 14138
rect 265858 14086 265860 14138
rect 265804 14084 265860 14086
rect 277228 55970 277284 55972
rect 277228 55918 277230 55970
rect 277230 55918 277282 55970
rect 277282 55918 277284 55970
rect 277228 55916 277284 55918
rect 279692 55916 279748 55972
rect 273196 12796 273252 12852
rect 281820 55970 281876 55972
rect 281820 55918 281822 55970
rect 281822 55918 281874 55970
rect 281874 55918 281876 55970
rect 281820 55916 281876 55918
rect 280956 55690 281012 55692
rect 280956 55638 280958 55690
rect 280958 55638 281010 55690
rect 281010 55638 281012 55690
rect 280956 55636 281012 55638
rect 281060 55690 281116 55692
rect 281060 55638 281062 55690
rect 281062 55638 281114 55690
rect 281114 55638 281116 55690
rect 281060 55636 281116 55638
rect 281164 55690 281220 55692
rect 281164 55638 281166 55690
rect 281166 55638 281218 55690
rect 281218 55638 281220 55690
rect 281164 55636 281220 55638
rect 280956 54122 281012 54124
rect 280956 54070 280958 54122
rect 280958 54070 281010 54122
rect 281010 54070 281012 54122
rect 280956 54068 281012 54070
rect 281060 54122 281116 54124
rect 281060 54070 281062 54122
rect 281062 54070 281114 54122
rect 281114 54070 281116 54122
rect 281060 54068 281116 54070
rect 281164 54122 281220 54124
rect 281164 54070 281166 54122
rect 281166 54070 281218 54122
rect 281218 54070 281220 54122
rect 281164 54068 281220 54070
rect 280956 52554 281012 52556
rect 280956 52502 280958 52554
rect 280958 52502 281010 52554
rect 281010 52502 281012 52554
rect 280956 52500 281012 52502
rect 281060 52554 281116 52556
rect 281060 52502 281062 52554
rect 281062 52502 281114 52554
rect 281114 52502 281116 52554
rect 281060 52500 281116 52502
rect 281164 52554 281220 52556
rect 281164 52502 281166 52554
rect 281166 52502 281218 52554
rect 281218 52502 281220 52554
rect 281164 52500 281220 52502
rect 280956 50986 281012 50988
rect 280956 50934 280958 50986
rect 280958 50934 281010 50986
rect 281010 50934 281012 50986
rect 280956 50932 281012 50934
rect 281060 50986 281116 50988
rect 281060 50934 281062 50986
rect 281062 50934 281114 50986
rect 281114 50934 281116 50986
rect 281060 50932 281116 50934
rect 281164 50986 281220 50988
rect 281164 50934 281166 50986
rect 281166 50934 281218 50986
rect 281218 50934 281220 50986
rect 281164 50932 281220 50934
rect 280956 49418 281012 49420
rect 280956 49366 280958 49418
rect 280958 49366 281010 49418
rect 281010 49366 281012 49418
rect 280956 49364 281012 49366
rect 281060 49418 281116 49420
rect 281060 49366 281062 49418
rect 281062 49366 281114 49418
rect 281114 49366 281116 49418
rect 281060 49364 281116 49366
rect 281164 49418 281220 49420
rect 281164 49366 281166 49418
rect 281166 49366 281218 49418
rect 281218 49366 281220 49418
rect 281164 49364 281220 49366
rect 280956 47850 281012 47852
rect 280956 47798 280958 47850
rect 280958 47798 281010 47850
rect 281010 47798 281012 47850
rect 280956 47796 281012 47798
rect 281060 47850 281116 47852
rect 281060 47798 281062 47850
rect 281062 47798 281114 47850
rect 281114 47798 281116 47850
rect 281060 47796 281116 47798
rect 281164 47850 281220 47852
rect 281164 47798 281166 47850
rect 281166 47798 281218 47850
rect 281218 47798 281220 47850
rect 281164 47796 281220 47798
rect 280956 46282 281012 46284
rect 280956 46230 280958 46282
rect 280958 46230 281010 46282
rect 281010 46230 281012 46282
rect 280956 46228 281012 46230
rect 281060 46282 281116 46284
rect 281060 46230 281062 46282
rect 281062 46230 281114 46282
rect 281114 46230 281116 46282
rect 281060 46228 281116 46230
rect 281164 46282 281220 46284
rect 281164 46230 281166 46282
rect 281166 46230 281218 46282
rect 281218 46230 281220 46282
rect 281164 46228 281220 46230
rect 280956 44714 281012 44716
rect 280956 44662 280958 44714
rect 280958 44662 281010 44714
rect 281010 44662 281012 44714
rect 280956 44660 281012 44662
rect 281060 44714 281116 44716
rect 281060 44662 281062 44714
rect 281062 44662 281114 44714
rect 281114 44662 281116 44714
rect 281060 44660 281116 44662
rect 281164 44714 281220 44716
rect 281164 44662 281166 44714
rect 281166 44662 281218 44714
rect 281218 44662 281220 44714
rect 281164 44660 281220 44662
rect 280956 43146 281012 43148
rect 280956 43094 280958 43146
rect 280958 43094 281010 43146
rect 281010 43094 281012 43146
rect 280956 43092 281012 43094
rect 281060 43146 281116 43148
rect 281060 43094 281062 43146
rect 281062 43094 281114 43146
rect 281114 43094 281116 43146
rect 281060 43092 281116 43094
rect 281164 43146 281220 43148
rect 281164 43094 281166 43146
rect 281166 43094 281218 43146
rect 281218 43094 281220 43146
rect 281164 43092 281220 43094
rect 280956 41578 281012 41580
rect 280956 41526 280958 41578
rect 280958 41526 281010 41578
rect 281010 41526 281012 41578
rect 280956 41524 281012 41526
rect 281060 41578 281116 41580
rect 281060 41526 281062 41578
rect 281062 41526 281114 41578
rect 281114 41526 281116 41578
rect 281060 41524 281116 41526
rect 281164 41578 281220 41580
rect 281164 41526 281166 41578
rect 281166 41526 281218 41578
rect 281218 41526 281220 41578
rect 281164 41524 281220 41526
rect 280956 40010 281012 40012
rect 280956 39958 280958 40010
rect 280958 39958 281010 40010
rect 281010 39958 281012 40010
rect 280956 39956 281012 39958
rect 281060 40010 281116 40012
rect 281060 39958 281062 40010
rect 281062 39958 281114 40010
rect 281114 39958 281116 40010
rect 281060 39956 281116 39958
rect 281164 40010 281220 40012
rect 281164 39958 281166 40010
rect 281166 39958 281218 40010
rect 281218 39958 281220 40010
rect 281164 39956 281220 39958
rect 280956 38442 281012 38444
rect 280956 38390 280958 38442
rect 280958 38390 281010 38442
rect 281010 38390 281012 38442
rect 280956 38388 281012 38390
rect 281060 38442 281116 38444
rect 281060 38390 281062 38442
rect 281062 38390 281114 38442
rect 281114 38390 281116 38442
rect 281060 38388 281116 38390
rect 281164 38442 281220 38444
rect 281164 38390 281166 38442
rect 281166 38390 281218 38442
rect 281218 38390 281220 38442
rect 281164 38388 281220 38390
rect 280956 36874 281012 36876
rect 280956 36822 280958 36874
rect 280958 36822 281010 36874
rect 281010 36822 281012 36874
rect 280956 36820 281012 36822
rect 281060 36874 281116 36876
rect 281060 36822 281062 36874
rect 281062 36822 281114 36874
rect 281114 36822 281116 36874
rect 281060 36820 281116 36822
rect 281164 36874 281220 36876
rect 281164 36822 281166 36874
rect 281166 36822 281218 36874
rect 281218 36822 281220 36874
rect 281164 36820 281220 36822
rect 280956 35306 281012 35308
rect 280956 35254 280958 35306
rect 280958 35254 281010 35306
rect 281010 35254 281012 35306
rect 280956 35252 281012 35254
rect 281060 35306 281116 35308
rect 281060 35254 281062 35306
rect 281062 35254 281114 35306
rect 281114 35254 281116 35306
rect 281060 35252 281116 35254
rect 281164 35306 281220 35308
rect 281164 35254 281166 35306
rect 281166 35254 281218 35306
rect 281218 35254 281220 35306
rect 281164 35252 281220 35254
rect 280956 33738 281012 33740
rect 280956 33686 280958 33738
rect 280958 33686 281010 33738
rect 281010 33686 281012 33738
rect 280956 33684 281012 33686
rect 281060 33738 281116 33740
rect 281060 33686 281062 33738
rect 281062 33686 281114 33738
rect 281114 33686 281116 33738
rect 281060 33684 281116 33686
rect 281164 33738 281220 33740
rect 281164 33686 281166 33738
rect 281166 33686 281218 33738
rect 281218 33686 281220 33738
rect 281164 33684 281220 33686
rect 280956 32170 281012 32172
rect 280956 32118 280958 32170
rect 280958 32118 281010 32170
rect 281010 32118 281012 32170
rect 280956 32116 281012 32118
rect 281060 32170 281116 32172
rect 281060 32118 281062 32170
rect 281062 32118 281114 32170
rect 281114 32118 281116 32170
rect 281060 32116 281116 32118
rect 281164 32170 281220 32172
rect 281164 32118 281166 32170
rect 281166 32118 281218 32170
rect 281218 32118 281220 32170
rect 281164 32116 281220 32118
rect 280956 30602 281012 30604
rect 280956 30550 280958 30602
rect 280958 30550 281010 30602
rect 281010 30550 281012 30602
rect 280956 30548 281012 30550
rect 281060 30602 281116 30604
rect 281060 30550 281062 30602
rect 281062 30550 281114 30602
rect 281114 30550 281116 30602
rect 281060 30548 281116 30550
rect 281164 30602 281220 30604
rect 281164 30550 281166 30602
rect 281166 30550 281218 30602
rect 281218 30550 281220 30602
rect 281164 30548 281220 30550
rect 280956 29034 281012 29036
rect 280956 28982 280958 29034
rect 280958 28982 281010 29034
rect 281010 28982 281012 29034
rect 280956 28980 281012 28982
rect 281060 29034 281116 29036
rect 281060 28982 281062 29034
rect 281062 28982 281114 29034
rect 281114 28982 281116 29034
rect 281060 28980 281116 28982
rect 281164 29034 281220 29036
rect 281164 28982 281166 29034
rect 281166 28982 281218 29034
rect 281218 28982 281220 29034
rect 281164 28980 281220 28982
rect 288092 27692 288148 27748
rect 280956 27466 281012 27468
rect 280956 27414 280958 27466
rect 280958 27414 281010 27466
rect 281010 27414 281012 27466
rect 280956 27412 281012 27414
rect 281060 27466 281116 27468
rect 281060 27414 281062 27466
rect 281062 27414 281114 27466
rect 281114 27414 281116 27466
rect 281060 27412 281116 27414
rect 281164 27466 281220 27468
rect 281164 27414 281166 27466
rect 281166 27414 281218 27466
rect 281218 27414 281220 27466
rect 281164 27412 281220 27414
rect 280956 25898 281012 25900
rect 280956 25846 280958 25898
rect 280958 25846 281010 25898
rect 281010 25846 281012 25898
rect 280956 25844 281012 25846
rect 281060 25898 281116 25900
rect 281060 25846 281062 25898
rect 281062 25846 281114 25898
rect 281114 25846 281116 25898
rect 281060 25844 281116 25846
rect 281164 25898 281220 25900
rect 281164 25846 281166 25898
rect 281166 25846 281218 25898
rect 281218 25846 281220 25898
rect 281164 25844 281220 25846
rect 280956 24330 281012 24332
rect 280956 24278 280958 24330
rect 280958 24278 281010 24330
rect 281010 24278 281012 24330
rect 280956 24276 281012 24278
rect 281060 24330 281116 24332
rect 281060 24278 281062 24330
rect 281062 24278 281114 24330
rect 281114 24278 281116 24330
rect 281060 24276 281116 24278
rect 281164 24330 281220 24332
rect 281164 24278 281166 24330
rect 281166 24278 281218 24330
rect 281218 24278 281220 24330
rect 281164 24276 281220 24278
rect 280956 22762 281012 22764
rect 280956 22710 280958 22762
rect 280958 22710 281010 22762
rect 281010 22710 281012 22762
rect 280956 22708 281012 22710
rect 281060 22762 281116 22764
rect 281060 22710 281062 22762
rect 281062 22710 281114 22762
rect 281114 22710 281116 22762
rect 281060 22708 281116 22710
rect 281164 22762 281220 22764
rect 281164 22710 281166 22762
rect 281166 22710 281218 22762
rect 281218 22710 281220 22762
rect 281164 22708 281220 22710
rect 280956 21194 281012 21196
rect 280956 21142 280958 21194
rect 280958 21142 281010 21194
rect 281010 21142 281012 21194
rect 280956 21140 281012 21142
rect 281060 21194 281116 21196
rect 281060 21142 281062 21194
rect 281062 21142 281114 21194
rect 281114 21142 281116 21194
rect 281060 21140 281116 21142
rect 281164 21194 281220 21196
rect 281164 21142 281166 21194
rect 281166 21142 281218 21194
rect 281218 21142 281220 21194
rect 281164 21140 281220 21142
rect 296316 54906 296372 54908
rect 296316 54854 296318 54906
rect 296318 54854 296370 54906
rect 296370 54854 296372 54906
rect 296316 54852 296372 54854
rect 296420 54906 296476 54908
rect 296420 54854 296422 54906
rect 296422 54854 296474 54906
rect 296474 54854 296476 54906
rect 296420 54852 296476 54854
rect 296524 54906 296580 54908
rect 296524 54854 296526 54906
rect 296526 54854 296578 54906
rect 296578 54854 296580 54906
rect 296524 54852 296580 54854
rect 296316 53338 296372 53340
rect 296316 53286 296318 53338
rect 296318 53286 296370 53338
rect 296370 53286 296372 53338
rect 296316 53284 296372 53286
rect 296420 53338 296476 53340
rect 296420 53286 296422 53338
rect 296422 53286 296474 53338
rect 296474 53286 296476 53338
rect 296420 53284 296476 53286
rect 296524 53338 296580 53340
rect 296524 53286 296526 53338
rect 296526 53286 296578 53338
rect 296578 53286 296580 53338
rect 296524 53284 296580 53286
rect 296316 51770 296372 51772
rect 296316 51718 296318 51770
rect 296318 51718 296370 51770
rect 296370 51718 296372 51770
rect 296316 51716 296372 51718
rect 296420 51770 296476 51772
rect 296420 51718 296422 51770
rect 296422 51718 296474 51770
rect 296474 51718 296476 51770
rect 296420 51716 296476 51718
rect 296524 51770 296580 51772
rect 296524 51718 296526 51770
rect 296526 51718 296578 51770
rect 296578 51718 296580 51770
rect 296524 51716 296580 51718
rect 296316 50202 296372 50204
rect 296316 50150 296318 50202
rect 296318 50150 296370 50202
rect 296370 50150 296372 50202
rect 296316 50148 296372 50150
rect 296420 50202 296476 50204
rect 296420 50150 296422 50202
rect 296422 50150 296474 50202
rect 296474 50150 296476 50202
rect 296420 50148 296476 50150
rect 296524 50202 296580 50204
rect 296524 50150 296526 50202
rect 296526 50150 296578 50202
rect 296578 50150 296580 50202
rect 296524 50148 296580 50150
rect 296316 48634 296372 48636
rect 296316 48582 296318 48634
rect 296318 48582 296370 48634
rect 296370 48582 296372 48634
rect 296316 48580 296372 48582
rect 296420 48634 296476 48636
rect 296420 48582 296422 48634
rect 296422 48582 296474 48634
rect 296474 48582 296476 48634
rect 296420 48580 296476 48582
rect 296524 48634 296580 48636
rect 296524 48582 296526 48634
rect 296526 48582 296578 48634
rect 296578 48582 296580 48634
rect 296524 48580 296580 48582
rect 296316 47066 296372 47068
rect 296316 47014 296318 47066
rect 296318 47014 296370 47066
rect 296370 47014 296372 47066
rect 296316 47012 296372 47014
rect 296420 47066 296476 47068
rect 296420 47014 296422 47066
rect 296422 47014 296474 47066
rect 296474 47014 296476 47066
rect 296420 47012 296476 47014
rect 296524 47066 296580 47068
rect 296524 47014 296526 47066
rect 296526 47014 296578 47066
rect 296578 47014 296580 47066
rect 296524 47012 296580 47014
rect 296316 45498 296372 45500
rect 296316 45446 296318 45498
rect 296318 45446 296370 45498
rect 296370 45446 296372 45498
rect 296316 45444 296372 45446
rect 296420 45498 296476 45500
rect 296420 45446 296422 45498
rect 296422 45446 296474 45498
rect 296474 45446 296476 45498
rect 296420 45444 296476 45446
rect 296524 45498 296580 45500
rect 296524 45446 296526 45498
rect 296526 45446 296578 45498
rect 296578 45446 296580 45498
rect 296524 45444 296580 45446
rect 296316 43930 296372 43932
rect 296316 43878 296318 43930
rect 296318 43878 296370 43930
rect 296370 43878 296372 43930
rect 296316 43876 296372 43878
rect 296420 43930 296476 43932
rect 296420 43878 296422 43930
rect 296422 43878 296474 43930
rect 296474 43878 296476 43930
rect 296420 43876 296476 43878
rect 296524 43930 296580 43932
rect 296524 43878 296526 43930
rect 296526 43878 296578 43930
rect 296578 43878 296580 43930
rect 296524 43876 296580 43878
rect 296316 42362 296372 42364
rect 296316 42310 296318 42362
rect 296318 42310 296370 42362
rect 296370 42310 296372 42362
rect 296316 42308 296372 42310
rect 296420 42362 296476 42364
rect 296420 42310 296422 42362
rect 296422 42310 296474 42362
rect 296474 42310 296476 42362
rect 296420 42308 296476 42310
rect 296524 42362 296580 42364
rect 296524 42310 296526 42362
rect 296526 42310 296578 42362
rect 296578 42310 296580 42362
rect 296524 42308 296580 42310
rect 296316 40794 296372 40796
rect 296316 40742 296318 40794
rect 296318 40742 296370 40794
rect 296370 40742 296372 40794
rect 296316 40740 296372 40742
rect 296420 40794 296476 40796
rect 296420 40742 296422 40794
rect 296422 40742 296474 40794
rect 296474 40742 296476 40794
rect 296420 40740 296476 40742
rect 296524 40794 296580 40796
rect 296524 40742 296526 40794
rect 296526 40742 296578 40794
rect 296578 40742 296580 40794
rect 296524 40740 296580 40742
rect 296316 39226 296372 39228
rect 296316 39174 296318 39226
rect 296318 39174 296370 39226
rect 296370 39174 296372 39226
rect 296316 39172 296372 39174
rect 296420 39226 296476 39228
rect 296420 39174 296422 39226
rect 296422 39174 296474 39226
rect 296474 39174 296476 39226
rect 296420 39172 296476 39174
rect 296524 39226 296580 39228
rect 296524 39174 296526 39226
rect 296526 39174 296578 39226
rect 296578 39174 296580 39226
rect 296524 39172 296580 39174
rect 296316 37658 296372 37660
rect 296316 37606 296318 37658
rect 296318 37606 296370 37658
rect 296370 37606 296372 37658
rect 296316 37604 296372 37606
rect 296420 37658 296476 37660
rect 296420 37606 296422 37658
rect 296422 37606 296474 37658
rect 296474 37606 296476 37658
rect 296420 37604 296476 37606
rect 296524 37658 296580 37660
rect 296524 37606 296526 37658
rect 296526 37606 296578 37658
rect 296578 37606 296580 37658
rect 296524 37604 296580 37606
rect 296316 36090 296372 36092
rect 296316 36038 296318 36090
rect 296318 36038 296370 36090
rect 296370 36038 296372 36090
rect 296316 36036 296372 36038
rect 296420 36090 296476 36092
rect 296420 36038 296422 36090
rect 296422 36038 296474 36090
rect 296474 36038 296476 36090
rect 296420 36036 296476 36038
rect 296524 36090 296580 36092
rect 296524 36038 296526 36090
rect 296526 36038 296578 36090
rect 296578 36038 296580 36090
rect 296524 36036 296580 36038
rect 296316 34522 296372 34524
rect 296316 34470 296318 34522
rect 296318 34470 296370 34522
rect 296370 34470 296372 34522
rect 296316 34468 296372 34470
rect 296420 34522 296476 34524
rect 296420 34470 296422 34522
rect 296422 34470 296474 34522
rect 296474 34470 296476 34522
rect 296420 34468 296476 34470
rect 296524 34522 296580 34524
rect 296524 34470 296526 34522
rect 296526 34470 296578 34522
rect 296578 34470 296580 34522
rect 296524 34468 296580 34470
rect 296316 32954 296372 32956
rect 296316 32902 296318 32954
rect 296318 32902 296370 32954
rect 296370 32902 296372 32954
rect 296316 32900 296372 32902
rect 296420 32954 296476 32956
rect 296420 32902 296422 32954
rect 296422 32902 296474 32954
rect 296474 32902 296476 32954
rect 296420 32900 296476 32902
rect 296524 32954 296580 32956
rect 296524 32902 296526 32954
rect 296526 32902 296578 32954
rect 296578 32902 296580 32954
rect 296524 32900 296580 32902
rect 296316 31386 296372 31388
rect 296316 31334 296318 31386
rect 296318 31334 296370 31386
rect 296370 31334 296372 31386
rect 296316 31332 296372 31334
rect 296420 31386 296476 31388
rect 296420 31334 296422 31386
rect 296422 31334 296474 31386
rect 296474 31334 296476 31386
rect 296420 31332 296476 31334
rect 296524 31386 296580 31388
rect 296524 31334 296526 31386
rect 296526 31334 296578 31386
rect 296578 31334 296580 31386
rect 296524 31332 296580 31334
rect 296316 29818 296372 29820
rect 296316 29766 296318 29818
rect 296318 29766 296370 29818
rect 296370 29766 296372 29818
rect 296316 29764 296372 29766
rect 296420 29818 296476 29820
rect 296420 29766 296422 29818
rect 296422 29766 296474 29818
rect 296474 29766 296476 29818
rect 296420 29764 296476 29766
rect 296524 29818 296580 29820
rect 296524 29766 296526 29818
rect 296526 29766 296578 29818
rect 296578 29766 296580 29818
rect 296524 29764 296580 29766
rect 296316 28250 296372 28252
rect 296316 28198 296318 28250
rect 296318 28198 296370 28250
rect 296370 28198 296372 28250
rect 296316 28196 296372 28198
rect 296420 28250 296476 28252
rect 296420 28198 296422 28250
rect 296422 28198 296474 28250
rect 296474 28198 296476 28250
rect 296420 28196 296476 28198
rect 296524 28250 296580 28252
rect 296524 28198 296526 28250
rect 296526 28198 296578 28250
rect 296578 28198 296580 28250
rect 296524 28196 296580 28198
rect 296316 26682 296372 26684
rect 296316 26630 296318 26682
rect 296318 26630 296370 26682
rect 296370 26630 296372 26682
rect 296316 26628 296372 26630
rect 296420 26682 296476 26684
rect 296420 26630 296422 26682
rect 296422 26630 296474 26682
rect 296474 26630 296476 26682
rect 296420 26628 296476 26630
rect 296524 26682 296580 26684
rect 296524 26630 296526 26682
rect 296526 26630 296578 26682
rect 296578 26630 296580 26682
rect 296524 26628 296580 26630
rect 296316 25114 296372 25116
rect 296316 25062 296318 25114
rect 296318 25062 296370 25114
rect 296370 25062 296372 25114
rect 296316 25060 296372 25062
rect 296420 25114 296476 25116
rect 296420 25062 296422 25114
rect 296422 25062 296474 25114
rect 296474 25062 296476 25114
rect 296420 25060 296476 25062
rect 296524 25114 296580 25116
rect 296524 25062 296526 25114
rect 296526 25062 296578 25114
rect 296578 25062 296580 25114
rect 296524 25060 296580 25062
rect 296316 23546 296372 23548
rect 296316 23494 296318 23546
rect 296318 23494 296370 23546
rect 296370 23494 296372 23546
rect 296316 23492 296372 23494
rect 296420 23546 296476 23548
rect 296420 23494 296422 23546
rect 296422 23494 296474 23546
rect 296474 23494 296476 23546
rect 296420 23492 296476 23494
rect 296524 23546 296580 23548
rect 296524 23494 296526 23546
rect 296526 23494 296578 23546
rect 296578 23494 296580 23546
rect 296524 23492 296580 23494
rect 296316 21978 296372 21980
rect 296316 21926 296318 21978
rect 296318 21926 296370 21978
rect 296370 21926 296372 21978
rect 296316 21924 296372 21926
rect 296420 21978 296476 21980
rect 296420 21926 296422 21978
rect 296422 21926 296474 21978
rect 296474 21926 296476 21978
rect 296420 21924 296476 21926
rect 296524 21978 296580 21980
rect 296524 21926 296526 21978
rect 296526 21926 296578 21978
rect 296578 21926 296580 21978
rect 296524 21924 296580 21926
rect 293356 20972 293412 21028
rect 296316 20410 296372 20412
rect 296316 20358 296318 20410
rect 296318 20358 296370 20410
rect 296370 20358 296372 20410
rect 296316 20356 296372 20358
rect 296420 20410 296476 20412
rect 296420 20358 296422 20410
rect 296422 20358 296474 20410
rect 296474 20358 296476 20410
rect 296420 20356 296476 20358
rect 296524 20410 296580 20412
rect 296524 20358 296526 20410
rect 296526 20358 296578 20410
rect 296578 20358 296580 20410
rect 296524 20356 296580 20358
rect 280956 19626 281012 19628
rect 280956 19574 280958 19626
rect 280958 19574 281010 19626
rect 281010 19574 281012 19626
rect 280956 19572 281012 19574
rect 281060 19626 281116 19628
rect 281060 19574 281062 19626
rect 281062 19574 281114 19626
rect 281114 19574 281116 19626
rect 281060 19572 281116 19574
rect 281164 19626 281220 19628
rect 281164 19574 281166 19626
rect 281166 19574 281218 19626
rect 281218 19574 281220 19626
rect 281164 19572 281220 19574
rect 296316 18842 296372 18844
rect 296316 18790 296318 18842
rect 296318 18790 296370 18842
rect 296370 18790 296372 18842
rect 296316 18788 296372 18790
rect 296420 18842 296476 18844
rect 296420 18790 296422 18842
rect 296422 18790 296474 18842
rect 296474 18790 296476 18842
rect 296420 18788 296476 18790
rect 296524 18842 296580 18844
rect 296524 18790 296526 18842
rect 296526 18790 296578 18842
rect 296578 18790 296580 18842
rect 296524 18788 296580 18790
rect 280956 18058 281012 18060
rect 280956 18006 280958 18058
rect 280958 18006 281010 18058
rect 281010 18006 281012 18058
rect 280956 18004 281012 18006
rect 281060 18058 281116 18060
rect 281060 18006 281062 18058
rect 281062 18006 281114 18058
rect 281114 18006 281116 18058
rect 281060 18004 281116 18006
rect 281164 18058 281220 18060
rect 281164 18006 281166 18058
rect 281166 18006 281218 18058
rect 281218 18006 281220 18058
rect 281164 18004 281220 18006
rect 296316 17274 296372 17276
rect 296316 17222 296318 17274
rect 296318 17222 296370 17274
rect 296370 17222 296372 17274
rect 296316 17220 296372 17222
rect 296420 17274 296476 17276
rect 296420 17222 296422 17274
rect 296422 17222 296474 17274
rect 296474 17222 296476 17274
rect 296420 17220 296476 17222
rect 296524 17274 296580 17276
rect 296524 17222 296526 17274
rect 296526 17222 296578 17274
rect 296578 17222 296580 17274
rect 296524 17220 296580 17222
rect 280956 16490 281012 16492
rect 280956 16438 280958 16490
rect 280958 16438 281010 16490
rect 281010 16438 281012 16490
rect 280956 16436 281012 16438
rect 281060 16490 281116 16492
rect 281060 16438 281062 16490
rect 281062 16438 281114 16490
rect 281114 16438 281116 16490
rect 281060 16436 281116 16438
rect 281164 16490 281220 16492
rect 281164 16438 281166 16490
rect 281166 16438 281218 16490
rect 281218 16438 281220 16490
rect 281164 16436 281220 16438
rect 296316 15706 296372 15708
rect 296316 15654 296318 15706
rect 296318 15654 296370 15706
rect 296370 15654 296372 15706
rect 296316 15652 296372 15654
rect 296420 15706 296476 15708
rect 296420 15654 296422 15706
rect 296422 15654 296474 15706
rect 296474 15654 296476 15706
rect 296420 15652 296476 15654
rect 296524 15706 296580 15708
rect 296524 15654 296526 15706
rect 296526 15654 296578 15706
rect 296578 15654 296580 15706
rect 296524 15652 296580 15654
rect 280956 14922 281012 14924
rect 280956 14870 280958 14922
rect 280958 14870 281010 14922
rect 281010 14870 281012 14922
rect 280956 14868 281012 14870
rect 281060 14922 281116 14924
rect 281060 14870 281062 14922
rect 281062 14870 281114 14922
rect 281114 14870 281116 14922
rect 281060 14868 281116 14870
rect 281164 14922 281220 14924
rect 281164 14870 281166 14922
rect 281166 14870 281218 14922
rect 281218 14870 281220 14922
rect 281164 14868 281220 14870
rect 296316 14138 296372 14140
rect 296316 14086 296318 14138
rect 296318 14086 296370 14138
rect 296370 14086 296372 14138
rect 296316 14084 296372 14086
rect 296420 14138 296476 14140
rect 296420 14086 296422 14138
rect 296422 14086 296474 14138
rect 296474 14086 296476 14138
rect 296420 14084 296476 14086
rect 296524 14138 296580 14140
rect 296524 14086 296526 14138
rect 296526 14086 296578 14138
rect 296578 14086 296580 14138
rect 296524 14084 296580 14086
rect 280956 13354 281012 13356
rect 280956 13302 280958 13354
rect 280958 13302 281010 13354
rect 281010 13302 281012 13354
rect 280956 13300 281012 13302
rect 281060 13354 281116 13356
rect 281060 13302 281062 13354
rect 281062 13302 281114 13354
rect 281114 13302 281116 13354
rect 281060 13300 281116 13302
rect 281164 13354 281220 13356
rect 281164 13302 281166 13354
rect 281166 13302 281218 13354
rect 281218 13302 281220 13354
rect 281164 13300 281220 13302
rect 279692 12684 279748 12740
rect 265596 12570 265652 12572
rect 265596 12518 265598 12570
rect 265598 12518 265650 12570
rect 265650 12518 265652 12570
rect 265596 12516 265652 12518
rect 265700 12570 265756 12572
rect 265700 12518 265702 12570
rect 265702 12518 265754 12570
rect 265754 12518 265756 12570
rect 265700 12516 265756 12518
rect 265804 12570 265860 12572
rect 265804 12518 265806 12570
rect 265806 12518 265858 12570
rect 265858 12518 265860 12570
rect 265804 12516 265860 12518
rect 296316 12570 296372 12572
rect 296316 12518 296318 12570
rect 296318 12518 296370 12570
rect 296370 12518 296372 12570
rect 296316 12516 296372 12518
rect 296420 12570 296476 12572
rect 296420 12518 296422 12570
rect 296422 12518 296474 12570
rect 296474 12518 296476 12570
rect 296420 12516 296476 12518
rect 296524 12570 296580 12572
rect 296524 12518 296526 12570
rect 296526 12518 296578 12570
rect 296578 12518 296580 12570
rect 296524 12516 296580 12518
rect 280956 11786 281012 11788
rect 280956 11734 280958 11786
rect 280958 11734 281010 11786
rect 281010 11734 281012 11786
rect 280956 11732 281012 11734
rect 281060 11786 281116 11788
rect 281060 11734 281062 11786
rect 281062 11734 281114 11786
rect 281114 11734 281116 11786
rect 281060 11732 281116 11734
rect 281164 11786 281220 11788
rect 281164 11734 281166 11786
rect 281166 11734 281218 11786
rect 281218 11734 281220 11786
rect 281164 11732 281220 11734
rect 261772 11116 261828 11172
rect 234876 11002 234932 11004
rect 234876 10950 234878 11002
rect 234878 10950 234930 11002
rect 234930 10950 234932 11002
rect 234876 10948 234932 10950
rect 234980 11002 235036 11004
rect 234980 10950 234982 11002
rect 234982 10950 235034 11002
rect 235034 10950 235036 11002
rect 234980 10948 235036 10950
rect 235084 11002 235140 11004
rect 235084 10950 235086 11002
rect 235086 10950 235138 11002
rect 235138 10950 235140 11002
rect 235084 10948 235140 10950
rect 265596 11002 265652 11004
rect 265596 10950 265598 11002
rect 265598 10950 265650 11002
rect 265650 10950 265652 11002
rect 265596 10948 265652 10950
rect 265700 11002 265756 11004
rect 265700 10950 265702 11002
rect 265702 10950 265754 11002
rect 265754 10950 265756 11002
rect 265700 10948 265756 10950
rect 265804 11002 265860 11004
rect 265804 10950 265806 11002
rect 265806 10950 265858 11002
rect 265858 10950 265860 11002
rect 265804 10948 265860 10950
rect 296316 11002 296372 11004
rect 296316 10950 296318 11002
rect 296318 10950 296370 11002
rect 296370 10950 296372 11002
rect 296316 10948 296372 10950
rect 296420 11002 296476 11004
rect 296420 10950 296422 11002
rect 296422 10950 296474 11002
rect 296474 10950 296476 11002
rect 296420 10948 296476 10950
rect 296524 11002 296580 11004
rect 296524 10950 296526 11002
rect 296526 10950 296578 11002
rect 296578 10950 296580 11002
rect 296524 10948 296580 10950
rect 250236 10218 250292 10220
rect 250236 10166 250238 10218
rect 250238 10166 250290 10218
rect 250290 10166 250292 10218
rect 250236 10164 250292 10166
rect 250340 10218 250396 10220
rect 250340 10166 250342 10218
rect 250342 10166 250394 10218
rect 250394 10166 250396 10218
rect 250340 10164 250396 10166
rect 250444 10218 250500 10220
rect 250444 10166 250446 10218
rect 250446 10166 250498 10218
rect 250498 10166 250500 10218
rect 250444 10164 250500 10166
rect 280956 10218 281012 10220
rect 280956 10166 280958 10218
rect 280958 10166 281010 10218
rect 281010 10166 281012 10218
rect 280956 10164 281012 10166
rect 281060 10218 281116 10220
rect 281060 10166 281062 10218
rect 281062 10166 281114 10218
rect 281114 10166 281116 10218
rect 281060 10164 281116 10166
rect 281164 10218 281220 10220
rect 281164 10166 281166 10218
rect 281166 10166 281218 10218
rect 281218 10166 281220 10218
rect 281164 10164 281220 10166
rect 270620 9884 270676 9940
rect 234876 9434 234932 9436
rect 234876 9382 234878 9434
rect 234878 9382 234930 9434
rect 234930 9382 234932 9434
rect 234876 9380 234932 9382
rect 234980 9434 235036 9436
rect 234980 9382 234982 9434
rect 234982 9382 235034 9434
rect 235034 9382 235036 9434
rect 234980 9380 235036 9382
rect 235084 9434 235140 9436
rect 235084 9382 235086 9434
rect 235086 9382 235138 9434
rect 235138 9382 235140 9434
rect 235084 9380 235140 9382
rect 265596 9434 265652 9436
rect 265596 9382 265598 9434
rect 265598 9382 265650 9434
rect 265650 9382 265652 9434
rect 265596 9380 265652 9382
rect 265700 9434 265756 9436
rect 265700 9382 265702 9434
rect 265702 9382 265754 9434
rect 265754 9382 265756 9434
rect 265700 9380 265756 9382
rect 265804 9434 265860 9436
rect 265804 9382 265806 9434
rect 265806 9382 265858 9434
rect 265858 9382 265860 9434
rect 265804 9380 265860 9382
rect 250236 8650 250292 8652
rect 250236 8598 250238 8650
rect 250238 8598 250290 8650
rect 250290 8598 250292 8650
rect 250236 8596 250292 8598
rect 250340 8650 250396 8652
rect 250340 8598 250342 8650
rect 250342 8598 250394 8650
rect 250394 8598 250396 8650
rect 250340 8596 250396 8598
rect 250444 8650 250500 8652
rect 250444 8598 250446 8650
rect 250446 8598 250498 8650
rect 250498 8598 250500 8650
rect 250444 8596 250500 8598
rect 225932 8316 225988 8372
rect 234876 7866 234932 7868
rect 234876 7814 234878 7866
rect 234878 7814 234930 7866
rect 234930 7814 234932 7866
rect 234876 7812 234932 7814
rect 234980 7866 235036 7868
rect 234980 7814 234982 7866
rect 234982 7814 235034 7866
rect 235034 7814 235036 7866
rect 234980 7812 235036 7814
rect 235084 7866 235140 7868
rect 235084 7814 235086 7866
rect 235086 7814 235138 7866
rect 235138 7814 235140 7866
rect 235084 7812 235140 7814
rect 265596 7866 265652 7868
rect 265596 7814 265598 7866
rect 265598 7814 265650 7866
rect 265650 7814 265652 7866
rect 265596 7812 265652 7814
rect 265700 7866 265756 7868
rect 265700 7814 265702 7866
rect 265702 7814 265754 7866
rect 265754 7814 265756 7866
rect 265700 7812 265756 7814
rect 265804 7866 265860 7868
rect 265804 7814 265806 7866
rect 265806 7814 265858 7866
rect 265858 7814 265860 7866
rect 265804 7812 265860 7814
rect 221788 7644 221844 7700
rect 250236 7082 250292 7084
rect 250236 7030 250238 7082
rect 250238 7030 250290 7082
rect 250290 7030 250292 7082
rect 250236 7028 250292 7030
rect 250340 7082 250396 7084
rect 250340 7030 250342 7082
rect 250342 7030 250394 7082
rect 250394 7030 250396 7082
rect 250340 7028 250396 7030
rect 250444 7082 250500 7084
rect 250444 7030 250446 7082
rect 250446 7030 250498 7082
rect 250498 7030 250500 7082
rect 250444 7028 250500 7030
rect 234876 6298 234932 6300
rect 234876 6246 234878 6298
rect 234878 6246 234930 6298
rect 234930 6246 234932 6298
rect 234876 6244 234932 6246
rect 234980 6298 235036 6300
rect 234980 6246 234982 6298
rect 234982 6246 235034 6298
rect 235034 6246 235036 6298
rect 234980 6244 235036 6246
rect 235084 6298 235140 6300
rect 235084 6246 235086 6298
rect 235086 6246 235138 6298
rect 235138 6246 235140 6298
rect 235084 6244 235140 6246
rect 265596 6298 265652 6300
rect 265596 6246 265598 6298
rect 265598 6246 265650 6298
rect 265650 6246 265652 6298
rect 265596 6244 265652 6246
rect 265700 6298 265756 6300
rect 265700 6246 265702 6298
rect 265702 6246 265754 6298
rect 265754 6246 265756 6298
rect 265700 6244 265756 6246
rect 265804 6298 265860 6300
rect 265804 6246 265806 6298
rect 265806 6246 265858 6298
rect 265858 6246 265860 6298
rect 265804 6244 265860 6246
rect 263004 6076 263060 6132
rect 222572 5180 222628 5236
rect 221564 5122 221620 5124
rect 221564 5070 221566 5122
rect 221566 5070 221618 5122
rect 221618 5070 221620 5122
rect 221564 5068 221620 5070
rect 220892 3948 220948 4004
rect 220556 3612 220612 3668
rect 220444 3500 220500 3556
rect 220108 2716 220164 2772
rect 221788 4844 221844 4900
rect 222124 4844 222180 4900
rect 221900 4338 221956 4340
rect 221900 4286 221902 4338
rect 221902 4286 221954 4338
rect 221954 4286 221956 4338
rect 221900 4284 221956 4286
rect 221452 3612 221508 3668
rect 221228 3442 221284 3444
rect 221228 3390 221230 3442
rect 221230 3390 221282 3442
rect 221282 3390 221284 3442
rect 221228 3388 221284 3390
rect 223468 5180 223524 5236
rect 223132 4898 223188 4900
rect 223132 4846 223134 4898
rect 223134 4846 223186 4898
rect 223186 4846 223188 4898
rect 223132 4844 223188 4846
rect 234332 5740 234388 5796
rect 224028 5122 224084 5124
rect 224028 5070 224030 5122
rect 224030 5070 224082 5122
rect 224082 5070 224084 5122
rect 224028 5068 224084 5070
rect 223020 4732 223076 4788
rect 223244 4338 223300 4340
rect 223244 4286 223246 4338
rect 223246 4286 223298 4338
rect 223298 4286 223300 4338
rect 223244 4284 223300 4286
rect 223132 4226 223188 4228
rect 223132 4174 223134 4226
rect 223134 4174 223186 4226
rect 223186 4174 223188 4226
rect 223132 4172 223188 4174
rect 223916 4732 223972 4788
rect 223692 4338 223748 4340
rect 223692 4286 223694 4338
rect 223694 4286 223746 4338
rect 223746 4286 223748 4338
rect 223692 4284 223748 4286
rect 223356 4060 223412 4116
rect 230748 4508 230804 4564
rect 224700 3612 224756 3668
rect 228508 4396 228564 4452
rect 222012 2828 222068 2884
rect 223916 3500 223972 3556
rect 221116 2044 221172 2100
rect 225932 3500 225988 3556
rect 225932 2940 225988 2996
rect 227164 3330 227220 3332
rect 227164 3278 227166 3330
rect 227166 3278 227218 3330
rect 227218 3278 227220 3330
rect 227164 3276 227220 3278
rect 228508 2492 228564 2548
rect 250236 5514 250292 5516
rect 250236 5462 250238 5514
rect 250238 5462 250290 5514
rect 250290 5462 250292 5514
rect 250236 5460 250292 5462
rect 250340 5514 250396 5516
rect 250340 5462 250342 5514
rect 250342 5462 250394 5514
rect 250394 5462 250396 5514
rect 250340 5460 250396 5462
rect 250444 5514 250500 5516
rect 250444 5462 250446 5514
rect 250446 5462 250498 5514
rect 250498 5462 250500 5514
rect 250444 5460 250500 5462
rect 245420 5180 245476 5236
rect 241612 4956 241668 5012
rect 234876 4730 234932 4732
rect 234876 4678 234878 4730
rect 234878 4678 234930 4730
rect 234930 4678 234932 4730
rect 234876 4676 234932 4678
rect 234980 4730 235036 4732
rect 234980 4678 234982 4730
rect 234982 4678 235034 4730
rect 235034 4678 235036 4730
rect 234980 4676 235036 4678
rect 235084 4730 235140 4732
rect 235084 4678 235086 4730
rect 235086 4678 235138 4730
rect 235138 4678 235140 4730
rect 235084 4676 235140 4678
rect 237916 3724 237972 3780
rect 234876 3162 234932 3164
rect 234876 3110 234878 3162
rect 234878 3110 234930 3162
rect 234930 3110 234932 3162
rect 234876 3108 234932 3110
rect 234980 3162 235036 3164
rect 234980 3110 234982 3162
rect 234982 3110 235034 3162
rect 235034 3110 235036 3162
rect 234980 3108 235036 3110
rect 235084 3162 235140 3164
rect 235084 3110 235086 3162
rect 235086 3110 235138 3162
rect 235138 3110 235140 3162
rect 235084 3108 235140 3110
rect 244972 3442 245028 3444
rect 244972 3390 244974 3442
rect 244974 3390 245026 3442
rect 245026 3390 245028 3442
rect 244972 3388 245028 3390
rect 249228 4284 249284 4340
rect 245644 3388 245700 3444
rect 248780 3442 248836 3444
rect 248780 3390 248782 3442
rect 248782 3390 248834 3442
rect 248834 3390 248836 3442
rect 248780 3388 248836 3390
rect 253036 4060 253092 4116
rect 250236 3946 250292 3948
rect 250236 3894 250238 3946
rect 250238 3894 250290 3946
rect 250290 3894 250292 3946
rect 250236 3892 250292 3894
rect 250340 3946 250396 3948
rect 250340 3894 250342 3946
rect 250342 3894 250394 3946
rect 250394 3894 250396 3946
rect 250340 3892 250396 3894
rect 250444 3946 250500 3948
rect 250444 3894 250446 3946
rect 250446 3894 250498 3946
rect 250498 3894 250500 3946
rect 250444 3892 250500 3894
rect 249340 3612 249396 3668
rect 249452 3388 249508 3444
rect 255836 3724 255892 3780
rect 249340 1260 249396 1316
rect 259420 2716 259476 2772
rect 265596 4730 265652 4732
rect 265596 4678 265598 4730
rect 265598 4678 265650 4730
rect 265650 4678 265652 4730
rect 265596 4676 265652 4678
rect 265700 4730 265756 4732
rect 265700 4678 265702 4730
rect 265702 4678 265754 4730
rect 265754 4678 265756 4730
rect 265700 4676 265756 4678
rect 265804 4730 265860 4732
rect 265804 4678 265806 4730
rect 265806 4678 265858 4730
rect 265858 4678 265860 4730
rect 265804 4676 265860 4678
rect 265356 3388 265412 3444
rect 265596 3162 265652 3164
rect 265596 3110 265598 3162
rect 265598 3110 265650 3162
rect 265650 3110 265652 3162
rect 265596 3108 265652 3110
rect 265700 3162 265756 3164
rect 265700 3110 265702 3162
rect 265702 3110 265754 3162
rect 265754 3110 265756 3162
rect 265700 3108 265756 3110
rect 265804 3162 265860 3164
rect 265804 3110 265806 3162
rect 265806 3110 265858 3162
rect 265858 3110 265860 3162
rect 265804 3108 265860 3110
rect 265356 1596 265412 1652
rect 296316 9434 296372 9436
rect 296316 9382 296318 9434
rect 296318 9382 296370 9434
rect 296370 9382 296372 9434
rect 296316 9380 296372 9382
rect 296420 9434 296476 9436
rect 296420 9382 296422 9434
rect 296422 9382 296474 9434
rect 296474 9382 296476 9434
rect 296420 9380 296476 9382
rect 296524 9434 296580 9436
rect 296524 9382 296526 9434
rect 296526 9382 296578 9434
rect 296578 9382 296580 9434
rect 296524 9380 296580 9382
rect 280956 8650 281012 8652
rect 280956 8598 280958 8650
rect 280958 8598 281010 8650
rect 281010 8598 281012 8650
rect 280956 8596 281012 8598
rect 281060 8650 281116 8652
rect 281060 8598 281062 8650
rect 281062 8598 281114 8650
rect 281114 8598 281116 8650
rect 281060 8596 281116 8598
rect 281164 8650 281220 8652
rect 281164 8598 281166 8650
rect 281166 8598 281218 8650
rect 281218 8598 281220 8650
rect 281164 8596 281220 8598
rect 296316 7866 296372 7868
rect 296316 7814 296318 7866
rect 296318 7814 296370 7866
rect 296370 7814 296372 7866
rect 296316 7812 296372 7814
rect 296420 7866 296476 7868
rect 296420 7814 296422 7866
rect 296422 7814 296474 7866
rect 296474 7814 296476 7866
rect 296420 7812 296476 7814
rect 296524 7866 296580 7868
rect 296524 7814 296526 7866
rect 296526 7814 296578 7866
rect 296578 7814 296580 7866
rect 296524 7812 296580 7814
rect 280956 7082 281012 7084
rect 280956 7030 280958 7082
rect 280958 7030 281010 7082
rect 281010 7030 281012 7082
rect 280956 7028 281012 7030
rect 281060 7082 281116 7084
rect 281060 7030 281062 7082
rect 281062 7030 281114 7082
rect 281114 7030 281116 7082
rect 281060 7028 281116 7030
rect 281164 7082 281220 7084
rect 281164 7030 281166 7082
rect 281166 7030 281218 7082
rect 281218 7030 281220 7082
rect 281164 7028 281220 7030
rect 296316 6298 296372 6300
rect 296316 6246 296318 6298
rect 296318 6246 296370 6298
rect 296370 6246 296372 6298
rect 296316 6244 296372 6246
rect 296420 6298 296476 6300
rect 296420 6246 296422 6298
rect 296422 6246 296474 6298
rect 296474 6246 296476 6298
rect 296420 6244 296476 6246
rect 296524 6298 296580 6300
rect 296524 6246 296526 6298
rect 296526 6246 296578 6298
rect 296578 6246 296580 6298
rect 296524 6244 296580 6246
rect 292124 5964 292180 6020
rect 280956 5514 281012 5516
rect 280956 5462 280958 5514
rect 280958 5462 281010 5514
rect 281010 5462 281012 5514
rect 280956 5460 281012 5462
rect 281060 5514 281116 5516
rect 281060 5462 281062 5514
rect 281062 5462 281114 5514
rect 281114 5462 281116 5514
rect 281060 5460 281116 5462
rect 281164 5514 281220 5516
rect 281164 5462 281166 5514
rect 281166 5462 281218 5514
rect 281218 5462 281220 5514
rect 281164 5460 281220 5462
rect 288540 4396 288596 4452
rect 280956 3946 281012 3948
rect 280956 3894 280958 3946
rect 280958 3894 281010 3946
rect 281010 3894 281012 3946
rect 280956 3892 281012 3894
rect 281060 3946 281116 3948
rect 281060 3894 281062 3946
rect 281062 3894 281114 3946
rect 281114 3894 281116 3946
rect 281060 3892 281116 3894
rect 281164 3946 281220 3948
rect 281164 3894 281166 3946
rect 281166 3894 281218 3946
rect 281218 3894 281220 3946
rect 281164 3892 281220 3894
rect 281372 3724 281428 3780
rect 296316 4730 296372 4732
rect 296316 4678 296318 4730
rect 296318 4678 296370 4730
rect 296370 4678 296372 4730
rect 296316 4676 296372 4678
rect 296420 4730 296476 4732
rect 296420 4678 296422 4730
rect 296422 4678 296474 4730
rect 296474 4678 296476 4730
rect 296420 4676 296476 4678
rect 296524 4730 296580 4732
rect 296524 4678 296526 4730
rect 296526 4678 296578 4730
rect 296578 4678 296580 4730
rect 296524 4676 296580 4678
rect 285068 3554 285124 3556
rect 285068 3502 285070 3554
rect 285070 3502 285122 3554
rect 285122 3502 285124 3554
rect 285068 3500 285124 3502
rect 267036 3388 267092 3444
rect 274316 1372 274372 1428
rect 277900 3276 277956 3332
rect 296316 3162 296372 3164
rect 296316 3110 296318 3162
rect 296318 3110 296370 3162
rect 296370 3110 296372 3162
rect 296316 3108 296372 3110
rect 296420 3162 296476 3164
rect 296420 3110 296422 3162
rect 296422 3110 296474 3162
rect 296474 3110 296476 3162
rect 296420 3108 296476 3110
rect 296524 3162 296580 3164
rect 296524 3110 296526 3162
rect 296526 3110 296578 3162
rect 296578 3110 296580 3162
rect 296524 3108 296580 3110
<< metal3 >>
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 81266 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81550 56476
rect 111986 56420 111996 56476
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 112260 56420 112270 56476
rect 142706 56420 142716 56476
rect 142772 56420 142820 56476
rect 142876 56420 142924 56476
rect 142980 56420 142990 56476
rect 173426 56420 173436 56476
rect 173492 56420 173540 56476
rect 173596 56420 173644 56476
rect 173700 56420 173710 56476
rect 204146 56420 204156 56476
rect 204212 56420 204260 56476
rect 204316 56420 204364 56476
rect 204420 56420 204430 56476
rect 234866 56420 234876 56476
rect 234932 56420 234980 56476
rect 235036 56420 235084 56476
rect 235140 56420 235150 56476
rect 265586 56420 265596 56476
rect 265652 56420 265700 56476
rect 265756 56420 265804 56476
rect 265860 56420 265870 56476
rect 296306 56420 296316 56476
rect 296372 56420 296420 56476
rect 296476 56420 296524 56476
rect 296580 56420 296590 56476
rect 19170 56252 19180 56308
rect 19236 56252 173068 56308
rect 206322 56252 206332 56308
rect 206388 56252 208348 56308
rect 208404 56252 208414 56308
rect 233538 56252 233548 56308
rect 233604 56252 234220 56308
rect 234276 56252 234286 56308
rect 126242 56140 126252 56196
rect 126308 56140 127820 56196
rect 127876 56140 127886 56196
rect 135762 56140 135772 56196
rect 135828 56140 136668 56196
rect 136724 56140 136734 56196
rect 142146 56140 142156 56196
rect 142212 56140 142828 56196
rect 142884 56140 142894 56196
rect 84914 56028 84924 56084
rect 84980 56028 85708 56084
rect 85764 56028 85774 56084
rect 173012 55972 173068 56252
rect 184034 56140 184044 56196
rect 184100 56140 185052 56196
rect 185108 56140 185118 56196
rect 187170 56140 187180 56196
rect 187236 56140 189868 56196
rect 189924 56140 189934 56196
rect 193890 56140 193900 56196
rect 193956 56140 195916 56196
rect 195972 56140 195982 56196
rect 190866 56028 190876 56084
rect 190932 56028 191772 56084
rect 191828 56028 191838 56084
rect 260082 56028 260092 56084
rect 260148 56028 260764 56084
rect 260820 56028 260830 56084
rect 271506 56028 271516 56084
rect 271572 56028 272188 56084
rect 272244 56028 272254 56084
rect 281586 56028 281596 56084
rect 281652 56028 282716 56084
rect 282772 56028 283612 56084
rect 283668 56028 283678 56084
rect 51762 55916 51772 55972
rect 51828 55916 52892 55972
rect 52948 55916 52958 55972
rect 69346 55916 69356 55972
rect 69412 55916 70476 55972
rect 70532 55916 73052 55972
rect 73108 55916 73118 55972
rect 80434 55916 80444 55972
rect 80500 55916 81004 55972
rect 81060 55916 83132 55972
rect 83188 55916 83198 55972
rect 88050 55916 88060 55972
rect 88116 55916 89516 55972
rect 89572 55916 89582 55972
rect 96226 55916 96236 55972
rect 96292 55916 97132 55972
rect 97188 55916 99932 55972
rect 99988 55916 99998 55972
rect 121090 55916 121100 55972
rect 121156 55916 126028 55972
rect 173012 55916 187852 55972
rect 187908 55916 189084 55972
rect 189140 55916 189150 55972
rect 202962 55916 202972 55972
rect 203028 55916 203756 55972
rect 203812 55916 205772 55972
rect 205828 55916 205838 55972
rect 264562 55916 264572 55972
rect 264628 55916 266364 55972
rect 266420 55916 266430 55972
rect 267092 55916 277228 55972
rect 277284 55916 277294 55972
rect 279682 55916 279692 55972
rect 279748 55916 281820 55972
rect 281876 55916 281886 55972
rect 125972 55860 126028 55916
rect 267092 55860 267148 55916
rect 125972 55804 183372 55860
rect 183428 55804 183438 55860
rect 209122 55804 209132 55860
rect 209188 55804 267148 55860
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 96626 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96910 55692
rect 127346 55636 127356 55692
rect 127412 55636 127460 55692
rect 127516 55636 127564 55692
rect 127620 55636 127630 55692
rect 158066 55636 158076 55692
rect 158132 55636 158180 55692
rect 158236 55636 158284 55692
rect 158340 55636 158350 55692
rect 188786 55636 188796 55692
rect 188852 55636 188900 55692
rect 188956 55636 189004 55692
rect 189060 55636 189070 55692
rect 219506 55636 219516 55692
rect 219572 55636 219620 55692
rect 219676 55636 219724 55692
rect 219780 55636 219790 55692
rect 250226 55636 250236 55692
rect 250292 55636 250340 55692
rect 250396 55636 250444 55692
rect 250500 55636 250510 55692
rect 280946 55636 280956 55692
rect 281012 55636 281060 55692
rect 281116 55636 281164 55692
rect 281220 55636 281230 55692
rect 61954 55468 61964 55524
rect 62020 55468 91644 55524
rect 91700 55468 91710 55524
rect 98802 55356 98812 55412
rect 98868 55356 100044 55412
rect 100100 55356 100110 55412
rect 141250 55356 141260 55412
rect 141316 55356 142604 55412
rect 142660 55356 142670 55412
rect 153906 55356 153916 55412
rect 153972 55356 156268 55412
rect 156324 55356 156716 55412
rect 156772 55356 161868 55412
rect 161924 55356 162428 55412
rect 162484 55356 162494 55412
rect 182354 55356 182364 55412
rect 182420 55356 186172 55412
rect 186228 55356 186238 55412
rect 186386 55356 186396 55412
rect 186452 55356 188300 55412
rect 188356 55356 188366 55412
rect 132962 55244 132972 55300
rect 133028 55244 135100 55300
rect 135156 55244 138348 55300
rect 138404 55244 140476 55300
rect 140532 55244 143836 55300
rect 143892 55244 147868 55300
rect 147924 55244 147934 55300
rect 169698 55244 169708 55300
rect 169764 55244 170380 55300
rect 170436 55244 174972 55300
rect 175028 55244 175532 55300
rect 175588 55244 179452 55300
rect 179508 55244 179518 55300
rect 110338 55132 110348 55188
rect 110404 55132 186956 55188
rect 187012 55132 187516 55188
rect 187572 55132 187582 55188
rect 152674 55020 152684 55076
rect 152740 55020 153244 55076
rect 153300 55020 166236 55076
rect 166292 55020 166302 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 81266 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81550 54908
rect 111986 54852 111996 54908
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 112260 54852 112270 54908
rect 142706 54852 142716 54908
rect 142772 54852 142820 54908
rect 142876 54852 142924 54908
rect 142980 54852 142990 54908
rect 173426 54852 173436 54908
rect 173492 54852 173540 54908
rect 173596 54852 173644 54908
rect 173700 54852 173710 54908
rect 204146 54852 204156 54908
rect 204212 54852 204260 54908
rect 204316 54852 204364 54908
rect 204420 54852 204430 54908
rect 234866 54852 234876 54908
rect 234932 54852 234980 54908
rect 235036 54852 235084 54908
rect 235140 54852 235150 54908
rect 265586 54852 265596 54908
rect 265652 54852 265700 54908
rect 265756 54852 265804 54908
rect 265860 54852 265870 54908
rect 296306 54852 296316 54908
rect 296372 54852 296420 54908
rect 296476 54852 296524 54908
rect 296580 54852 296590 54908
rect 148082 54684 148092 54740
rect 148148 54684 148652 54740
rect 148708 54684 150108 54740
rect 150164 54684 153916 54740
rect 153972 54684 153982 54740
rect 162306 54684 162316 54740
rect 162372 54684 163212 54740
rect 163268 54684 163278 54740
rect 167906 54684 167916 54740
rect 167972 54684 168924 54740
rect 168980 54684 168990 54740
rect 172722 54684 172732 54740
rect 172788 54684 174300 54740
rect 174356 54684 174366 54740
rect 220658 54572 220668 54628
rect 220724 54572 239260 54628
rect 239316 54572 239326 54628
rect 190418 54460 190428 54516
rect 190484 54460 191436 54516
rect 191492 54460 194572 54516
rect 194628 54460 194638 54516
rect 130274 54348 130284 54404
rect 130340 54348 131740 54404
rect 131796 54348 131806 54404
rect 145954 54348 145964 54404
rect 146020 54348 147420 54404
rect 147476 54348 147486 54404
rect 151554 54348 151564 54404
rect 151620 54348 153132 54404
rect 153188 54348 153198 54404
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 96626 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96910 54124
rect 127346 54068 127356 54124
rect 127412 54068 127460 54124
rect 127516 54068 127564 54124
rect 127620 54068 127630 54124
rect 158066 54068 158076 54124
rect 158132 54068 158180 54124
rect 158236 54068 158284 54124
rect 158340 54068 158350 54124
rect 188786 54068 188796 54124
rect 188852 54068 188900 54124
rect 188956 54068 189004 54124
rect 189060 54068 189070 54124
rect 219506 54068 219516 54124
rect 219572 54068 219620 54124
rect 219676 54068 219724 54124
rect 219780 54068 219790 54124
rect 250226 54068 250236 54124
rect 250292 54068 250340 54124
rect 250396 54068 250444 54124
rect 250500 54068 250510 54124
rect 280946 54068 280956 54124
rect 281012 54068 281060 54124
rect 281116 54068 281164 54124
rect 281220 54068 281230 54124
rect 225922 53900 225932 53956
rect 225988 53900 233996 53956
rect 234052 53900 234062 53956
rect 179442 53788 179452 53844
rect 179508 53788 180124 53844
rect 180180 53788 182140 53844
rect 182196 53788 182812 53844
rect 182868 53788 182878 53844
rect 193218 53788 193228 53844
rect 193284 53788 195804 53844
rect 195860 53788 195870 53844
rect 224242 53788 224252 53844
rect 224308 53788 228060 53844
rect 228116 53788 228126 53844
rect 186498 53676 186508 53732
rect 186564 53676 187964 53732
rect 188020 53676 189756 53732
rect 189812 53676 190428 53732
rect 190484 53676 190494 53732
rect 166226 53564 166236 53620
rect 166292 53564 167468 53620
rect 167524 53564 177660 53620
rect 177716 53564 178108 53620
rect 178164 53564 178174 53620
rect 183362 53452 183372 53508
rect 183428 53452 189420 53508
rect 189476 53452 191100 53508
rect 191156 53452 191166 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 81266 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81550 53340
rect 111986 53284 111996 53340
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 112260 53284 112270 53340
rect 142706 53284 142716 53340
rect 142772 53284 142820 53340
rect 142876 53284 142924 53340
rect 142980 53284 142990 53340
rect 173426 53284 173436 53340
rect 173492 53284 173540 53340
rect 173596 53284 173644 53340
rect 173700 53284 173710 53340
rect 204146 53284 204156 53340
rect 204212 53284 204260 53340
rect 204316 53284 204364 53340
rect 204420 53284 204430 53340
rect 234866 53284 234876 53340
rect 234932 53284 234980 53340
rect 235036 53284 235084 53340
rect 235140 53284 235150 53340
rect 265586 53284 265596 53340
rect 265652 53284 265700 53340
rect 265756 53284 265804 53340
rect 265860 53284 265870 53340
rect 296306 53284 296316 53340
rect 296372 53284 296420 53340
rect 296476 53284 296524 53340
rect 296580 53284 296590 53340
rect 182466 53116 182476 53172
rect 182532 53116 185836 53172
rect 185892 53116 186508 53172
rect 186564 53116 186574 53172
rect 127810 52780 127820 52836
rect 127876 52780 181468 52836
rect 181524 52780 183260 52836
rect 183316 52780 183326 52836
rect 186162 52780 186172 52836
rect 186228 52780 187180 52836
rect 187236 52780 187246 52836
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 96626 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96910 52556
rect 127346 52500 127356 52556
rect 127412 52500 127460 52556
rect 127516 52500 127564 52556
rect 127620 52500 127630 52556
rect 158066 52500 158076 52556
rect 158132 52500 158180 52556
rect 158236 52500 158284 52556
rect 158340 52500 158350 52556
rect 188786 52500 188796 52556
rect 188852 52500 188900 52556
rect 188956 52500 189004 52556
rect 189060 52500 189070 52556
rect 219506 52500 219516 52556
rect 219572 52500 219620 52556
rect 219676 52500 219724 52556
rect 219780 52500 219790 52556
rect 250226 52500 250236 52556
rect 250292 52500 250340 52556
rect 250396 52500 250444 52556
rect 250500 52500 250510 52556
rect 280946 52500 280956 52556
rect 281012 52500 281060 52556
rect 281116 52500 281164 52556
rect 281220 52500 281230 52556
rect 173012 52220 186172 52276
rect 186228 52220 186238 52276
rect 173012 52164 173068 52220
rect 116498 52108 116508 52164
rect 116564 52108 173068 52164
rect 189298 52108 189308 52164
rect 189364 52108 190652 52164
rect 190708 52108 190718 52164
rect 7410 51996 7420 52052
rect 7476 51996 161980 52052
rect 162036 51996 162046 52052
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 81266 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81550 51772
rect 111986 51716 111996 51772
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 112260 51716 112270 51772
rect 142706 51716 142716 51772
rect 142772 51716 142820 51772
rect 142876 51716 142924 51772
rect 142980 51716 142990 51772
rect 173426 51716 173436 51772
rect 173492 51716 173540 51772
rect 173596 51716 173644 51772
rect 173700 51716 173710 51772
rect 204146 51716 204156 51772
rect 204212 51716 204260 51772
rect 204316 51716 204364 51772
rect 204420 51716 204430 51772
rect 234866 51716 234876 51772
rect 234932 51716 234980 51772
rect 235036 51716 235084 51772
rect 235140 51716 235150 51772
rect 265586 51716 265596 51772
rect 265652 51716 265700 51772
rect 265756 51716 265804 51772
rect 265860 51716 265870 51772
rect 296306 51716 296316 51772
rect 296372 51716 296420 51772
rect 296476 51716 296524 51772
rect 296580 51716 296590 51772
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 96626 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96910 50988
rect 127346 50932 127356 50988
rect 127412 50932 127460 50988
rect 127516 50932 127564 50988
rect 127620 50932 127630 50988
rect 158066 50932 158076 50988
rect 158132 50932 158180 50988
rect 158236 50932 158284 50988
rect 158340 50932 158350 50988
rect 188786 50932 188796 50988
rect 188852 50932 188900 50988
rect 188956 50932 189004 50988
rect 189060 50932 189070 50988
rect 219506 50932 219516 50988
rect 219572 50932 219620 50988
rect 219676 50932 219724 50988
rect 219780 50932 219790 50988
rect 250226 50932 250236 50988
rect 250292 50932 250340 50988
rect 250396 50932 250444 50988
rect 250500 50932 250510 50988
rect 280946 50932 280956 50988
rect 281012 50932 281060 50988
rect 281116 50932 281164 50988
rect 281220 50932 281230 50988
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 81266 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81550 50204
rect 111986 50148 111996 50204
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 112260 50148 112270 50204
rect 142706 50148 142716 50204
rect 142772 50148 142820 50204
rect 142876 50148 142924 50204
rect 142980 50148 142990 50204
rect 173426 50148 173436 50204
rect 173492 50148 173540 50204
rect 173596 50148 173644 50204
rect 173700 50148 173710 50204
rect 204146 50148 204156 50204
rect 204212 50148 204260 50204
rect 204316 50148 204364 50204
rect 204420 50148 204430 50204
rect 234866 50148 234876 50204
rect 234932 50148 234980 50204
rect 235036 50148 235084 50204
rect 235140 50148 235150 50204
rect 265586 50148 265596 50204
rect 265652 50148 265700 50204
rect 265756 50148 265804 50204
rect 265860 50148 265870 50204
rect 296306 50148 296316 50204
rect 296372 50148 296420 50204
rect 296476 50148 296524 50204
rect 296580 50148 296590 50204
rect 102498 49532 102508 49588
rect 102564 49532 187292 49588
rect 187348 49532 187358 49588
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 96626 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96910 49420
rect 127346 49364 127356 49420
rect 127412 49364 127460 49420
rect 127516 49364 127564 49420
rect 127620 49364 127630 49420
rect 158066 49364 158076 49420
rect 158132 49364 158180 49420
rect 158236 49364 158284 49420
rect 158340 49364 158350 49420
rect 188786 49364 188796 49420
rect 188852 49364 188900 49420
rect 188956 49364 189004 49420
rect 189060 49364 189070 49420
rect 219506 49364 219516 49420
rect 219572 49364 219620 49420
rect 219676 49364 219724 49420
rect 219780 49364 219790 49420
rect 250226 49364 250236 49420
rect 250292 49364 250340 49420
rect 250396 49364 250444 49420
rect 250500 49364 250510 49420
rect 280946 49364 280956 49420
rect 281012 49364 281060 49420
rect 281116 49364 281164 49420
rect 281220 49364 281230 49420
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 81266 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81550 48636
rect 111986 48580 111996 48636
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 112260 48580 112270 48636
rect 142706 48580 142716 48636
rect 142772 48580 142820 48636
rect 142876 48580 142924 48636
rect 142980 48580 142990 48636
rect 173426 48580 173436 48636
rect 173492 48580 173540 48636
rect 173596 48580 173644 48636
rect 173700 48580 173710 48636
rect 204146 48580 204156 48636
rect 204212 48580 204260 48636
rect 204316 48580 204364 48636
rect 204420 48580 204430 48636
rect 234866 48580 234876 48636
rect 234932 48580 234980 48636
rect 235036 48580 235084 48636
rect 235140 48580 235150 48636
rect 265586 48580 265596 48636
rect 265652 48580 265700 48636
rect 265756 48580 265804 48636
rect 265860 48580 265870 48636
rect 296306 48580 296316 48636
rect 296372 48580 296420 48636
rect 296476 48580 296524 48636
rect 296580 48580 296590 48636
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 96626 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96910 47852
rect 127346 47796 127356 47852
rect 127412 47796 127460 47852
rect 127516 47796 127564 47852
rect 127620 47796 127630 47852
rect 158066 47796 158076 47852
rect 158132 47796 158180 47852
rect 158236 47796 158284 47852
rect 158340 47796 158350 47852
rect 188786 47796 188796 47852
rect 188852 47796 188900 47852
rect 188956 47796 189004 47852
rect 189060 47796 189070 47852
rect 219506 47796 219516 47852
rect 219572 47796 219620 47852
rect 219676 47796 219724 47852
rect 219780 47796 219790 47852
rect 250226 47796 250236 47852
rect 250292 47796 250340 47852
rect 250396 47796 250444 47852
rect 250500 47796 250510 47852
rect 280946 47796 280956 47852
rect 281012 47796 281060 47852
rect 281116 47796 281164 47852
rect 281220 47796 281230 47852
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 81266 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81550 47068
rect 111986 47012 111996 47068
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 112260 47012 112270 47068
rect 142706 47012 142716 47068
rect 142772 47012 142820 47068
rect 142876 47012 142924 47068
rect 142980 47012 142990 47068
rect 173426 47012 173436 47068
rect 173492 47012 173540 47068
rect 173596 47012 173644 47068
rect 173700 47012 173710 47068
rect 204146 47012 204156 47068
rect 204212 47012 204260 47068
rect 204316 47012 204364 47068
rect 204420 47012 204430 47068
rect 234866 47012 234876 47068
rect 234932 47012 234980 47068
rect 235036 47012 235084 47068
rect 235140 47012 235150 47068
rect 265586 47012 265596 47068
rect 265652 47012 265700 47068
rect 265756 47012 265804 47068
rect 265860 47012 265870 47068
rect 296306 47012 296316 47068
rect 296372 47012 296420 47068
rect 296476 47012 296524 47068
rect 296580 47012 296590 47068
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 96626 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96910 46284
rect 127346 46228 127356 46284
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127620 46228 127630 46284
rect 158066 46228 158076 46284
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158340 46228 158350 46284
rect 188786 46228 188796 46284
rect 188852 46228 188900 46284
rect 188956 46228 189004 46284
rect 189060 46228 189070 46284
rect 219506 46228 219516 46284
rect 219572 46228 219620 46284
rect 219676 46228 219724 46284
rect 219780 46228 219790 46284
rect 250226 46228 250236 46284
rect 250292 46228 250340 46284
rect 250396 46228 250444 46284
rect 250500 46228 250510 46284
rect 280946 46228 280956 46284
rect 281012 46228 281060 46284
rect 281116 46228 281164 46284
rect 281220 46228 281230 46284
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 81266 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81550 45500
rect 111986 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112270 45500
rect 142706 45444 142716 45500
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142980 45444 142990 45500
rect 173426 45444 173436 45500
rect 173492 45444 173540 45500
rect 173596 45444 173644 45500
rect 173700 45444 173710 45500
rect 204146 45444 204156 45500
rect 204212 45444 204260 45500
rect 204316 45444 204364 45500
rect 204420 45444 204430 45500
rect 234866 45444 234876 45500
rect 234932 45444 234980 45500
rect 235036 45444 235084 45500
rect 235140 45444 235150 45500
rect 265586 45444 265596 45500
rect 265652 45444 265700 45500
rect 265756 45444 265804 45500
rect 265860 45444 265870 45500
rect 296306 45444 296316 45500
rect 296372 45444 296420 45500
rect 296476 45444 296524 45500
rect 296580 45444 296590 45500
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 96626 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96910 44716
rect 127346 44660 127356 44716
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127620 44660 127630 44716
rect 158066 44660 158076 44716
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158340 44660 158350 44716
rect 188786 44660 188796 44716
rect 188852 44660 188900 44716
rect 188956 44660 189004 44716
rect 189060 44660 189070 44716
rect 219506 44660 219516 44716
rect 219572 44660 219620 44716
rect 219676 44660 219724 44716
rect 219780 44660 219790 44716
rect 250226 44660 250236 44716
rect 250292 44660 250340 44716
rect 250396 44660 250444 44716
rect 250500 44660 250510 44716
rect 280946 44660 280956 44716
rect 281012 44660 281060 44716
rect 281116 44660 281164 44716
rect 281220 44660 281230 44716
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 81266 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81550 43932
rect 111986 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112270 43932
rect 142706 43876 142716 43932
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142980 43876 142990 43932
rect 173426 43876 173436 43932
rect 173492 43876 173540 43932
rect 173596 43876 173644 43932
rect 173700 43876 173710 43932
rect 204146 43876 204156 43932
rect 204212 43876 204260 43932
rect 204316 43876 204364 43932
rect 204420 43876 204430 43932
rect 234866 43876 234876 43932
rect 234932 43876 234980 43932
rect 235036 43876 235084 43932
rect 235140 43876 235150 43932
rect 265586 43876 265596 43932
rect 265652 43876 265700 43932
rect 265756 43876 265804 43932
rect 265860 43876 265870 43932
rect 296306 43876 296316 43932
rect 296372 43876 296420 43932
rect 296476 43876 296524 43932
rect 296580 43876 296590 43932
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 96626 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96910 43148
rect 127346 43092 127356 43148
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127620 43092 127630 43148
rect 158066 43092 158076 43148
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158340 43092 158350 43148
rect 188786 43092 188796 43148
rect 188852 43092 188900 43148
rect 188956 43092 189004 43148
rect 189060 43092 189070 43148
rect 219506 43092 219516 43148
rect 219572 43092 219620 43148
rect 219676 43092 219724 43148
rect 219780 43092 219790 43148
rect 250226 43092 250236 43148
rect 250292 43092 250340 43148
rect 250396 43092 250444 43148
rect 250500 43092 250510 43148
rect 280946 43092 280956 43148
rect 281012 43092 281060 43148
rect 281116 43092 281164 43148
rect 281220 43092 281230 43148
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 81266 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81550 42364
rect 111986 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112270 42364
rect 142706 42308 142716 42364
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142980 42308 142990 42364
rect 173426 42308 173436 42364
rect 173492 42308 173540 42364
rect 173596 42308 173644 42364
rect 173700 42308 173710 42364
rect 204146 42308 204156 42364
rect 204212 42308 204260 42364
rect 204316 42308 204364 42364
rect 204420 42308 204430 42364
rect 234866 42308 234876 42364
rect 234932 42308 234980 42364
rect 235036 42308 235084 42364
rect 235140 42308 235150 42364
rect 265586 42308 265596 42364
rect 265652 42308 265700 42364
rect 265756 42308 265804 42364
rect 265860 42308 265870 42364
rect 296306 42308 296316 42364
rect 296372 42308 296420 42364
rect 296476 42308 296524 42364
rect 296580 42308 296590 42364
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 96626 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96910 41580
rect 127346 41524 127356 41580
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127620 41524 127630 41580
rect 158066 41524 158076 41580
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158340 41524 158350 41580
rect 188786 41524 188796 41580
rect 188852 41524 188900 41580
rect 188956 41524 189004 41580
rect 189060 41524 189070 41580
rect 219506 41524 219516 41580
rect 219572 41524 219620 41580
rect 219676 41524 219724 41580
rect 219780 41524 219790 41580
rect 250226 41524 250236 41580
rect 250292 41524 250340 41580
rect 250396 41524 250444 41580
rect 250500 41524 250510 41580
rect 280946 41524 280956 41580
rect 281012 41524 281060 41580
rect 281116 41524 281164 41580
rect 281220 41524 281230 41580
rect 54338 41132 54348 41188
rect 54404 41132 145180 41188
rect 145236 41132 145246 41188
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 81266 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81550 40796
rect 111986 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112270 40796
rect 142706 40740 142716 40796
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142980 40740 142990 40796
rect 173426 40740 173436 40796
rect 173492 40740 173540 40796
rect 173596 40740 173644 40796
rect 173700 40740 173710 40796
rect 204146 40740 204156 40796
rect 204212 40740 204260 40796
rect 204316 40740 204364 40796
rect 204420 40740 204430 40796
rect 234866 40740 234876 40796
rect 234932 40740 234980 40796
rect 235036 40740 235084 40796
rect 235140 40740 235150 40796
rect 265586 40740 265596 40796
rect 265652 40740 265700 40796
rect 265756 40740 265804 40796
rect 265860 40740 265870 40796
rect 296306 40740 296316 40796
rect 296372 40740 296420 40796
rect 296476 40740 296524 40796
rect 296580 40740 296590 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 96626 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96910 40012
rect 127346 39956 127356 40012
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127620 39956 127630 40012
rect 158066 39956 158076 40012
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158340 39956 158350 40012
rect 188786 39956 188796 40012
rect 188852 39956 188900 40012
rect 188956 39956 189004 40012
rect 189060 39956 189070 40012
rect 219506 39956 219516 40012
rect 219572 39956 219620 40012
rect 219676 39956 219724 40012
rect 219780 39956 219790 40012
rect 250226 39956 250236 40012
rect 250292 39956 250340 40012
rect 250396 39956 250444 40012
rect 250500 39956 250510 40012
rect 280946 39956 280956 40012
rect 281012 39956 281060 40012
rect 281116 39956 281164 40012
rect 281220 39956 281230 40012
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 81266 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81550 39228
rect 111986 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112270 39228
rect 142706 39172 142716 39228
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142980 39172 142990 39228
rect 173426 39172 173436 39228
rect 173492 39172 173540 39228
rect 173596 39172 173644 39228
rect 173700 39172 173710 39228
rect 204146 39172 204156 39228
rect 204212 39172 204260 39228
rect 204316 39172 204364 39228
rect 204420 39172 204430 39228
rect 234866 39172 234876 39228
rect 234932 39172 234980 39228
rect 235036 39172 235084 39228
rect 235140 39172 235150 39228
rect 265586 39172 265596 39228
rect 265652 39172 265700 39228
rect 265756 39172 265804 39228
rect 265860 39172 265870 39228
rect 296306 39172 296316 39228
rect 296372 39172 296420 39228
rect 296476 39172 296524 39228
rect 296580 39172 296590 39228
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 96626 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96910 38444
rect 127346 38388 127356 38444
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127620 38388 127630 38444
rect 158066 38388 158076 38444
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158340 38388 158350 38444
rect 188786 38388 188796 38444
rect 188852 38388 188900 38444
rect 188956 38388 189004 38444
rect 189060 38388 189070 38444
rect 219506 38388 219516 38444
rect 219572 38388 219620 38444
rect 219676 38388 219724 38444
rect 219780 38388 219790 38444
rect 250226 38388 250236 38444
rect 250292 38388 250340 38444
rect 250396 38388 250444 38444
rect 250500 38388 250510 38444
rect 280946 38388 280956 38444
rect 281012 38388 281060 38444
rect 281116 38388 281164 38444
rect 281220 38388 281230 38444
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 81266 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81550 37660
rect 111986 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112270 37660
rect 142706 37604 142716 37660
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142980 37604 142990 37660
rect 173426 37604 173436 37660
rect 173492 37604 173540 37660
rect 173596 37604 173644 37660
rect 173700 37604 173710 37660
rect 204146 37604 204156 37660
rect 204212 37604 204260 37660
rect 204316 37604 204364 37660
rect 204420 37604 204430 37660
rect 234866 37604 234876 37660
rect 234932 37604 234980 37660
rect 235036 37604 235084 37660
rect 235140 37604 235150 37660
rect 265586 37604 265596 37660
rect 265652 37604 265700 37660
rect 265756 37604 265804 37660
rect 265860 37604 265870 37660
rect 296306 37604 296316 37660
rect 296372 37604 296420 37660
rect 296476 37604 296524 37660
rect 296580 37604 296590 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 96626 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96910 36876
rect 127346 36820 127356 36876
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127620 36820 127630 36876
rect 158066 36820 158076 36876
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158340 36820 158350 36876
rect 188786 36820 188796 36876
rect 188852 36820 188900 36876
rect 188956 36820 189004 36876
rect 189060 36820 189070 36876
rect 219506 36820 219516 36876
rect 219572 36820 219620 36876
rect 219676 36820 219724 36876
rect 219780 36820 219790 36876
rect 250226 36820 250236 36876
rect 250292 36820 250340 36876
rect 250396 36820 250444 36876
rect 250500 36820 250510 36876
rect 280946 36820 280956 36876
rect 281012 36820 281060 36876
rect 281116 36820 281164 36876
rect 281220 36820 281230 36876
rect 68226 36204 68236 36260
rect 68292 36204 161532 36260
rect 161588 36204 161598 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 81266 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81550 36092
rect 111986 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112270 36092
rect 142706 36036 142716 36092
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142980 36036 142990 36092
rect 173426 36036 173436 36092
rect 173492 36036 173540 36092
rect 173596 36036 173644 36092
rect 173700 36036 173710 36092
rect 204146 36036 204156 36092
rect 204212 36036 204260 36092
rect 204316 36036 204364 36092
rect 204420 36036 204430 36092
rect 234866 36036 234876 36092
rect 234932 36036 234980 36092
rect 235036 36036 235084 36092
rect 235140 36036 235150 36092
rect 265586 36036 265596 36092
rect 265652 36036 265700 36092
rect 265756 36036 265804 36092
rect 265860 36036 265870 36092
rect 296306 36036 296316 36092
rect 296372 36036 296420 36092
rect 296476 36036 296524 36092
rect 296580 36036 296590 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 96626 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96910 35308
rect 127346 35252 127356 35308
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127620 35252 127630 35308
rect 158066 35252 158076 35308
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158340 35252 158350 35308
rect 188786 35252 188796 35308
rect 188852 35252 188900 35308
rect 188956 35252 189004 35308
rect 189060 35252 189070 35308
rect 219506 35252 219516 35308
rect 219572 35252 219620 35308
rect 219676 35252 219724 35308
rect 219780 35252 219790 35308
rect 250226 35252 250236 35308
rect 250292 35252 250340 35308
rect 250396 35252 250444 35308
rect 250500 35252 250510 35308
rect 280946 35252 280956 35308
rect 281012 35252 281060 35308
rect 281116 35252 281164 35308
rect 281220 35252 281230 35308
rect 69570 34636 69580 34692
rect 69636 34636 167132 34692
rect 167188 34636 167198 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 81266 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81550 34524
rect 111986 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112270 34524
rect 142706 34468 142716 34524
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142980 34468 142990 34524
rect 173426 34468 173436 34524
rect 173492 34468 173540 34524
rect 173596 34468 173644 34524
rect 173700 34468 173710 34524
rect 204146 34468 204156 34524
rect 204212 34468 204260 34524
rect 204316 34468 204364 34524
rect 204420 34468 204430 34524
rect 234866 34468 234876 34524
rect 234932 34468 234980 34524
rect 235036 34468 235084 34524
rect 235140 34468 235150 34524
rect 265586 34468 265596 34524
rect 265652 34468 265700 34524
rect 265756 34468 265804 34524
rect 265860 34468 265870 34524
rect 296306 34468 296316 34524
rect 296372 34468 296420 34524
rect 296476 34468 296524 34524
rect 296580 34468 296590 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 96626 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96910 33740
rect 127346 33684 127356 33740
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127620 33684 127630 33740
rect 158066 33684 158076 33740
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158340 33684 158350 33740
rect 188786 33684 188796 33740
rect 188852 33684 188900 33740
rect 188956 33684 189004 33740
rect 189060 33684 189070 33740
rect 219506 33684 219516 33740
rect 219572 33684 219620 33740
rect 219676 33684 219724 33740
rect 219780 33684 219790 33740
rect 250226 33684 250236 33740
rect 250292 33684 250340 33740
rect 250396 33684 250444 33740
rect 250500 33684 250510 33740
rect 280946 33684 280956 33740
rect 281012 33684 281060 33740
rect 281116 33684 281164 33740
rect 281220 33684 281230 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 81266 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81550 32956
rect 111986 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112270 32956
rect 142706 32900 142716 32956
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142980 32900 142990 32956
rect 173426 32900 173436 32956
rect 173492 32900 173540 32956
rect 173596 32900 173644 32956
rect 173700 32900 173710 32956
rect 204146 32900 204156 32956
rect 204212 32900 204260 32956
rect 204316 32900 204364 32956
rect 204420 32900 204430 32956
rect 234866 32900 234876 32956
rect 234932 32900 234980 32956
rect 235036 32900 235084 32956
rect 235140 32900 235150 32956
rect 265586 32900 265596 32956
rect 265652 32900 265700 32956
rect 265756 32900 265804 32956
rect 265860 32900 265870 32956
rect 296306 32900 296316 32956
rect 296372 32900 296420 32956
rect 296476 32900 296524 32956
rect 296580 32900 296590 32956
rect 60946 32732 60956 32788
rect 61012 32732 156380 32788
rect 156436 32732 156446 32788
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 96626 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96910 32172
rect 127346 32116 127356 32172
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127620 32116 127630 32172
rect 158066 32116 158076 32172
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158340 32116 158350 32172
rect 188786 32116 188796 32172
rect 188852 32116 188900 32172
rect 188956 32116 189004 32172
rect 189060 32116 189070 32172
rect 219506 32116 219516 32172
rect 219572 32116 219620 32172
rect 219676 32116 219724 32172
rect 219780 32116 219790 32172
rect 250226 32116 250236 32172
rect 250292 32116 250340 32172
rect 250396 32116 250444 32172
rect 250500 32116 250510 32172
rect 280946 32116 280956 32172
rect 281012 32116 281060 32172
rect 281116 32116 281164 32172
rect 281220 32116 281230 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 81266 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81550 31388
rect 111986 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112270 31388
rect 142706 31332 142716 31388
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142980 31332 142990 31388
rect 173426 31332 173436 31388
rect 173492 31332 173540 31388
rect 173596 31332 173644 31388
rect 173700 31332 173710 31388
rect 204146 31332 204156 31388
rect 204212 31332 204260 31388
rect 204316 31332 204364 31388
rect 204420 31332 204430 31388
rect 234866 31332 234876 31388
rect 234932 31332 234980 31388
rect 235036 31332 235084 31388
rect 235140 31332 235150 31388
rect 265586 31332 265596 31388
rect 265652 31332 265700 31388
rect 265756 31332 265804 31388
rect 265860 31332 265870 31388
rect 296306 31332 296316 31388
rect 296372 31332 296420 31388
rect 296476 31332 296524 31388
rect 296580 31332 296590 31388
rect 57250 31052 57260 31108
rect 57316 31052 150780 31108
rect 150836 31052 150846 31108
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 96626 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96910 30604
rect 127346 30548 127356 30604
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127620 30548 127630 30604
rect 158066 30548 158076 30604
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158340 30548 158350 30604
rect 188786 30548 188796 30604
rect 188852 30548 188900 30604
rect 188956 30548 189004 30604
rect 189060 30548 189070 30604
rect 219506 30548 219516 30604
rect 219572 30548 219620 30604
rect 219676 30548 219724 30604
rect 219780 30548 219790 30604
rect 250226 30548 250236 30604
rect 250292 30548 250340 30604
rect 250396 30548 250444 30604
rect 250500 30548 250510 30604
rect 280946 30548 280956 30604
rect 281012 30548 281060 30604
rect 281116 30548 281164 30604
rect 281220 30548 281230 30604
rect 205762 30268 205772 30324
rect 205828 30268 210028 30324
rect 210084 30268 210094 30324
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 81266 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81550 29820
rect 111986 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112270 29820
rect 142706 29764 142716 29820
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142980 29764 142990 29820
rect 173426 29764 173436 29820
rect 173492 29764 173540 29820
rect 173596 29764 173644 29820
rect 173700 29764 173710 29820
rect 204146 29764 204156 29820
rect 204212 29764 204260 29820
rect 204316 29764 204364 29820
rect 204420 29764 204430 29820
rect 234866 29764 234876 29820
rect 234932 29764 234980 29820
rect 235036 29764 235084 29820
rect 235140 29764 235150 29820
rect 265586 29764 265596 29820
rect 265652 29764 265700 29820
rect 265756 29764 265804 29820
rect 265860 29764 265870 29820
rect 296306 29764 296316 29820
rect 296372 29764 296420 29820
rect 296476 29764 296524 29820
rect 296580 29764 296590 29820
rect 59602 29372 59612 29428
rect 59668 29372 140252 29428
rect 140308 29372 140318 29428
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 96626 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96910 29036
rect 127346 28980 127356 29036
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127620 28980 127630 29036
rect 158066 28980 158076 29036
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158340 28980 158350 29036
rect 188786 28980 188796 29036
rect 188852 28980 188900 29036
rect 188956 28980 189004 29036
rect 189060 28980 189070 29036
rect 219506 28980 219516 29036
rect 219572 28980 219620 29036
rect 219676 28980 219724 29036
rect 219780 28980 219790 29036
rect 250226 28980 250236 29036
rect 250292 28980 250340 29036
rect 250396 28980 250444 29036
rect 250500 28980 250510 29036
rect 280946 28980 280956 29036
rect 281012 28980 281060 29036
rect 281116 28980 281164 29036
rect 281220 28980 281230 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 81266 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81550 28252
rect 111986 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112270 28252
rect 142706 28196 142716 28252
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142980 28196 142990 28252
rect 173426 28196 173436 28252
rect 173492 28196 173540 28252
rect 173596 28196 173644 28252
rect 173700 28196 173710 28252
rect 204146 28196 204156 28252
rect 204212 28196 204260 28252
rect 204316 28196 204364 28252
rect 204420 28196 204430 28252
rect 234866 28196 234876 28252
rect 234932 28196 234980 28252
rect 235036 28196 235084 28252
rect 235140 28196 235150 28252
rect 265586 28196 265596 28252
rect 265652 28196 265700 28252
rect 265756 28196 265804 28252
rect 265860 28196 265870 28252
rect 296306 28196 296316 28252
rect 296372 28196 296420 28252
rect 296476 28196 296524 28252
rect 296580 28196 296590 28252
rect 202290 27692 202300 27748
rect 202356 27692 288092 27748
rect 288148 27692 288158 27748
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 96626 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96910 27468
rect 127346 27412 127356 27468
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127620 27412 127630 27468
rect 158066 27412 158076 27468
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158340 27412 158350 27468
rect 188786 27412 188796 27468
rect 188852 27412 188900 27468
rect 188956 27412 189004 27468
rect 189060 27412 189070 27468
rect 219506 27412 219516 27468
rect 219572 27412 219620 27468
rect 219676 27412 219724 27468
rect 219780 27412 219790 27468
rect 250226 27412 250236 27468
rect 250292 27412 250340 27468
rect 250396 27412 250444 27468
rect 250500 27412 250510 27468
rect 280946 27412 280956 27468
rect 281012 27412 281060 27468
rect 281116 27412 281164 27468
rect 281220 27412 281230 27468
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 81266 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81550 26684
rect 111986 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112270 26684
rect 142706 26628 142716 26684
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142980 26628 142990 26684
rect 173426 26628 173436 26684
rect 173492 26628 173540 26684
rect 173596 26628 173644 26684
rect 173700 26628 173710 26684
rect 204146 26628 204156 26684
rect 204212 26628 204260 26684
rect 204316 26628 204364 26684
rect 204420 26628 204430 26684
rect 234866 26628 234876 26684
rect 234932 26628 234980 26684
rect 235036 26628 235084 26684
rect 235140 26628 235150 26684
rect 265586 26628 265596 26684
rect 265652 26628 265700 26684
rect 265756 26628 265804 26684
rect 265860 26628 265870 26684
rect 296306 26628 296316 26684
rect 296372 26628 296420 26684
rect 296476 26628 296524 26684
rect 296580 26628 296590 26684
rect 47618 26012 47628 26068
rect 47684 26012 134876 26068
rect 134932 26012 134942 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 96626 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96910 25900
rect 127346 25844 127356 25900
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127620 25844 127630 25900
rect 158066 25844 158076 25900
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158340 25844 158350 25900
rect 188786 25844 188796 25900
rect 188852 25844 188900 25900
rect 188956 25844 189004 25900
rect 189060 25844 189070 25900
rect 219506 25844 219516 25900
rect 219572 25844 219620 25900
rect 219676 25844 219724 25900
rect 219780 25844 219790 25900
rect 250226 25844 250236 25900
rect 250292 25844 250340 25900
rect 250396 25844 250444 25900
rect 250500 25844 250510 25900
rect 280946 25844 280956 25900
rect 281012 25844 281060 25900
rect 281116 25844 281164 25900
rect 281220 25844 281230 25900
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 81266 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81550 25116
rect 111986 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112270 25116
rect 142706 25060 142716 25116
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142980 25060 142990 25116
rect 173426 25060 173436 25116
rect 173492 25060 173540 25116
rect 173596 25060 173644 25116
rect 173700 25060 173710 25116
rect 204146 25060 204156 25116
rect 204212 25060 204260 25116
rect 204316 25060 204364 25116
rect 204420 25060 204430 25116
rect 234866 25060 234876 25116
rect 234932 25060 234980 25116
rect 235036 25060 235084 25116
rect 235140 25060 235150 25116
rect 265586 25060 265596 25116
rect 265652 25060 265700 25116
rect 265756 25060 265804 25116
rect 265860 25060 265870 25116
rect 296306 25060 296316 25116
rect 296372 25060 296420 25116
rect 296476 25060 296524 25116
rect 296580 25060 296590 25116
rect 43810 24444 43820 24500
rect 43876 24444 129388 24500
rect 129444 24444 129454 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 96626 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96910 24332
rect 127346 24276 127356 24332
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127620 24276 127630 24332
rect 158066 24276 158076 24332
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158340 24276 158350 24332
rect 188786 24276 188796 24332
rect 188852 24276 188900 24332
rect 188956 24276 189004 24332
rect 189060 24276 189070 24332
rect 219506 24276 219516 24332
rect 219572 24276 219620 24332
rect 219676 24276 219724 24332
rect 219780 24276 219790 24332
rect 250226 24276 250236 24332
rect 250292 24276 250340 24332
rect 250396 24276 250444 24332
rect 250500 24276 250510 24332
rect 280946 24276 280956 24332
rect 281012 24276 281060 24332
rect 281116 24276 281164 24332
rect 281220 24276 281230 24332
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 81266 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81550 23548
rect 111986 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112270 23548
rect 142706 23492 142716 23548
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142980 23492 142990 23548
rect 173426 23492 173436 23548
rect 173492 23492 173540 23548
rect 173596 23492 173644 23548
rect 173700 23492 173710 23548
rect 204146 23492 204156 23548
rect 204212 23492 204260 23548
rect 204316 23492 204364 23548
rect 204420 23492 204430 23548
rect 234866 23492 234876 23548
rect 234932 23492 234980 23548
rect 235036 23492 235084 23548
rect 235140 23492 235150 23548
rect 265586 23492 265596 23548
rect 265652 23492 265700 23548
rect 265756 23492 265804 23548
rect 265860 23492 265870 23548
rect 296306 23492 296316 23548
rect 296372 23492 296420 23548
rect 296476 23492 296524 23548
rect 296580 23492 296590 23548
rect 52882 22876 52892 22932
rect 52948 22876 88732 22932
rect 88788 22876 88798 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 96626 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96910 22764
rect 127346 22708 127356 22764
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127620 22708 127630 22764
rect 158066 22708 158076 22764
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158340 22708 158350 22764
rect 188786 22708 188796 22764
rect 188852 22708 188900 22764
rect 188956 22708 189004 22764
rect 189060 22708 189070 22764
rect 219506 22708 219516 22764
rect 219572 22708 219620 22764
rect 219676 22708 219724 22764
rect 219780 22708 219790 22764
rect 250226 22708 250236 22764
rect 250292 22708 250340 22764
rect 250396 22708 250444 22764
rect 250500 22708 250510 22764
rect 280946 22708 280956 22764
rect 281012 22708 281060 22764
rect 281116 22708 281164 22764
rect 281220 22708 281230 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 81266 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81550 21980
rect 111986 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112270 21980
rect 142706 21924 142716 21980
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142980 21924 142990 21980
rect 173426 21924 173436 21980
rect 173492 21924 173540 21980
rect 173596 21924 173644 21980
rect 173700 21924 173710 21980
rect 204146 21924 204156 21980
rect 204212 21924 204260 21980
rect 204316 21924 204364 21980
rect 204420 21924 204430 21980
rect 234866 21924 234876 21980
rect 234932 21924 234980 21980
rect 235036 21924 235084 21980
rect 235140 21924 235150 21980
rect 265586 21924 265596 21980
rect 265652 21924 265700 21980
rect 265756 21924 265804 21980
rect 265860 21924 265870 21980
rect 296306 21924 296316 21980
rect 296372 21924 296420 21980
rect 296476 21924 296524 21980
rect 296580 21924 296590 21980
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 96626 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96910 21196
rect 127346 21140 127356 21196
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127620 21140 127630 21196
rect 158066 21140 158076 21196
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158340 21140 158350 21196
rect 188786 21140 188796 21196
rect 188852 21140 188900 21196
rect 188956 21140 189004 21196
rect 189060 21140 189070 21196
rect 219506 21140 219516 21196
rect 219572 21140 219620 21196
rect 219676 21140 219724 21196
rect 219780 21140 219790 21196
rect 250226 21140 250236 21196
rect 250292 21140 250340 21196
rect 250396 21140 250444 21196
rect 250500 21140 250510 21196
rect 280946 21140 280956 21196
rect 281012 21140 281060 21196
rect 281116 21140 281164 21196
rect 281220 21140 281230 21196
rect 45826 20972 45836 21028
rect 45892 20972 85036 21028
rect 85092 20972 85102 21028
rect 92418 20972 92428 21028
rect 92484 20972 178892 21028
rect 178948 20972 178958 21028
rect 207890 20972 207900 21028
rect 207956 20972 293356 21028
rect 293412 20972 293422 21028
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 81266 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81550 20412
rect 111986 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112270 20412
rect 142706 20356 142716 20412
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142980 20356 142990 20412
rect 173426 20356 173436 20412
rect 173492 20356 173540 20412
rect 173596 20356 173644 20412
rect 173700 20356 173710 20412
rect 204146 20356 204156 20412
rect 204212 20356 204260 20412
rect 204316 20356 204364 20412
rect 204420 20356 204430 20412
rect 234866 20356 234876 20412
rect 234932 20356 234980 20412
rect 235036 20356 235084 20412
rect 235140 20356 235150 20412
rect 265586 20356 265596 20412
rect 265652 20356 265700 20412
rect 265756 20356 265804 20412
rect 265860 20356 265870 20412
rect 296306 20356 296316 20412
rect 296372 20356 296420 20412
rect 296476 20356 296524 20412
rect 296580 20356 296590 20412
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 96626 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96910 19628
rect 127346 19572 127356 19628
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127620 19572 127630 19628
rect 158066 19572 158076 19628
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158340 19572 158350 19628
rect 188786 19572 188796 19628
rect 188852 19572 188900 19628
rect 188956 19572 189004 19628
rect 189060 19572 189070 19628
rect 219506 19572 219516 19628
rect 219572 19572 219620 19628
rect 219676 19572 219724 19628
rect 219780 19572 219790 19628
rect 250226 19572 250236 19628
rect 250292 19572 250340 19628
rect 250396 19572 250444 19628
rect 250500 19572 250510 19628
rect 280946 19572 280956 19628
rect 281012 19572 281060 19628
rect 281116 19572 281164 19628
rect 281220 19572 281230 19628
rect 35074 19292 35084 19348
rect 35140 19292 78652 19348
rect 78708 19292 78718 19348
rect 185378 19292 185388 19348
rect 185444 19292 198492 19348
rect 198548 19292 198558 19348
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 81266 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81550 18844
rect 111986 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112270 18844
rect 142706 18788 142716 18844
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142980 18788 142990 18844
rect 173426 18788 173436 18844
rect 173492 18788 173540 18844
rect 173596 18788 173644 18844
rect 173700 18788 173710 18844
rect 204146 18788 204156 18844
rect 204212 18788 204260 18844
rect 204316 18788 204364 18844
rect 204420 18788 204430 18844
rect 234866 18788 234876 18844
rect 234932 18788 234980 18844
rect 235036 18788 235084 18844
rect 235140 18788 235150 18844
rect 265586 18788 265596 18844
rect 265652 18788 265700 18844
rect 265756 18788 265804 18844
rect 265860 18788 265870 18844
rect 296306 18788 296316 18844
rect 296372 18788 296420 18844
rect 296476 18788 296524 18844
rect 296580 18788 296590 18844
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 96626 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96910 18060
rect 127346 18004 127356 18060
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127620 18004 127630 18060
rect 158066 18004 158076 18060
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158340 18004 158350 18060
rect 188786 18004 188796 18060
rect 188852 18004 188900 18060
rect 188956 18004 189004 18060
rect 189060 18004 189070 18060
rect 219506 18004 219516 18060
rect 219572 18004 219620 18060
rect 219676 18004 219724 18060
rect 219780 18004 219790 18060
rect 250226 18004 250236 18060
rect 250292 18004 250340 18060
rect 250396 18004 250444 18060
rect 250500 18004 250510 18060
rect 280946 18004 280956 18060
rect 281012 18004 281060 18060
rect 281116 18004 281164 18060
rect 281220 18004 281230 18060
rect 83122 17612 83132 17668
rect 83188 17612 183372 17668
rect 183428 17612 183438 17668
rect 191314 17612 191324 17668
rect 191380 17612 206892 17668
rect 206948 17612 206958 17668
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 81266 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81550 17276
rect 111986 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112270 17276
rect 142706 17220 142716 17276
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142980 17220 142990 17276
rect 173426 17220 173436 17276
rect 173492 17220 173540 17276
rect 173596 17220 173644 17276
rect 173700 17220 173710 17276
rect 204146 17220 204156 17276
rect 204212 17220 204260 17276
rect 204316 17220 204364 17276
rect 204420 17220 204430 17276
rect 234866 17220 234876 17276
rect 234932 17220 234980 17276
rect 235036 17220 235084 17276
rect 235140 17220 235150 17276
rect 265586 17220 265596 17276
rect 265652 17220 265700 17276
rect 265756 17220 265804 17276
rect 265860 17220 265870 17276
rect 296306 17220 296316 17276
rect 296372 17220 296420 17276
rect 296476 17220 296524 17276
rect 296580 17220 296590 17276
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 96626 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96910 16492
rect 127346 16436 127356 16492
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127620 16436 127630 16492
rect 158066 16436 158076 16492
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158340 16436 158350 16492
rect 188786 16436 188796 16492
rect 188852 16436 188900 16492
rect 188956 16436 189004 16492
rect 189060 16436 189070 16492
rect 219506 16436 219516 16492
rect 219572 16436 219620 16492
rect 219676 16436 219724 16492
rect 219780 16436 219790 16492
rect 250226 16436 250236 16492
rect 250292 16436 250340 16492
rect 250396 16436 250444 16492
rect 250500 16436 250510 16492
rect 280946 16436 280956 16492
rect 281012 16436 281060 16492
rect 281116 16436 281164 16492
rect 281220 16436 281230 16492
rect 40450 15932 40460 15988
rect 40516 15932 83132 15988
rect 83188 15932 83198 15988
rect 107650 15932 107660 15988
rect 107716 15932 182252 15988
rect 182308 15932 182318 15988
rect 193218 15932 193228 15988
rect 193284 15932 264572 15988
rect 264628 15932 264638 15988
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 81266 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81550 15708
rect 111986 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112270 15708
rect 142706 15652 142716 15708
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142980 15652 142990 15708
rect 173426 15652 173436 15708
rect 173492 15652 173540 15708
rect 173596 15652 173644 15708
rect 173700 15652 173710 15708
rect 204146 15652 204156 15708
rect 204212 15652 204260 15708
rect 204316 15652 204364 15708
rect 204420 15652 204430 15708
rect 234866 15652 234876 15708
rect 234932 15652 234980 15708
rect 235036 15652 235084 15708
rect 235140 15652 235150 15708
rect 265586 15652 265596 15708
rect 265652 15652 265700 15708
rect 265756 15652 265804 15708
rect 265860 15652 265870 15708
rect 296306 15652 296316 15708
rect 296372 15652 296420 15708
rect 296476 15652 296524 15708
rect 296580 15652 296590 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 96626 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96910 14924
rect 127346 14868 127356 14924
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127620 14868 127630 14924
rect 158066 14868 158076 14924
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158340 14868 158350 14924
rect 188786 14868 188796 14924
rect 188852 14868 188900 14924
rect 188956 14868 189004 14924
rect 189060 14868 189070 14924
rect 219506 14868 219516 14924
rect 219572 14868 219620 14924
rect 219676 14868 219724 14924
rect 219780 14868 219790 14924
rect 250226 14868 250236 14924
rect 250292 14868 250340 14924
rect 250396 14868 250444 14924
rect 250500 14868 250510 14924
rect 280946 14868 280956 14924
rect 281012 14868 281060 14924
rect 281116 14868 281164 14924
rect 281220 14868 281230 14924
rect 75170 14252 75180 14308
rect 75236 14252 184828 14308
rect 184884 14252 184894 14308
rect 196690 14252 196700 14308
rect 196756 14252 256060 14308
rect 256116 14252 256126 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 81266 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81550 14140
rect 111986 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112270 14140
rect 142706 14084 142716 14140
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142980 14084 142990 14140
rect 173426 14084 173436 14140
rect 173492 14084 173540 14140
rect 173596 14084 173644 14140
rect 173700 14084 173710 14140
rect 204146 14084 204156 14140
rect 204212 14084 204260 14140
rect 204316 14084 204364 14140
rect 204420 14084 204430 14140
rect 234866 14084 234876 14140
rect 234932 14084 234980 14140
rect 235036 14084 235084 14140
rect 235140 14084 235150 14140
rect 265586 14084 265596 14140
rect 265652 14084 265700 14140
rect 265756 14084 265804 14140
rect 265860 14084 265870 14140
rect 296306 14084 296316 14140
rect 296372 14084 296420 14140
rect 296476 14084 296524 14140
rect 296580 14084 296590 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 96626 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96910 13356
rect 127346 13300 127356 13356
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127620 13300 127630 13356
rect 158066 13300 158076 13356
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158340 13300 158350 13356
rect 188786 13300 188796 13356
rect 188852 13300 188900 13356
rect 188956 13300 189004 13356
rect 189060 13300 189070 13356
rect 219506 13300 219516 13356
rect 219572 13300 219620 13356
rect 219676 13300 219724 13356
rect 219780 13300 219790 13356
rect 250226 13300 250236 13356
rect 250292 13300 250340 13356
rect 250396 13300 250444 13356
rect 250500 13300 250510 13356
rect 280946 13300 280956 13356
rect 281012 13300 281060 13356
rect 281116 13300 281164 13356
rect 281220 13300 281230 13356
rect 217410 12908 217420 12964
rect 217476 12908 250124 12964
rect 250180 12908 250190 12964
rect 208226 12796 208236 12852
rect 208292 12796 273196 12852
rect 273252 12796 273262 12852
rect 73042 12684 73052 12740
rect 73108 12684 185276 12740
rect 185332 12684 185342 12740
rect 203634 12684 203644 12740
rect 203700 12684 279692 12740
rect 279748 12684 279758 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 81266 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81550 12572
rect 111986 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112270 12572
rect 142706 12516 142716 12572
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142980 12516 142990 12572
rect 173426 12516 173436 12572
rect 173492 12516 173540 12572
rect 173596 12516 173644 12572
rect 173700 12516 173710 12572
rect 204146 12516 204156 12572
rect 204212 12516 204260 12572
rect 204316 12516 204364 12572
rect 204420 12516 204430 12572
rect 234866 12516 234876 12572
rect 234932 12516 234980 12572
rect 235036 12516 235084 12572
rect 235140 12516 235150 12572
rect 265586 12516 265596 12572
rect 265652 12516 265700 12572
rect 265756 12516 265804 12572
rect 265860 12516 265870 12572
rect 296306 12516 296316 12572
rect 296372 12516 296420 12572
rect 296476 12516 296524 12572
rect 296580 12516 296590 12572
rect 213388 11788 217308 11844
rect 217364 11788 217374 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 96626 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96910 11788
rect 127346 11732 127356 11788
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127620 11732 127630 11788
rect 158066 11732 158076 11788
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158340 11732 158350 11788
rect 188786 11732 188796 11788
rect 188852 11732 188900 11788
rect 188956 11732 189004 11788
rect 189060 11732 189070 11788
rect 213388 11732 213444 11788
rect 219506 11732 219516 11788
rect 219572 11732 219620 11788
rect 219676 11732 219724 11788
rect 219780 11732 219790 11788
rect 250226 11732 250236 11788
rect 250292 11732 250340 11788
rect 250396 11732 250444 11788
rect 250500 11732 250510 11788
rect 280946 11732 280956 11788
rect 281012 11732 281060 11788
rect 281116 11732 281164 11788
rect 281220 11732 281230 11788
rect 211922 11676 211932 11732
rect 211988 11676 213444 11732
rect 73378 11228 73388 11284
rect 73444 11228 171948 11284
rect 172004 11228 172014 11284
rect 221778 11228 221788 11284
rect 221844 11228 244748 11284
rect 244804 11228 244814 11284
rect 85698 11116 85708 11172
rect 85764 11116 192556 11172
rect 192612 11116 192622 11172
rect 195010 11116 195020 11172
rect 195076 11116 261772 11172
rect 261828 11116 261838 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 81266 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81550 11004
rect 111986 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112270 11004
rect 142706 10948 142716 11004
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142980 10948 142990 11004
rect 173426 10948 173436 11004
rect 173492 10948 173540 11004
rect 173596 10948 173644 11004
rect 173700 10948 173710 11004
rect 204146 10948 204156 11004
rect 204212 10948 204260 11004
rect 204316 10948 204364 11004
rect 204420 10948 204430 11004
rect 234866 10948 234876 11004
rect 234932 10948 234980 11004
rect 235036 10948 235084 11004
rect 235140 10948 235150 11004
rect 265586 10948 265596 11004
rect 265652 10948 265700 11004
rect 265756 10948 265804 11004
rect 265860 10948 265870 11004
rect 296306 10948 296316 11004
rect 296372 10948 296420 11004
rect 296476 10948 296524 11004
rect 296580 10948 296590 11004
rect 196532 10444 220780 10500
rect 220836 10444 220846 10500
rect 196532 10388 196588 10444
rect 196130 10332 196140 10388
rect 196196 10332 196588 10388
rect 213602 10332 213612 10388
rect 213668 10332 222684 10388
rect 222740 10332 222750 10388
rect 190642 10220 190652 10276
rect 190708 10220 199164 10276
rect 199220 10220 199230 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 96626 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96910 10220
rect 127346 10164 127356 10220
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127620 10164 127630 10220
rect 158066 10164 158076 10220
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158340 10164 158350 10220
rect 188786 10164 188796 10220
rect 188852 10164 188900 10220
rect 188956 10164 189004 10220
rect 189060 10164 189070 10220
rect 219506 10164 219516 10220
rect 219572 10164 219620 10220
rect 219676 10164 219724 10220
rect 219780 10164 219790 10220
rect 250226 10164 250236 10220
rect 250292 10164 250340 10220
rect 250396 10164 250444 10220
rect 250500 10164 250510 10220
rect 280946 10164 280956 10220
rect 281012 10164 281060 10220
rect 281116 10164 281164 10220
rect 281220 10164 281230 10220
rect 195794 10108 195804 10164
rect 195860 10108 199724 10164
rect 199780 10108 199790 10164
rect 196242 9996 196252 10052
rect 196308 9996 220556 10052
rect 220612 9996 220622 10052
rect 195458 9884 195468 9940
rect 195524 9884 270620 9940
rect 270676 9884 270686 9940
rect 196018 9772 196028 9828
rect 196084 9772 218316 9828
rect 218372 9772 218382 9828
rect 210690 9660 210700 9716
rect 210756 9660 211036 9716
rect 211092 9660 211102 9716
rect 218418 9660 218428 9716
rect 218484 9660 219548 9716
rect 219604 9660 221788 9716
rect 221844 9660 221854 9716
rect 199714 9548 199724 9604
rect 199780 9548 200956 9604
rect 201012 9548 201022 9604
rect 203074 9548 203084 9604
rect 203140 9548 212492 9604
rect 212548 9548 216748 9604
rect 216804 9548 217532 9604
rect 217588 9548 217598 9604
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 81266 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81550 9436
rect 111986 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112270 9436
rect 142706 9380 142716 9436
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142980 9380 142990 9436
rect 173426 9380 173436 9436
rect 173492 9380 173540 9436
rect 173596 9380 173644 9436
rect 173700 9380 173710 9436
rect 204146 9380 204156 9436
rect 204212 9380 204260 9436
rect 204316 9380 204364 9436
rect 204420 9380 204430 9436
rect 234866 9380 234876 9436
rect 234932 9380 234980 9436
rect 235036 9380 235084 9436
rect 235140 9380 235150 9436
rect 265586 9380 265596 9436
rect 265652 9380 265700 9436
rect 265756 9380 265804 9436
rect 265860 9380 265870 9436
rect 296306 9380 296316 9436
rect 296372 9380 296420 9436
rect 296476 9380 296524 9436
rect 296580 9380 296590 9436
rect 29698 9212 29708 9268
rect 29764 9212 74844 9268
rect 74900 9212 74910 9268
rect 99922 9212 99932 9268
rect 99988 9212 193564 9268
rect 193620 9212 193630 9268
rect 197586 9212 197596 9268
rect 197652 9212 202300 9268
rect 202356 9212 202366 9268
rect 217746 9212 217756 9268
rect 217812 9212 219100 9268
rect 219156 9212 219996 9268
rect 220052 9212 221228 9268
rect 221284 9212 221294 9268
rect 221890 9212 221900 9268
rect 221956 9212 222348 9268
rect 222404 9212 224252 9268
rect 224308 9212 224318 9268
rect 220332 9156 220388 9212
rect 119186 9100 119196 9156
rect 119252 9100 209916 9156
rect 209972 9100 209982 9156
rect 210690 9100 210700 9156
rect 210756 9100 211260 9156
rect 211316 9100 211708 9156
rect 211764 9100 213388 9156
rect 213444 9100 213454 9156
rect 220322 9100 220332 9156
rect 220388 9100 220398 9156
rect 187282 8988 187292 9044
rect 187348 8988 192668 9044
rect 192724 8988 192734 9044
rect 201282 8988 201292 9044
rect 201348 8988 203644 9044
rect 203700 8988 203710 9044
rect 207676 8988 213836 9044
rect 213892 8988 216524 9044
rect 216580 8988 218764 9044
rect 218820 8988 218830 9044
rect 207676 8932 207732 8988
rect 206322 8876 206332 8932
rect 206388 8876 207676 8932
rect 207732 8876 207742 8932
rect 208292 8876 209132 8932
rect 209188 8876 209198 8932
rect 208292 8820 208348 8876
rect 199042 8764 199052 8820
rect 199108 8764 199500 8820
rect 199556 8764 199566 8820
rect 203858 8764 203868 8820
rect 203924 8764 208348 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 96626 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96910 8652
rect 127346 8596 127356 8652
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127620 8596 127630 8652
rect 158066 8596 158076 8652
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158340 8596 158350 8652
rect 188786 8596 188796 8652
rect 188852 8596 188900 8652
rect 188956 8596 189004 8652
rect 189060 8596 189070 8652
rect 219506 8596 219516 8652
rect 219572 8596 219620 8652
rect 219676 8596 219724 8652
rect 219780 8596 219790 8652
rect 250226 8596 250236 8652
rect 250292 8596 250340 8652
rect 250396 8596 250444 8652
rect 250500 8596 250510 8652
rect 280946 8596 280956 8652
rect 281012 8596 281060 8652
rect 281116 8596 281164 8652
rect 281220 8596 281230 8652
rect 191090 8540 191100 8596
rect 191156 8540 215740 8596
rect 215796 8540 215806 8596
rect 203970 8428 203980 8484
rect 204036 8428 217308 8484
rect 217364 8428 217374 8484
rect 189746 8316 189756 8372
rect 189812 8316 196588 8372
rect 198818 8316 198828 8372
rect 198884 8316 199612 8372
rect 199668 8316 199678 8372
rect 201842 8316 201852 8372
rect 201908 8316 202972 8372
rect 203028 8316 203038 8372
rect 205202 8316 205212 8372
rect 205268 8316 205884 8372
rect 205940 8316 205950 8372
rect 208114 8316 208124 8372
rect 208180 8316 212156 8372
rect 212212 8316 212222 8372
rect 216962 8316 216972 8372
rect 217028 8316 218204 8372
rect 218260 8316 218270 8372
rect 221442 8316 221452 8372
rect 221508 8316 222012 8372
rect 222068 8316 225932 8372
rect 225988 8316 225998 8372
rect 196532 8260 196588 8316
rect 188626 8204 188636 8260
rect 188692 8204 189084 8260
rect 189140 8204 190764 8260
rect 190820 8204 190830 8260
rect 196532 8204 209468 8260
rect 209524 8204 210140 8260
rect 210196 8204 210206 8260
rect 210354 8204 210364 8260
rect 210420 8204 211148 8260
rect 211204 8204 211214 8260
rect 212370 8204 212380 8260
rect 212436 8204 213388 8260
rect 213444 8204 213454 8260
rect 200050 8092 200060 8148
rect 200116 8092 200844 8148
rect 200900 8092 202188 8148
rect 202244 8092 202254 8148
rect 202402 8092 202412 8148
rect 202468 8092 207340 8148
rect 207396 8092 207406 8148
rect 211362 8092 211372 8148
rect 211428 8092 212828 8148
rect 212884 8092 212894 8148
rect 217746 8092 217756 8148
rect 217812 8092 218092 8148
rect 218148 8092 220220 8148
rect 220276 8092 221004 8148
rect 221060 8092 221564 8148
rect 221620 8092 221630 8148
rect 187842 7980 187852 8036
rect 187908 7980 190428 8036
rect 190484 7980 199724 8036
rect 199780 7980 199790 8036
rect 200946 7980 200956 8036
rect 201012 7980 203420 8036
rect 203476 7980 204876 8036
rect 204932 7980 205772 8036
rect 205828 7980 205838 8036
rect 205986 7980 205996 8036
rect 206052 7980 206062 8036
rect 211250 7980 211260 8036
rect 211316 7980 211932 8036
rect 211988 7980 212716 8036
rect 212772 7980 212782 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 81266 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81550 7868
rect 111986 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112270 7868
rect 142706 7812 142716 7868
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142980 7812 142990 7868
rect 173426 7812 173436 7868
rect 173492 7812 173540 7868
rect 173596 7812 173644 7868
rect 173700 7812 173710 7868
rect 204146 7812 204156 7868
rect 204212 7812 204260 7868
rect 204316 7812 204364 7868
rect 204420 7812 204430 7868
rect 184772 7756 193340 7812
rect 193396 7756 193900 7812
rect 193956 7756 193966 7812
rect 184772 7700 184828 7756
rect 137890 7644 137900 7700
rect 137956 7644 184828 7700
rect 187618 7644 187628 7700
rect 187684 7644 188636 7700
rect 188692 7644 188702 7700
rect 189298 7644 189308 7700
rect 189364 7644 191324 7700
rect 191380 7644 191390 7700
rect 195346 7644 195356 7700
rect 195412 7644 199388 7700
rect 199444 7644 199454 7700
rect 205996 7588 206052 7980
rect 212146 7868 212156 7924
rect 212212 7868 220220 7924
rect 220276 7868 221228 7924
rect 221284 7868 221676 7924
rect 221732 7868 221742 7924
rect 234866 7812 234876 7868
rect 234932 7812 234980 7868
rect 235036 7812 235084 7868
rect 235140 7812 235150 7868
rect 265586 7812 265596 7868
rect 265652 7812 265700 7868
rect 265756 7812 265804 7868
rect 265860 7812 265870 7868
rect 296306 7812 296316 7868
rect 296372 7812 296420 7868
rect 296476 7812 296524 7868
rect 296580 7812 296590 7868
rect 206882 7756 206892 7812
rect 206948 7756 209804 7812
rect 209860 7756 216972 7812
rect 217028 7756 217038 7812
rect 220742 7756 220780 7812
rect 220836 7756 220846 7812
rect 220658 7644 220668 7700
rect 220724 7644 221788 7700
rect 221844 7644 221854 7700
rect 25106 7532 25116 7588
rect 25172 7532 71148 7588
rect 71204 7532 71214 7588
rect 182242 7532 182252 7588
rect 182308 7532 185388 7588
rect 185444 7532 185454 7588
rect 188066 7532 188076 7588
rect 188132 7532 191100 7588
rect 191156 7532 191166 7588
rect 195234 7532 195244 7588
rect 195300 7532 206052 7588
rect 211586 7532 211596 7588
rect 211652 7532 214060 7588
rect 214116 7532 214732 7588
rect 214788 7532 214798 7588
rect 184482 7420 184492 7476
rect 184548 7420 185612 7476
rect 185668 7420 185678 7476
rect 186274 7420 186284 7476
rect 186340 7420 187516 7476
rect 187572 7420 187582 7476
rect 190642 7420 190652 7476
rect 190708 7420 198548 7476
rect 199266 7420 199276 7476
rect 199332 7420 200396 7476
rect 200452 7420 202412 7476
rect 202468 7420 202478 7476
rect 202962 7420 202972 7476
rect 203028 7420 204652 7476
rect 204708 7420 204718 7476
rect 209458 7420 209468 7476
rect 209524 7420 210924 7476
rect 210980 7420 210990 7476
rect 216402 7420 216412 7476
rect 216468 7420 217756 7476
rect 217812 7420 217822 7476
rect 198492 7364 198548 7420
rect 198482 7308 198492 7364
rect 198548 7308 202860 7364
rect 202916 7308 202926 7364
rect 204866 7308 204876 7364
rect 204932 7308 214508 7364
rect 214564 7308 217196 7364
rect 217252 7308 217262 7364
rect 188290 7196 188300 7252
rect 188356 7196 189868 7252
rect 189924 7196 189934 7252
rect 199602 7196 199612 7252
rect 199668 7196 200172 7252
rect 200228 7196 209524 7252
rect 209468 7140 209524 7196
rect 209458 7084 209468 7140
rect 209524 7084 209534 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 96626 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96910 7084
rect 127346 7028 127356 7084
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127620 7028 127630 7084
rect 158066 7028 158076 7084
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158340 7028 158350 7084
rect 188786 7028 188796 7084
rect 188852 7028 188900 7084
rect 188956 7028 189004 7084
rect 189060 7028 189070 7084
rect 219506 7028 219516 7084
rect 219572 7028 219620 7084
rect 219676 7028 219724 7084
rect 219780 7028 219790 7084
rect 250226 7028 250236 7084
rect 250292 7028 250340 7084
rect 250396 7028 250444 7084
rect 250500 7028 250510 7084
rect 280946 7028 280956 7084
rect 281012 7028 281060 7084
rect 281116 7028 281164 7084
rect 281220 7028 281230 7084
rect 206098 6972 206108 7028
rect 206164 6972 216748 7028
rect 216804 6972 216814 7028
rect 145058 6860 145068 6916
rect 145124 6860 173068 6916
rect 186722 6860 186732 6916
rect 186788 6860 196588 6916
rect 201170 6860 201180 6916
rect 201236 6860 204988 6916
rect 205044 6860 213836 6916
rect 213892 6860 214620 6916
rect 214676 6860 214686 6916
rect 173012 6804 173068 6860
rect 196532 6804 196588 6860
rect 173012 6748 190708 6804
rect 190866 6748 190876 6804
rect 190932 6748 192892 6804
rect 192948 6748 192958 6804
rect 196532 6748 210588 6804
rect 210644 6748 210654 6804
rect 217186 6748 217196 6804
rect 217252 6748 218204 6804
rect 218260 6748 218270 6804
rect 190652 6580 190708 6748
rect 190978 6636 190988 6692
rect 191044 6636 193228 6692
rect 193284 6636 193294 6692
rect 196532 6636 199836 6692
rect 199892 6636 201628 6692
rect 201684 6636 201694 6692
rect 202962 6636 202972 6692
rect 203028 6636 204428 6692
rect 204484 6636 204494 6692
rect 204642 6636 204652 6692
rect 204708 6636 207452 6692
rect 207508 6636 207518 6692
rect 190652 6524 192668 6580
rect 192724 6524 192734 6580
rect 196532 6468 196588 6636
rect 202850 6524 202860 6580
rect 202916 6524 205100 6580
rect 205156 6524 205166 6580
rect 148642 6412 148652 6468
rect 148708 6412 184044 6468
rect 184100 6412 184110 6468
rect 190306 6412 190316 6468
rect 190372 6412 192780 6468
rect 192836 6412 193116 6468
rect 193172 6412 193182 6468
rect 196018 6412 196028 6468
rect 196084 6412 196588 6468
rect 203074 6412 203084 6468
rect 203140 6412 207900 6468
rect 207956 6412 207966 6468
rect 213602 6412 213612 6468
rect 213668 6412 217644 6468
rect 217700 6412 218876 6468
rect 218932 6412 218942 6468
rect 187506 6300 187516 6356
rect 187572 6300 189420 6356
rect 189476 6300 195244 6356
rect 195300 6300 195310 6356
rect 204530 6300 204540 6356
rect 204596 6300 204764 6356
rect 204820 6300 207004 6356
rect 207060 6300 207070 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 81266 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81550 6300
rect 111986 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112270 6300
rect 142706 6244 142716 6300
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142980 6244 142990 6300
rect 173426 6244 173436 6300
rect 173492 6244 173540 6300
rect 173596 6244 173644 6300
rect 173700 6244 173710 6300
rect 204146 6244 204156 6300
rect 204212 6244 204260 6300
rect 204316 6244 204364 6300
rect 204420 6244 204430 6300
rect 234866 6244 234876 6300
rect 234932 6244 234980 6300
rect 235036 6244 235084 6300
rect 235140 6244 235150 6300
rect 265586 6244 265596 6300
rect 265652 6244 265700 6300
rect 265756 6244 265804 6300
rect 265860 6244 265870 6300
rect 296306 6244 296316 6300
rect 296372 6244 296420 6300
rect 296476 6244 296524 6300
rect 296580 6244 296590 6300
rect 141474 6076 141484 6132
rect 141540 6076 191660 6132
rect 191716 6076 191726 6132
rect 195346 6076 195356 6132
rect 195412 6076 197708 6132
rect 197764 6076 197774 6132
rect 203522 6076 203532 6132
rect 203588 6076 204540 6132
rect 204596 6076 205548 6132
rect 205604 6076 205614 6132
rect 217858 6076 217868 6132
rect 217924 6076 219100 6132
rect 219156 6076 263004 6132
rect 263060 6076 263070 6132
rect 187506 5964 187516 6020
rect 187572 5964 187964 6020
rect 188020 5964 188030 6020
rect 191762 5964 191772 6020
rect 191828 5964 192892 6020
rect 192948 5964 192958 6020
rect 199714 5964 199724 6020
rect 199780 5964 204652 6020
rect 204708 5964 204718 6020
rect 207442 5964 207452 6020
rect 207508 5964 292124 6020
rect 292180 5964 292190 6020
rect 56578 5852 56588 5908
rect 56644 5852 93548 5908
rect 93604 5852 93614 5908
rect 182354 5852 182364 5908
rect 182420 5852 183708 5908
rect 183764 5852 183774 5908
rect 184594 5852 184604 5908
rect 184660 5852 186732 5908
rect 186788 5852 186798 5908
rect 191090 5852 191100 5908
rect 191156 5852 196028 5908
rect 196084 5852 196094 5908
rect 200610 5852 200620 5908
rect 200676 5852 204876 5908
rect 204932 5852 204942 5908
rect 205762 5852 205772 5908
rect 205828 5852 206556 5908
rect 206612 5852 206622 5908
rect 209458 5852 209468 5908
rect 209524 5852 210364 5908
rect 210420 5852 210430 5908
rect 211250 5852 211260 5908
rect 211316 5852 215292 5908
rect 215348 5852 215358 5908
rect 210364 5796 210420 5852
rect 189186 5740 189196 5796
rect 189252 5740 190428 5796
rect 190484 5740 192332 5796
rect 192388 5740 192398 5796
rect 199714 5740 199724 5796
rect 199780 5740 203980 5796
rect 204036 5740 204046 5796
rect 204978 5740 204988 5796
rect 205044 5740 205548 5796
rect 205604 5740 206444 5796
rect 206500 5740 206510 5796
rect 210364 5740 215852 5796
rect 215908 5740 215918 5796
rect 216402 5740 216412 5796
rect 216468 5740 217084 5796
rect 217140 5740 234332 5796
rect 234388 5740 234398 5796
rect 186386 5628 186396 5684
rect 186452 5628 188860 5684
rect 188916 5628 190652 5684
rect 190708 5628 190718 5684
rect 198146 5628 198156 5684
rect 198212 5628 202972 5684
rect 203028 5628 203038 5684
rect 206210 5628 206220 5684
rect 206276 5628 207564 5684
rect 207620 5628 207630 5684
rect 203858 5516 203868 5572
rect 203924 5516 205212 5572
rect 205268 5516 205772 5572
rect 205828 5516 205838 5572
rect 205996 5516 208796 5572
rect 208852 5516 210700 5572
rect 210756 5516 210766 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 96626 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96910 5516
rect 127346 5460 127356 5516
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127620 5460 127630 5516
rect 158066 5460 158076 5516
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158340 5460 158350 5516
rect 188786 5460 188796 5516
rect 188852 5460 188900 5516
rect 188956 5460 189004 5516
rect 189060 5460 189070 5516
rect 205996 5460 206052 5516
rect 219506 5460 219516 5516
rect 219572 5460 219620 5516
rect 219676 5460 219724 5516
rect 219780 5460 219790 5516
rect 250226 5460 250236 5516
rect 250292 5460 250340 5516
rect 250396 5460 250444 5516
rect 250500 5460 250510 5516
rect 280946 5460 280956 5516
rect 281012 5460 281060 5516
rect 281116 5460 281164 5516
rect 281220 5460 281230 5516
rect 185378 5404 185388 5460
rect 185444 5404 187068 5460
rect 187124 5404 187134 5460
rect 192658 5404 192668 5460
rect 192724 5404 195020 5460
rect 195076 5404 195086 5460
rect 200946 5404 200956 5460
rect 201012 5404 203980 5460
rect 204036 5404 205996 5460
rect 206052 5404 206062 5460
rect 206556 5404 211596 5460
rect 211652 5404 211662 5460
rect 184706 5292 184716 5348
rect 184772 5292 187404 5348
rect 187460 5292 187470 5348
rect 190306 5292 190316 5348
rect 190372 5292 195468 5348
rect 195524 5292 195534 5348
rect 200834 5292 200844 5348
rect 200900 5292 202972 5348
rect 203028 5292 203038 5348
rect 206556 5236 206612 5404
rect 207330 5292 207340 5348
rect 207396 5292 208348 5348
rect 215954 5292 215964 5348
rect 216020 5292 231868 5348
rect 173012 5180 185948 5236
rect 186004 5180 186014 5236
rect 190642 5180 190652 5236
rect 190708 5180 191660 5236
rect 191716 5180 191726 5236
rect 192322 5180 192332 5236
rect 192388 5180 193676 5236
rect 193732 5180 193742 5236
rect 194562 5180 194572 5236
rect 194628 5180 195244 5236
rect 195300 5180 195310 5236
rect 196802 5180 196812 5236
rect 196868 5180 201068 5236
rect 201124 5180 201852 5236
rect 201908 5180 201918 5236
rect 206546 5180 206556 5236
rect 206612 5180 206622 5236
rect 173012 5124 173068 5180
rect 208292 5124 208348 5292
rect 231812 5236 231868 5292
rect 214722 5180 214732 5236
rect 214788 5180 215628 5236
rect 215684 5180 215694 5236
rect 218530 5180 218540 5236
rect 218596 5180 222572 5236
rect 222628 5180 223468 5236
rect 223524 5180 223534 5236
rect 231812 5180 245420 5236
rect 245476 5180 245486 5236
rect 122546 5068 122556 5124
rect 122612 5068 173068 5124
rect 186162 5068 186172 5124
rect 186228 5068 189868 5124
rect 189924 5068 189934 5124
rect 190978 5068 190988 5124
rect 191044 5068 194348 5124
rect 194404 5068 194414 5124
rect 195122 5068 195132 5124
rect 195188 5068 197708 5124
rect 197764 5068 197774 5124
rect 201730 5068 201740 5124
rect 201796 5068 203084 5124
rect 203140 5068 203150 5124
rect 206322 5068 206332 5124
rect 206388 5068 207340 5124
rect 207396 5068 207406 5124
rect 208292 5068 209468 5124
rect 209524 5068 209534 5124
rect 209906 5068 209916 5124
rect 209972 5068 216188 5124
rect 216244 5068 216254 5124
rect 217746 5068 217756 5124
rect 217812 5068 218988 5124
rect 219044 5068 219054 5124
rect 221554 5068 221564 5124
rect 221620 5068 224028 5124
rect 224084 5068 224094 5124
rect 183586 4956 183596 5012
rect 183652 4956 184604 5012
rect 184660 4956 184670 5012
rect 186610 4956 186620 5012
rect 186676 4956 187628 5012
rect 187684 4956 187694 5012
rect 197586 4956 197596 5012
rect 197652 4956 199164 5012
rect 199220 4956 199230 5012
rect 205986 4956 205996 5012
rect 206052 4956 207228 5012
rect 207284 4956 213612 5012
rect 213668 4956 213678 5012
rect 215170 4956 215180 5012
rect 215236 4956 216076 5012
rect 216132 4956 216636 5012
rect 216692 4956 217084 5012
rect 217140 4956 217150 5012
rect 217308 4956 241612 5012
rect 241668 4956 241678 5012
rect 217308 4900 217364 4956
rect 134306 4844 134316 4900
rect 134372 4844 184828 4900
rect 186162 4844 186172 4900
rect 186228 4844 187404 4900
rect 187460 4844 187470 4900
rect 194786 4844 194796 4900
rect 194852 4844 196140 4900
rect 196196 4844 196206 4900
rect 200396 4844 204092 4900
rect 204148 4844 204652 4900
rect 204708 4844 204718 4900
rect 206210 4844 206220 4900
rect 206276 4844 207004 4900
rect 207060 4844 207070 4900
rect 208898 4844 208908 4900
rect 208964 4844 210252 4900
rect 210308 4844 210318 4900
rect 216290 4844 216300 4900
rect 216356 4844 216860 4900
rect 216916 4844 216926 4900
rect 217074 4844 217084 4900
rect 217140 4844 217364 4900
rect 220658 4844 220668 4900
rect 220724 4844 221788 4900
rect 221844 4844 221854 4900
rect 222114 4844 222124 4900
rect 222180 4844 223132 4900
rect 223188 4844 223198 4900
rect 184772 4788 184828 4844
rect 184772 4732 190316 4788
rect 190372 4732 190382 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 81266 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81550 4732
rect 111986 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112270 4732
rect 142706 4676 142716 4732
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142980 4676 142990 4732
rect 173426 4676 173436 4732
rect 173492 4676 173540 4732
rect 173596 4676 173644 4732
rect 173700 4676 173710 4732
rect 189410 4620 189420 4676
rect 189476 4620 196364 4676
rect 196420 4620 198156 4676
rect 198212 4620 198222 4676
rect 91634 4508 91644 4564
rect 91700 4508 96236 4564
rect 96292 4508 96302 4564
rect 173730 4508 173740 4564
rect 173796 4508 196980 4564
rect 197138 4508 197148 4564
rect 197204 4508 197932 4564
rect 197988 4508 199500 4564
rect 199556 4508 199566 4564
rect 196924 4452 196980 4508
rect 200396 4452 200452 4844
rect 208908 4788 208964 4844
rect 208226 4732 208236 4788
rect 208292 4732 208964 4788
rect 211026 4732 211036 4788
rect 211092 4732 212492 4788
rect 212548 4732 220108 4788
rect 220164 4732 220556 4788
rect 220612 4732 220622 4788
rect 223010 4732 223020 4788
rect 223076 4732 223916 4788
rect 223972 4732 223982 4788
rect 204146 4676 204156 4732
rect 204212 4676 204260 4732
rect 204316 4676 204364 4732
rect 204420 4676 204430 4732
rect 223020 4676 223076 4732
rect 234866 4676 234876 4732
rect 234932 4676 234980 4732
rect 235036 4676 235084 4732
rect 235140 4676 235150 4732
rect 265586 4676 265596 4732
rect 265652 4676 265700 4732
rect 265756 4676 265804 4732
rect 265860 4676 265870 4732
rect 296306 4676 296316 4732
rect 296372 4676 296420 4732
rect 296476 4676 296524 4732
rect 296580 4676 296590 4732
rect 214498 4620 214508 4676
rect 214564 4620 215292 4676
rect 215348 4620 223076 4676
rect 200610 4508 200620 4564
rect 200676 4508 208012 4564
rect 208068 4508 208078 4564
rect 212370 4508 212380 4564
rect 212436 4508 215404 4564
rect 215460 4508 215470 4564
rect 215954 4508 215964 4564
rect 216020 4508 217084 4564
rect 217140 4508 217150 4564
rect 217298 4508 217308 4564
rect 217364 4508 230748 4564
rect 230804 4508 230814 4564
rect 85026 4396 85036 4452
rect 85092 4396 86716 4452
rect 86772 4396 86782 4452
rect 96786 4396 96796 4452
rect 96852 4396 97580 4452
rect 97636 4396 97646 4452
rect 187954 4396 187964 4452
rect 188020 4396 188300 4452
rect 188356 4396 188860 4452
rect 188916 4396 190540 4452
rect 190596 4396 190606 4452
rect 193452 4396 196700 4452
rect 196756 4396 196766 4452
rect 196924 4396 200452 4452
rect 201730 4396 201740 4452
rect 201796 4396 202076 4452
rect 202132 4396 202972 4452
rect 203028 4396 204540 4452
rect 204596 4396 205100 4452
rect 205156 4396 205166 4452
rect 209794 4396 209804 4452
rect 209860 4396 210812 4452
rect 210868 4396 211596 4452
rect 211652 4396 211932 4452
rect 211988 4396 211998 4452
rect 216738 4396 216748 4452
rect 216804 4396 217532 4452
rect 217588 4396 219548 4452
rect 219604 4396 219614 4452
rect 219772 4396 220668 4452
rect 220724 4396 220734 4452
rect 228498 4396 228508 4452
rect 228564 4396 288540 4452
rect 288596 4396 288606 4452
rect 193452 4340 193508 4396
rect 219772 4340 219828 4396
rect 75394 4284 75404 4340
rect 75460 4284 76636 4340
rect 76692 4284 76702 4340
rect 87042 4284 87052 4340
rect 87108 4284 87948 4340
rect 88004 4284 88014 4340
rect 89618 4284 89628 4340
rect 89684 4284 90972 4340
rect 91028 4284 91038 4340
rect 182802 4284 182812 4340
rect 182868 4284 183708 4340
rect 183764 4284 183774 4340
rect 193442 4284 193452 4340
rect 193508 4284 193518 4340
rect 196532 4284 197708 4340
rect 197764 4284 197774 4340
rect 205314 4284 205324 4340
rect 205380 4284 205548 4340
rect 205604 4284 206220 4340
rect 206276 4284 206286 4340
rect 208338 4284 208348 4340
rect 208404 4284 209020 4340
rect 209076 4284 210028 4340
rect 210084 4284 211148 4340
rect 211204 4284 211214 4340
rect 216514 4284 216524 4340
rect 216580 4284 217980 4340
rect 218036 4284 218046 4340
rect 218876 4284 219828 4340
rect 220770 4284 220780 4340
rect 220836 4284 221900 4340
rect 221956 4284 221966 4340
rect 223234 4284 223244 4340
rect 223300 4284 223692 4340
rect 223748 4284 249228 4340
rect 249284 4284 249294 4340
rect 196532 4228 196588 4284
rect 87154 4172 87164 4228
rect 87220 4172 89068 4228
rect 89124 4172 89134 4228
rect 152226 4172 152236 4228
rect 152292 4172 186284 4228
rect 186340 4172 186350 4228
rect 191650 4172 191660 4228
rect 191716 4172 196588 4228
rect 201170 4172 201180 4228
rect 201236 4172 205884 4228
rect 205940 4172 205950 4228
rect 218876 4116 218932 4284
rect 219090 4172 219100 4228
rect 219156 4172 219324 4228
rect 219380 4172 220108 4228
rect 220164 4172 220174 4228
rect 220322 4172 220332 4228
rect 220388 4172 223132 4228
rect 223188 4172 223198 4228
rect 76402 4060 76412 4116
rect 76468 4060 77644 4116
rect 77700 4060 77710 4116
rect 79986 4060 79996 4116
rect 80052 4060 81228 4116
rect 81284 4060 81294 4116
rect 83570 4060 83580 4116
rect 83636 4060 84812 4116
rect 84868 4060 84878 4116
rect 90738 4060 90748 4116
rect 90804 4060 91980 4116
rect 92036 4060 92046 4116
rect 123890 4060 123900 4116
rect 123956 4060 181580 4116
rect 181636 4060 182252 4116
rect 182308 4060 182318 4116
rect 192770 4060 192780 4116
rect 192836 4060 195804 4116
rect 195860 4060 195870 4116
rect 204530 4060 204540 4116
rect 204596 4060 218932 4116
rect 219538 4060 219548 4116
rect 219604 4060 220276 4116
rect 223346 4060 223356 4116
rect 223412 4060 253036 4116
rect 253092 4060 253102 4116
rect 220220 4004 220276 4060
rect 201282 3948 201292 4004
rect 201348 3948 208124 4004
rect 208180 3948 208190 4004
rect 220210 3948 220220 4004
rect 220276 3948 220892 4004
rect 220948 3948 220958 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 96626 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96910 3948
rect 127346 3892 127356 3948
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127620 3892 127630 3948
rect 158066 3892 158076 3948
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158340 3892 158350 3948
rect 188786 3892 188796 3948
rect 188852 3892 188900 3948
rect 188956 3892 189004 3948
rect 189060 3892 189070 3948
rect 219506 3892 219516 3948
rect 219572 3892 219620 3948
rect 219676 3892 219724 3948
rect 219780 3892 219790 3948
rect 250226 3892 250236 3948
rect 250292 3892 250340 3948
rect 250396 3892 250444 3948
rect 250500 3892 250510 3948
rect 280946 3892 280956 3948
rect 281012 3892 281060 3948
rect 281116 3892 281164 3948
rect 281220 3892 281230 3948
rect 170146 3836 170156 3892
rect 170212 3836 188692 3892
rect 201842 3836 201852 3892
rect 201908 3836 205660 3892
rect 205716 3836 206108 3892
rect 206164 3836 206174 3892
rect 188636 3780 188692 3836
rect 131506 3724 131516 3780
rect 131572 3724 182028 3780
rect 182084 3724 182094 3780
rect 183922 3724 183932 3780
rect 183988 3724 187516 3780
rect 187572 3724 187582 3780
rect 188636 3724 204204 3780
rect 204260 3724 206668 3780
rect 206724 3724 206734 3780
rect 208292 3724 212828 3780
rect 212884 3724 212894 3780
rect 216850 3724 216860 3780
rect 216916 3724 237916 3780
rect 237972 3724 237982 3780
rect 243572 3724 255836 3780
rect 255892 3724 255902 3780
rect 267092 3724 281372 3780
rect 281428 3724 281438 3780
rect 208292 3668 208348 3724
rect 243572 3668 243628 3724
rect 267092 3668 267148 3724
rect 43026 3612 43036 3668
rect 43092 3612 43820 3668
rect 43876 3612 43886 3668
rect 46834 3612 46844 3668
rect 46900 3612 47628 3668
rect 47684 3612 47694 3668
rect 62066 3612 62076 3668
rect 62132 3612 62860 3668
rect 62916 3612 62926 3668
rect 65202 3612 65212 3668
rect 65268 3612 65772 3668
rect 65828 3612 68236 3668
rect 68292 3612 68302 3668
rect 69234 3612 69244 3668
rect 69300 3612 70476 3668
rect 70532 3612 70542 3668
rect 181010 3612 181020 3668
rect 181076 3612 189868 3668
rect 189924 3612 189934 3668
rect 199042 3612 199052 3668
rect 199108 3612 201292 3668
rect 201348 3612 201358 3668
rect 205650 3612 205660 3668
rect 205716 3612 208348 3668
rect 220546 3612 220556 3668
rect 220612 3612 221452 3668
rect 221508 3612 221518 3668
rect 224690 3612 224700 3668
rect 224756 3612 243628 3668
rect 249330 3612 249340 3668
rect 249396 3612 267148 3668
rect 50530 3500 50540 3556
rect 50596 3500 59612 3556
rect 59668 3500 59678 3556
rect 68898 3500 68908 3556
rect 68964 3500 69580 3556
rect 69636 3500 69646 3556
rect 71698 3500 71708 3556
rect 71764 3500 74060 3556
rect 74116 3500 74126 3556
rect 88722 3500 88732 3556
rect 88788 3500 89404 3556
rect 89460 3500 89470 3556
rect 111458 3500 111468 3556
rect 111524 3500 111804 3556
rect 111860 3500 112812 3556
rect 112868 3500 112878 3556
rect 115042 3500 115052 3556
rect 115108 3500 115388 3556
rect 115444 3500 124348 3556
rect 124404 3500 124414 3556
rect 127698 3500 127708 3556
rect 127764 3500 182812 3556
rect 182868 3500 182878 3556
rect 185938 3500 185948 3556
rect 186004 3500 186732 3556
rect 186788 3500 186798 3556
rect 195346 3500 195356 3556
rect 195412 3500 197652 3556
rect 202402 3500 202412 3556
rect 202468 3500 203532 3556
rect 203588 3500 203598 3556
rect 204876 3500 210588 3556
rect 210644 3500 210654 3556
rect 210812 3500 212044 3556
rect 212100 3500 212110 3556
rect 212258 3500 212268 3556
rect 212324 3500 216468 3556
rect 220434 3500 220444 3556
rect 220500 3500 223916 3556
rect 223972 3500 223982 3556
rect 225922 3500 225932 3556
rect 225988 3500 285068 3556
rect 285124 3500 285134 3556
rect 197596 3444 197652 3500
rect 204876 3444 204932 3500
rect 210812 3444 210868 3500
rect 8306 3388 8316 3444
rect 8372 3388 10108 3444
rect 10164 3388 10174 3444
rect 65650 3388 65660 3444
rect 65716 3388 66668 3444
rect 66724 3388 66734 3444
rect 72930 3388 72940 3444
rect 72996 3388 75628 3444
rect 75684 3388 75694 3444
rect 103954 3388 103964 3444
rect 104020 3388 104748 3444
rect 104804 3388 107492 3444
rect 107762 3388 107772 3444
rect 107828 3388 108556 3444
rect 108612 3388 109340 3444
rect 109396 3388 109406 3444
rect 166562 3388 166572 3444
rect 166628 3388 169932 3444
rect 169988 3388 169998 3444
rect 187842 3388 187852 3444
rect 187908 3388 188524 3444
rect 188580 3388 188590 3444
rect 194674 3388 194684 3444
rect 194740 3388 195916 3444
rect 195972 3388 197148 3444
rect 197204 3388 197214 3444
rect 197586 3388 197596 3444
rect 197652 3388 197662 3444
rect 198706 3388 198716 3444
rect 198772 3388 200396 3444
rect 200452 3388 202748 3444
rect 202804 3388 202814 3444
rect 204866 3388 204876 3444
rect 204932 3388 204942 3444
rect 205650 3388 205660 3444
rect 205716 3388 207564 3444
rect 207620 3388 208460 3444
rect 208516 3388 208526 3444
rect 209122 3388 209132 3444
rect 209188 3388 210028 3444
rect 210084 3388 210868 3444
rect 211362 3388 211372 3444
rect 211428 3388 212828 3444
rect 212884 3388 212894 3444
rect 107436 3332 107492 3388
rect 216412 3332 216468 3500
rect 221218 3388 221228 3444
rect 221284 3388 227220 3444
rect 244962 3388 244972 3444
rect 245028 3388 245644 3444
rect 245700 3388 245710 3444
rect 248770 3388 248780 3444
rect 248836 3388 249452 3444
rect 249508 3388 249518 3444
rect 265346 3388 265356 3444
rect 265412 3388 267036 3444
rect 267092 3388 267102 3444
rect 227164 3332 227220 3388
rect 107436 3276 184828 3332
rect 184884 3276 184894 3332
rect 216402 3276 216412 3332
rect 216468 3276 216478 3332
rect 227154 3276 227164 3332
rect 227220 3276 227230 3332
rect 231812 3276 277900 3332
rect 277956 3276 277966 3332
rect 231812 3220 231868 3276
rect 208002 3164 208012 3220
rect 208068 3164 231868 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 81266 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81550 3164
rect 111986 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112270 3164
rect 142706 3108 142716 3164
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142980 3108 142990 3164
rect 173426 3108 173436 3164
rect 173492 3108 173540 3164
rect 173596 3108 173644 3164
rect 173700 3108 173710 3164
rect 204146 3108 204156 3164
rect 204212 3108 204260 3164
rect 204316 3108 204364 3164
rect 204420 3108 204430 3164
rect 234866 3108 234876 3164
rect 234932 3108 234980 3164
rect 235036 3108 235084 3164
rect 235140 3108 235150 3164
rect 265586 3108 265596 3164
rect 265652 3108 265700 3164
rect 265756 3108 265804 3164
rect 265860 3108 265870 3164
rect 296306 3108 296316 3164
rect 296372 3108 296420 3164
rect 296476 3108 296524 3164
rect 296580 3108 296590 3164
rect 204754 2940 204764 2996
rect 204820 2940 225932 2996
rect 225988 2940 225998 2996
rect 162978 2828 162988 2884
rect 163044 2828 198716 2884
rect 198772 2828 198782 2884
rect 203186 2828 203196 2884
rect 203252 2828 222012 2884
rect 222068 2828 222078 2884
rect 169922 2716 169932 2772
rect 169988 2716 200844 2772
rect 200900 2716 200910 2772
rect 203074 2716 203084 2772
rect 203140 2716 219100 2772
rect 219156 2716 219166 2772
rect 220098 2716 220108 2772
rect 220164 2716 259420 2772
rect 259476 2716 259486 2772
rect 186274 2604 186284 2660
rect 186340 2604 207340 2660
rect 207396 2604 207406 2660
rect 178882 2492 178892 2548
rect 178948 2492 193340 2548
rect 193396 2492 193406 2548
rect 198706 2492 198716 2548
rect 198772 2492 228508 2548
rect 228564 2492 228574 2548
rect 156258 2380 156268 2436
rect 156324 2380 205772 2436
rect 205828 2380 205838 2436
rect 112802 2268 112812 2324
rect 112868 2268 186844 2324
rect 186900 2268 186910 2324
rect 187058 2268 187068 2324
rect 187124 2268 211820 2324
rect 211876 2268 211886 2324
rect 186722 2156 186732 2212
rect 186788 2156 210476 2212
rect 210532 2156 210542 2212
rect 197586 2044 197596 2100
rect 197652 2044 221116 2100
rect 221172 2044 221182 2100
rect 159618 1932 159628 1988
rect 159684 1932 204876 1988
rect 204932 1932 204942 1988
rect 195794 1596 195804 1652
rect 195860 1596 265356 1652
rect 265412 1596 265422 1652
rect 124338 1484 124348 1540
rect 124404 1484 210364 1540
rect 210420 1484 210430 1540
rect 192994 1372 193004 1428
rect 193060 1372 274316 1428
rect 274372 1372 274382 1428
rect 201282 1260 201292 1316
rect 201348 1260 249340 1316
rect 249396 1260 249406 1316
rect 177314 1148 177324 1204
rect 177380 1148 205996 1204
rect 206052 1148 206062 1204
rect 109330 1036 109340 1092
rect 109396 1036 206892 1092
rect 206948 1036 206958 1092
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 81276 56420 81332 56476
rect 81380 56420 81436 56476
rect 81484 56420 81540 56476
rect 111996 56420 112052 56476
rect 112100 56420 112156 56476
rect 112204 56420 112260 56476
rect 142716 56420 142772 56476
rect 142820 56420 142876 56476
rect 142924 56420 142980 56476
rect 173436 56420 173492 56476
rect 173540 56420 173596 56476
rect 173644 56420 173700 56476
rect 204156 56420 204212 56476
rect 204260 56420 204316 56476
rect 204364 56420 204420 56476
rect 234876 56420 234932 56476
rect 234980 56420 235036 56476
rect 235084 56420 235140 56476
rect 265596 56420 265652 56476
rect 265700 56420 265756 56476
rect 265804 56420 265860 56476
rect 296316 56420 296372 56476
rect 296420 56420 296476 56476
rect 296524 56420 296580 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 96636 55636 96692 55692
rect 96740 55636 96796 55692
rect 96844 55636 96900 55692
rect 127356 55636 127412 55692
rect 127460 55636 127516 55692
rect 127564 55636 127620 55692
rect 158076 55636 158132 55692
rect 158180 55636 158236 55692
rect 158284 55636 158340 55692
rect 188796 55636 188852 55692
rect 188900 55636 188956 55692
rect 189004 55636 189060 55692
rect 219516 55636 219572 55692
rect 219620 55636 219676 55692
rect 219724 55636 219780 55692
rect 250236 55636 250292 55692
rect 250340 55636 250396 55692
rect 250444 55636 250500 55692
rect 280956 55636 281012 55692
rect 281060 55636 281116 55692
rect 281164 55636 281220 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 81276 54852 81332 54908
rect 81380 54852 81436 54908
rect 81484 54852 81540 54908
rect 111996 54852 112052 54908
rect 112100 54852 112156 54908
rect 112204 54852 112260 54908
rect 142716 54852 142772 54908
rect 142820 54852 142876 54908
rect 142924 54852 142980 54908
rect 173436 54852 173492 54908
rect 173540 54852 173596 54908
rect 173644 54852 173700 54908
rect 204156 54852 204212 54908
rect 204260 54852 204316 54908
rect 204364 54852 204420 54908
rect 234876 54852 234932 54908
rect 234980 54852 235036 54908
rect 235084 54852 235140 54908
rect 265596 54852 265652 54908
rect 265700 54852 265756 54908
rect 265804 54852 265860 54908
rect 296316 54852 296372 54908
rect 296420 54852 296476 54908
rect 296524 54852 296580 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 96636 54068 96692 54124
rect 96740 54068 96796 54124
rect 96844 54068 96900 54124
rect 127356 54068 127412 54124
rect 127460 54068 127516 54124
rect 127564 54068 127620 54124
rect 158076 54068 158132 54124
rect 158180 54068 158236 54124
rect 158284 54068 158340 54124
rect 188796 54068 188852 54124
rect 188900 54068 188956 54124
rect 189004 54068 189060 54124
rect 219516 54068 219572 54124
rect 219620 54068 219676 54124
rect 219724 54068 219780 54124
rect 250236 54068 250292 54124
rect 250340 54068 250396 54124
rect 250444 54068 250500 54124
rect 280956 54068 281012 54124
rect 281060 54068 281116 54124
rect 281164 54068 281220 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 81276 53284 81332 53340
rect 81380 53284 81436 53340
rect 81484 53284 81540 53340
rect 111996 53284 112052 53340
rect 112100 53284 112156 53340
rect 112204 53284 112260 53340
rect 142716 53284 142772 53340
rect 142820 53284 142876 53340
rect 142924 53284 142980 53340
rect 173436 53284 173492 53340
rect 173540 53284 173596 53340
rect 173644 53284 173700 53340
rect 204156 53284 204212 53340
rect 204260 53284 204316 53340
rect 204364 53284 204420 53340
rect 234876 53284 234932 53340
rect 234980 53284 235036 53340
rect 235084 53284 235140 53340
rect 265596 53284 265652 53340
rect 265700 53284 265756 53340
rect 265804 53284 265860 53340
rect 296316 53284 296372 53340
rect 296420 53284 296476 53340
rect 296524 53284 296580 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 96636 52500 96692 52556
rect 96740 52500 96796 52556
rect 96844 52500 96900 52556
rect 127356 52500 127412 52556
rect 127460 52500 127516 52556
rect 127564 52500 127620 52556
rect 158076 52500 158132 52556
rect 158180 52500 158236 52556
rect 158284 52500 158340 52556
rect 188796 52500 188852 52556
rect 188900 52500 188956 52556
rect 189004 52500 189060 52556
rect 219516 52500 219572 52556
rect 219620 52500 219676 52556
rect 219724 52500 219780 52556
rect 250236 52500 250292 52556
rect 250340 52500 250396 52556
rect 250444 52500 250500 52556
rect 280956 52500 281012 52556
rect 281060 52500 281116 52556
rect 281164 52500 281220 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 81276 51716 81332 51772
rect 81380 51716 81436 51772
rect 81484 51716 81540 51772
rect 111996 51716 112052 51772
rect 112100 51716 112156 51772
rect 112204 51716 112260 51772
rect 142716 51716 142772 51772
rect 142820 51716 142876 51772
rect 142924 51716 142980 51772
rect 173436 51716 173492 51772
rect 173540 51716 173596 51772
rect 173644 51716 173700 51772
rect 204156 51716 204212 51772
rect 204260 51716 204316 51772
rect 204364 51716 204420 51772
rect 234876 51716 234932 51772
rect 234980 51716 235036 51772
rect 235084 51716 235140 51772
rect 265596 51716 265652 51772
rect 265700 51716 265756 51772
rect 265804 51716 265860 51772
rect 296316 51716 296372 51772
rect 296420 51716 296476 51772
rect 296524 51716 296580 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 96636 50932 96692 50988
rect 96740 50932 96796 50988
rect 96844 50932 96900 50988
rect 127356 50932 127412 50988
rect 127460 50932 127516 50988
rect 127564 50932 127620 50988
rect 158076 50932 158132 50988
rect 158180 50932 158236 50988
rect 158284 50932 158340 50988
rect 188796 50932 188852 50988
rect 188900 50932 188956 50988
rect 189004 50932 189060 50988
rect 219516 50932 219572 50988
rect 219620 50932 219676 50988
rect 219724 50932 219780 50988
rect 250236 50932 250292 50988
rect 250340 50932 250396 50988
rect 250444 50932 250500 50988
rect 280956 50932 281012 50988
rect 281060 50932 281116 50988
rect 281164 50932 281220 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 81276 50148 81332 50204
rect 81380 50148 81436 50204
rect 81484 50148 81540 50204
rect 111996 50148 112052 50204
rect 112100 50148 112156 50204
rect 112204 50148 112260 50204
rect 142716 50148 142772 50204
rect 142820 50148 142876 50204
rect 142924 50148 142980 50204
rect 173436 50148 173492 50204
rect 173540 50148 173596 50204
rect 173644 50148 173700 50204
rect 204156 50148 204212 50204
rect 204260 50148 204316 50204
rect 204364 50148 204420 50204
rect 234876 50148 234932 50204
rect 234980 50148 235036 50204
rect 235084 50148 235140 50204
rect 265596 50148 265652 50204
rect 265700 50148 265756 50204
rect 265804 50148 265860 50204
rect 296316 50148 296372 50204
rect 296420 50148 296476 50204
rect 296524 50148 296580 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 96636 49364 96692 49420
rect 96740 49364 96796 49420
rect 96844 49364 96900 49420
rect 127356 49364 127412 49420
rect 127460 49364 127516 49420
rect 127564 49364 127620 49420
rect 158076 49364 158132 49420
rect 158180 49364 158236 49420
rect 158284 49364 158340 49420
rect 188796 49364 188852 49420
rect 188900 49364 188956 49420
rect 189004 49364 189060 49420
rect 219516 49364 219572 49420
rect 219620 49364 219676 49420
rect 219724 49364 219780 49420
rect 250236 49364 250292 49420
rect 250340 49364 250396 49420
rect 250444 49364 250500 49420
rect 280956 49364 281012 49420
rect 281060 49364 281116 49420
rect 281164 49364 281220 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 81276 48580 81332 48636
rect 81380 48580 81436 48636
rect 81484 48580 81540 48636
rect 111996 48580 112052 48636
rect 112100 48580 112156 48636
rect 112204 48580 112260 48636
rect 142716 48580 142772 48636
rect 142820 48580 142876 48636
rect 142924 48580 142980 48636
rect 173436 48580 173492 48636
rect 173540 48580 173596 48636
rect 173644 48580 173700 48636
rect 204156 48580 204212 48636
rect 204260 48580 204316 48636
rect 204364 48580 204420 48636
rect 234876 48580 234932 48636
rect 234980 48580 235036 48636
rect 235084 48580 235140 48636
rect 265596 48580 265652 48636
rect 265700 48580 265756 48636
rect 265804 48580 265860 48636
rect 296316 48580 296372 48636
rect 296420 48580 296476 48636
rect 296524 48580 296580 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 96636 47796 96692 47852
rect 96740 47796 96796 47852
rect 96844 47796 96900 47852
rect 127356 47796 127412 47852
rect 127460 47796 127516 47852
rect 127564 47796 127620 47852
rect 158076 47796 158132 47852
rect 158180 47796 158236 47852
rect 158284 47796 158340 47852
rect 188796 47796 188852 47852
rect 188900 47796 188956 47852
rect 189004 47796 189060 47852
rect 219516 47796 219572 47852
rect 219620 47796 219676 47852
rect 219724 47796 219780 47852
rect 250236 47796 250292 47852
rect 250340 47796 250396 47852
rect 250444 47796 250500 47852
rect 280956 47796 281012 47852
rect 281060 47796 281116 47852
rect 281164 47796 281220 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 81276 47012 81332 47068
rect 81380 47012 81436 47068
rect 81484 47012 81540 47068
rect 111996 47012 112052 47068
rect 112100 47012 112156 47068
rect 112204 47012 112260 47068
rect 142716 47012 142772 47068
rect 142820 47012 142876 47068
rect 142924 47012 142980 47068
rect 173436 47012 173492 47068
rect 173540 47012 173596 47068
rect 173644 47012 173700 47068
rect 204156 47012 204212 47068
rect 204260 47012 204316 47068
rect 204364 47012 204420 47068
rect 234876 47012 234932 47068
rect 234980 47012 235036 47068
rect 235084 47012 235140 47068
rect 265596 47012 265652 47068
rect 265700 47012 265756 47068
rect 265804 47012 265860 47068
rect 296316 47012 296372 47068
rect 296420 47012 296476 47068
rect 296524 47012 296580 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 96636 46228 96692 46284
rect 96740 46228 96796 46284
rect 96844 46228 96900 46284
rect 127356 46228 127412 46284
rect 127460 46228 127516 46284
rect 127564 46228 127620 46284
rect 158076 46228 158132 46284
rect 158180 46228 158236 46284
rect 158284 46228 158340 46284
rect 188796 46228 188852 46284
rect 188900 46228 188956 46284
rect 189004 46228 189060 46284
rect 219516 46228 219572 46284
rect 219620 46228 219676 46284
rect 219724 46228 219780 46284
rect 250236 46228 250292 46284
rect 250340 46228 250396 46284
rect 250444 46228 250500 46284
rect 280956 46228 281012 46284
rect 281060 46228 281116 46284
rect 281164 46228 281220 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 81276 45444 81332 45500
rect 81380 45444 81436 45500
rect 81484 45444 81540 45500
rect 111996 45444 112052 45500
rect 112100 45444 112156 45500
rect 112204 45444 112260 45500
rect 142716 45444 142772 45500
rect 142820 45444 142876 45500
rect 142924 45444 142980 45500
rect 173436 45444 173492 45500
rect 173540 45444 173596 45500
rect 173644 45444 173700 45500
rect 204156 45444 204212 45500
rect 204260 45444 204316 45500
rect 204364 45444 204420 45500
rect 234876 45444 234932 45500
rect 234980 45444 235036 45500
rect 235084 45444 235140 45500
rect 265596 45444 265652 45500
rect 265700 45444 265756 45500
rect 265804 45444 265860 45500
rect 296316 45444 296372 45500
rect 296420 45444 296476 45500
rect 296524 45444 296580 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 96636 44660 96692 44716
rect 96740 44660 96796 44716
rect 96844 44660 96900 44716
rect 127356 44660 127412 44716
rect 127460 44660 127516 44716
rect 127564 44660 127620 44716
rect 158076 44660 158132 44716
rect 158180 44660 158236 44716
rect 158284 44660 158340 44716
rect 188796 44660 188852 44716
rect 188900 44660 188956 44716
rect 189004 44660 189060 44716
rect 219516 44660 219572 44716
rect 219620 44660 219676 44716
rect 219724 44660 219780 44716
rect 250236 44660 250292 44716
rect 250340 44660 250396 44716
rect 250444 44660 250500 44716
rect 280956 44660 281012 44716
rect 281060 44660 281116 44716
rect 281164 44660 281220 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 81276 43876 81332 43932
rect 81380 43876 81436 43932
rect 81484 43876 81540 43932
rect 111996 43876 112052 43932
rect 112100 43876 112156 43932
rect 112204 43876 112260 43932
rect 142716 43876 142772 43932
rect 142820 43876 142876 43932
rect 142924 43876 142980 43932
rect 173436 43876 173492 43932
rect 173540 43876 173596 43932
rect 173644 43876 173700 43932
rect 204156 43876 204212 43932
rect 204260 43876 204316 43932
rect 204364 43876 204420 43932
rect 234876 43876 234932 43932
rect 234980 43876 235036 43932
rect 235084 43876 235140 43932
rect 265596 43876 265652 43932
rect 265700 43876 265756 43932
rect 265804 43876 265860 43932
rect 296316 43876 296372 43932
rect 296420 43876 296476 43932
rect 296524 43876 296580 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 96636 43092 96692 43148
rect 96740 43092 96796 43148
rect 96844 43092 96900 43148
rect 127356 43092 127412 43148
rect 127460 43092 127516 43148
rect 127564 43092 127620 43148
rect 158076 43092 158132 43148
rect 158180 43092 158236 43148
rect 158284 43092 158340 43148
rect 188796 43092 188852 43148
rect 188900 43092 188956 43148
rect 189004 43092 189060 43148
rect 219516 43092 219572 43148
rect 219620 43092 219676 43148
rect 219724 43092 219780 43148
rect 250236 43092 250292 43148
rect 250340 43092 250396 43148
rect 250444 43092 250500 43148
rect 280956 43092 281012 43148
rect 281060 43092 281116 43148
rect 281164 43092 281220 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 81276 42308 81332 42364
rect 81380 42308 81436 42364
rect 81484 42308 81540 42364
rect 111996 42308 112052 42364
rect 112100 42308 112156 42364
rect 112204 42308 112260 42364
rect 142716 42308 142772 42364
rect 142820 42308 142876 42364
rect 142924 42308 142980 42364
rect 173436 42308 173492 42364
rect 173540 42308 173596 42364
rect 173644 42308 173700 42364
rect 204156 42308 204212 42364
rect 204260 42308 204316 42364
rect 204364 42308 204420 42364
rect 234876 42308 234932 42364
rect 234980 42308 235036 42364
rect 235084 42308 235140 42364
rect 265596 42308 265652 42364
rect 265700 42308 265756 42364
rect 265804 42308 265860 42364
rect 296316 42308 296372 42364
rect 296420 42308 296476 42364
rect 296524 42308 296580 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 96636 41524 96692 41580
rect 96740 41524 96796 41580
rect 96844 41524 96900 41580
rect 127356 41524 127412 41580
rect 127460 41524 127516 41580
rect 127564 41524 127620 41580
rect 158076 41524 158132 41580
rect 158180 41524 158236 41580
rect 158284 41524 158340 41580
rect 188796 41524 188852 41580
rect 188900 41524 188956 41580
rect 189004 41524 189060 41580
rect 219516 41524 219572 41580
rect 219620 41524 219676 41580
rect 219724 41524 219780 41580
rect 250236 41524 250292 41580
rect 250340 41524 250396 41580
rect 250444 41524 250500 41580
rect 280956 41524 281012 41580
rect 281060 41524 281116 41580
rect 281164 41524 281220 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 81276 40740 81332 40796
rect 81380 40740 81436 40796
rect 81484 40740 81540 40796
rect 111996 40740 112052 40796
rect 112100 40740 112156 40796
rect 112204 40740 112260 40796
rect 142716 40740 142772 40796
rect 142820 40740 142876 40796
rect 142924 40740 142980 40796
rect 173436 40740 173492 40796
rect 173540 40740 173596 40796
rect 173644 40740 173700 40796
rect 204156 40740 204212 40796
rect 204260 40740 204316 40796
rect 204364 40740 204420 40796
rect 234876 40740 234932 40796
rect 234980 40740 235036 40796
rect 235084 40740 235140 40796
rect 265596 40740 265652 40796
rect 265700 40740 265756 40796
rect 265804 40740 265860 40796
rect 296316 40740 296372 40796
rect 296420 40740 296476 40796
rect 296524 40740 296580 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 96636 39956 96692 40012
rect 96740 39956 96796 40012
rect 96844 39956 96900 40012
rect 127356 39956 127412 40012
rect 127460 39956 127516 40012
rect 127564 39956 127620 40012
rect 158076 39956 158132 40012
rect 158180 39956 158236 40012
rect 158284 39956 158340 40012
rect 188796 39956 188852 40012
rect 188900 39956 188956 40012
rect 189004 39956 189060 40012
rect 219516 39956 219572 40012
rect 219620 39956 219676 40012
rect 219724 39956 219780 40012
rect 250236 39956 250292 40012
rect 250340 39956 250396 40012
rect 250444 39956 250500 40012
rect 280956 39956 281012 40012
rect 281060 39956 281116 40012
rect 281164 39956 281220 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 81276 39172 81332 39228
rect 81380 39172 81436 39228
rect 81484 39172 81540 39228
rect 111996 39172 112052 39228
rect 112100 39172 112156 39228
rect 112204 39172 112260 39228
rect 142716 39172 142772 39228
rect 142820 39172 142876 39228
rect 142924 39172 142980 39228
rect 173436 39172 173492 39228
rect 173540 39172 173596 39228
rect 173644 39172 173700 39228
rect 204156 39172 204212 39228
rect 204260 39172 204316 39228
rect 204364 39172 204420 39228
rect 234876 39172 234932 39228
rect 234980 39172 235036 39228
rect 235084 39172 235140 39228
rect 265596 39172 265652 39228
rect 265700 39172 265756 39228
rect 265804 39172 265860 39228
rect 296316 39172 296372 39228
rect 296420 39172 296476 39228
rect 296524 39172 296580 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 96636 38388 96692 38444
rect 96740 38388 96796 38444
rect 96844 38388 96900 38444
rect 127356 38388 127412 38444
rect 127460 38388 127516 38444
rect 127564 38388 127620 38444
rect 158076 38388 158132 38444
rect 158180 38388 158236 38444
rect 158284 38388 158340 38444
rect 188796 38388 188852 38444
rect 188900 38388 188956 38444
rect 189004 38388 189060 38444
rect 219516 38388 219572 38444
rect 219620 38388 219676 38444
rect 219724 38388 219780 38444
rect 250236 38388 250292 38444
rect 250340 38388 250396 38444
rect 250444 38388 250500 38444
rect 280956 38388 281012 38444
rect 281060 38388 281116 38444
rect 281164 38388 281220 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 81276 37604 81332 37660
rect 81380 37604 81436 37660
rect 81484 37604 81540 37660
rect 111996 37604 112052 37660
rect 112100 37604 112156 37660
rect 112204 37604 112260 37660
rect 142716 37604 142772 37660
rect 142820 37604 142876 37660
rect 142924 37604 142980 37660
rect 173436 37604 173492 37660
rect 173540 37604 173596 37660
rect 173644 37604 173700 37660
rect 204156 37604 204212 37660
rect 204260 37604 204316 37660
rect 204364 37604 204420 37660
rect 234876 37604 234932 37660
rect 234980 37604 235036 37660
rect 235084 37604 235140 37660
rect 265596 37604 265652 37660
rect 265700 37604 265756 37660
rect 265804 37604 265860 37660
rect 296316 37604 296372 37660
rect 296420 37604 296476 37660
rect 296524 37604 296580 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 96636 36820 96692 36876
rect 96740 36820 96796 36876
rect 96844 36820 96900 36876
rect 127356 36820 127412 36876
rect 127460 36820 127516 36876
rect 127564 36820 127620 36876
rect 158076 36820 158132 36876
rect 158180 36820 158236 36876
rect 158284 36820 158340 36876
rect 188796 36820 188852 36876
rect 188900 36820 188956 36876
rect 189004 36820 189060 36876
rect 219516 36820 219572 36876
rect 219620 36820 219676 36876
rect 219724 36820 219780 36876
rect 250236 36820 250292 36876
rect 250340 36820 250396 36876
rect 250444 36820 250500 36876
rect 280956 36820 281012 36876
rect 281060 36820 281116 36876
rect 281164 36820 281220 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 81276 36036 81332 36092
rect 81380 36036 81436 36092
rect 81484 36036 81540 36092
rect 111996 36036 112052 36092
rect 112100 36036 112156 36092
rect 112204 36036 112260 36092
rect 142716 36036 142772 36092
rect 142820 36036 142876 36092
rect 142924 36036 142980 36092
rect 173436 36036 173492 36092
rect 173540 36036 173596 36092
rect 173644 36036 173700 36092
rect 204156 36036 204212 36092
rect 204260 36036 204316 36092
rect 204364 36036 204420 36092
rect 234876 36036 234932 36092
rect 234980 36036 235036 36092
rect 235084 36036 235140 36092
rect 265596 36036 265652 36092
rect 265700 36036 265756 36092
rect 265804 36036 265860 36092
rect 296316 36036 296372 36092
rect 296420 36036 296476 36092
rect 296524 36036 296580 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 96636 35252 96692 35308
rect 96740 35252 96796 35308
rect 96844 35252 96900 35308
rect 127356 35252 127412 35308
rect 127460 35252 127516 35308
rect 127564 35252 127620 35308
rect 158076 35252 158132 35308
rect 158180 35252 158236 35308
rect 158284 35252 158340 35308
rect 188796 35252 188852 35308
rect 188900 35252 188956 35308
rect 189004 35252 189060 35308
rect 219516 35252 219572 35308
rect 219620 35252 219676 35308
rect 219724 35252 219780 35308
rect 250236 35252 250292 35308
rect 250340 35252 250396 35308
rect 250444 35252 250500 35308
rect 280956 35252 281012 35308
rect 281060 35252 281116 35308
rect 281164 35252 281220 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 81276 34468 81332 34524
rect 81380 34468 81436 34524
rect 81484 34468 81540 34524
rect 111996 34468 112052 34524
rect 112100 34468 112156 34524
rect 112204 34468 112260 34524
rect 142716 34468 142772 34524
rect 142820 34468 142876 34524
rect 142924 34468 142980 34524
rect 173436 34468 173492 34524
rect 173540 34468 173596 34524
rect 173644 34468 173700 34524
rect 204156 34468 204212 34524
rect 204260 34468 204316 34524
rect 204364 34468 204420 34524
rect 234876 34468 234932 34524
rect 234980 34468 235036 34524
rect 235084 34468 235140 34524
rect 265596 34468 265652 34524
rect 265700 34468 265756 34524
rect 265804 34468 265860 34524
rect 296316 34468 296372 34524
rect 296420 34468 296476 34524
rect 296524 34468 296580 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 96636 33684 96692 33740
rect 96740 33684 96796 33740
rect 96844 33684 96900 33740
rect 127356 33684 127412 33740
rect 127460 33684 127516 33740
rect 127564 33684 127620 33740
rect 158076 33684 158132 33740
rect 158180 33684 158236 33740
rect 158284 33684 158340 33740
rect 188796 33684 188852 33740
rect 188900 33684 188956 33740
rect 189004 33684 189060 33740
rect 219516 33684 219572 33740
rect 219620 33684 219676 33740
rect 219724 33684 219780 33740
rect 250236 33684 250292 33740
rect 250340 33684 250396 33740
rect 250444 33684 250500 33740
rect 280956 33684 281012 33740
rect 281060 33684 281116 33740
rect 281164 33684 281220 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 81276 32900 81332 32956
rect 81380 32900 81436 32956
rect 81484 32900 81540 32956
rect 111996 32900 112052 32956
rect 112100 32900 112156 32956
rect 112204 32900 112260 32956
rect 142716 32900 142772 32956
rect 142820 32900 142876 32956
rect 142924 32900 142980 32956
rect 173436 32900 173492 32956
rect 173540 32900 173596 32956
rect 173644 32900 173700 32956
rect 204156 32900 204212 32956
rect 204260 32900 204316 32956
rect 204364 32900 204420 32956
rect 234876 32900 234932 32956
rect 234980 32900 235036 32956
rect 235084 32900 235140 32956
rect 265596 32900 265652 32956
rect 265700 32900 265756 32956
rect 265804 32900 265860 32956
rect 296316 32900 296372 32956
rect 296420 32900 296476 32956
rect 296524 32900 296580 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 96636 32116 96692 32172
rect 96740 32116 96796 32172
rect 96844 32116 96900 32172
rect 127356 32116 127412 32172
rect 127460 32116 127516 32172
rect 127564 32116 127620 32172
rect 158076 32116 158132 32172
rect 158180 32116 158236 32172
rect 158284 32116 158340 32172
rect 188796 32116 188852 32172
rect 188900 32116 188956 32172
rect 189004 32116 189060 32172
rect 219516 32116 219572 32172
rect 219620 32116 219676 32172
rect 219724 32116 219780 32172
rect 250236 32116 250292 32172
rect 250340 32116 250396 32172
rect 250444 32116 250500 32172
rect 280956 32116 281012 32172
rect 281060 32116 281116 32172
rect 281164 32116 281220 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 81276 31332 81332 31388
rect 81380 31332 81436 31388
rect 81484 31332 81540 31388
rect 111996 31332 112052 31388
rect 112100 31332 112156 31388
rect 112204 31332 112260 31388
rect 142716 31332 142772 31388
rect 142820 31332 142876 31388
rect 142924 31332 142980 31388
rect 173436 31332 173492 31388
rect 173540 31332 173596 31388
rect 173644 31332 173700 31388
rect 204156 31332 204212 31388
rect 204260 31332 204316 31388
rect 204364 31332 204420 31388
rect 234876 31332 234932 31388
rect 234980 31332 235036 31388
rect 235084 31332 235140 31388
rect 265596 31332 265652 31388
rect 265700 31332 265756 31388
rect 265804 31332 265860 31388
rect 296316 31332 296372 31388
rect 296420 31332 296476 31388
rect 296524 31332 296580 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 96636 30548 96692 30604
rect 96740 30548 96796 30604
rect 96844 30548 96900 30604
rect 127356 30548 127412 30604
rect 127460 30548 127516 30604
rect 127564 30548 127620 30604
rect 158076 30548 158132 30604
rect 158180 30548 158236 30604
rect 158284 30548 158340 30604
rect 188796 30548 188852 30604
rect 188900 30548 188956 30604
rect 189004 30548 189060 30604
rect 219516 30548 219572 30604
rect 219620 30548 219676 30604
rect 219724 30548 219780 30604
rect 250236 30548 250292 30604
rect 250340 30548 250396 30604
rect 250444 30548 250500 30604
rect 280956 30548 281012 30604
rect 281060 30548 281116 30604
rect 281164 30548 281220 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 81276 29764 81332 29820
rect 81380 29764 81436 29820
rect 81484 29764 81540 29820
rect 111996 29764 112052 29820
rect 112100 29764 112156 29820
rect 112204 29764 112260 29820
rect 142716 29764 142772 29820
rect 142820 29764 142876 29820
rect 142924 29764 142980 29820
rect 173436 29764 173492 29820
rect 173540 29764 173596 29820
rect 173644 29764 173700 29820
rect 204156 29764 204212 29820
rect 204260 29764 204316 29820
rect 204364 29764 204420 29820
rect 234876 29764 234932 29820
rect 234980 29764 235036 29820
rect 235084 29764 235140 29820
rect 265596 29764 265652 29820
rect 265700 29764 265756 29820
rect 265804 29764 265860 29820
rect 296316 29764 296372 29820
rect 296420 29764 296476 29820
rect 296524 29764 296580 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 96636 28980 96692 29036
rect 96740 28980 96796 29036
rect 96844 28980 96900 29036
rect 127356 28980 127412 29036
rect 127460 28980 127516 29036
rect 127564 28980 127620 29036
rect 158076 28980 158132 29036
rect 158180 28980 158236 29036
rect 158284 28980 158340 29036
rect 188796 28980 188852 29036
rect 188900 28980 188956 29036
rect 189004 28980 189060 29036
rect 219516 28980 219572 29036
rect 219620 28980 219676 29036
rect 219724 28980 219780 29036
rect 250236 28980 250292 29036
rect 250340 28980 250396 29036
rect 250444 28980 250500 29036
rect 280956 28980 281012 29036
rect 281060 28980 281116 29036
rect 281164 28980 281220 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 81276 28196 81332 28252
rect 81380 28196 81436 28252
rect 81484 28196 81540 28252
rect 111996 28196 112052 28252
rect 112100 28196 112156 28252
rect 112204 28196 112260 28252
rect 142716 28196 142772 28252
rect 142820 28196 142876 28252
rect 142924 28196 142980 28252
rect 173436 28196 173492 28252
rect 173540 28196 173596 28252
rect 173644 28196 173700 28252
rect 204156 28196 204212 28252
rect 204260 28196 204316 28252
rect 204364 28196 204420 28252
rect 234876 28196 234932 28252
rect 234980 28196 235036 28252
rect 235084 28196 235140 28252
rect 265596 28196 265652 28252
rect 265700 28196 265756 28252
rect 265804 28196 265860 28252
rect 296316 28196 296372 28252
rect 296420 28196 296476 28252
rect 296524 28196 296580 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 96636 27412 96692 27468
rect 96740 27412 96796 27468
rect 96844 27412 96900 27468
rect 127356 27412 127412 27468
rect 127460 27412 127516 27468
rect 127564 27412 127620 27468
rect 158076 27412 158132 27468
rect 158180 27412 158236 27468
rect 158284 27412 158340 27468
rect 188796 27412 188852 27468
rect 188900 27412 188956 27468
rect 189004 27412 189060 27468
rect 219516 27412 219572 27468
rect 219620 27412 219676 27468
rect 219724 27412 219780 27468
rect 250236 27412 250292 27468
rect 250340 27412 250396 27468
rect 250444 27412 250500 27468
rect 280956 27412 281012 27468
rect 281060 27412 281116 27468
rect 281164 27412 281220 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 81276 26628 81332 26684
rect 81380 26628 81436 26684
rect 81484 26628 81540 26684
rect 111996 26628 112052 26684
rect 112100 26628 112156 26684
rect 112204 26628 112260 26684
rect 142716 26628 142772 26684
rect 142820 26628 142876 26684
rect 142924 26628 142980 26684
rect 173436 26628 173492 26684
rect 173540 26628 173596 26684
rect 173644 26628 173700 26684
rect 204156 26628 204212 26684
rect 204260 26628 204316 26684
rect 204364 26628 204420 26684
rect 234876 26628 234932 26684
rect 234980 26628 235036 26684
rect 235084 26628 235140 26684
rect 265596 26628 265652 26684
rect 265700 26628 265756 26684
rect 265804 26628 265860 26684
rect 296316 26628 296372 26684
rect 296420 26628 296476 26684
rect 296524 26628 296580 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 96636 25844 96692 25900
rect 96740 25844 96796 25900
rect 96844 25844 96900 25900
rect 127356 25844 127412 25900
rect 127460 25844 127516 25900
rect 127564 25844 127620 25900
rect 158076 25844 158132 25900
rect 158180 25844 158236 25900
rect 158284 25844 158340 25900
rect 188796 25844 188852 25900
rect 188900 25844 188956 25900
rect 189004 25844 189060 25900
rect 219516 25844 219572 25900
rect 219620 25844 219676 25900
rect 219724 25844 219780 25900
rect 250236 25844 250292 25900
rect 250340 25844 250396 25900
rect 250444 25844 250500 25900
rect 280956 25844 281012 25900
rect 281060 25844 281116 25900
rect 281164 25844 281220 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 81276 25060 81332 25116
rect 81380 25060 81436 25116
rect 81484 25060 81540 25116
rect 111996 25060 112052 25116
rect 112100 25060 112156 25116
rect 112204 25060 112260 25116
rect 142716 25060 142772 25116
rect 142820 25060 142876 25116
rect 142924 25060 142980 25116
rect 173436 25060 173492 25116
rect 173540 25060 173596 25116
rect 173644 25060 173700 25116
rect 204156 25060 204212 25116
rect 204260 25060 204316 25116
rect 204364 25060 204420 25116
rect 234876 25060 234932 25116
rect 234980 25060 235036 25116
rect 235084 25060 235140 25116
rect 265596 25060 265652 25116
rect 265700 25060 265756 25116
rect 265804 25060 265860 25116
rect 296316 25060 296372 25116
rect 296420 25060 296476 25116
rect 296524 25060 296580 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 96636 24276 96692 24332
rect 96740 24276 96796 24332
rect 96844 24276 96900 24332
rect 127356 24276 127412 24332
rect 127460 24276 127516 24332
rect 127564 24276 127620 24332
rect 158076 24276 158132 24332
rect 158180 24276 158236 24332
rect 158284 24276 158340 24332
rect 188796 24276 188852 24332
rect 188900 24276 188956 24332
rect 189004 24276 189060 24332
rect 219516 24276 219572 24332
rect 219620 24276 219676 24332
rect 219724 24276 219780 24332
rect 250236 24276 250292 24332
rect 250340 24276 250396 24332
rect 250444 24276 250500 24332
rect 280956 24276 281012 24332
rect 281060 24276 281116 24332
rect 281164 24276 281220 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 81276 23492 81332 23548
rect 81380 23492 81436 23548
rect 81484 23492 81540 23548
rect 111996 23492 112052 23548
rect 112100 23492 112156 23548
rect 112204 23492 112260 23548
rect 142716 23492 142772 23548
rect 142820 23492 142876 23548
rect 142924 23492 142980 23548
rect 173436 23492 173492 23548
rect 173540 23492 173596 23548
rect 173644 23492 173700 23548
rect 204156 23492 204212 23548
rect 204260 23492 204316 23548
rect 204364 23492 204420 23548
rect 234876 23492 234932 23548
rect 234980 23492 235036 23548
rect 235084 23492 235140 23548
rect 265596 23492 265652 23548
rect 265700 23492 265756 23548
rect 265804 23492 265860 23548
rect 296316 23492 296372 23548
rect 296420 23492 296476 23548
rect 296524 23492 296580 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 96636 22708 96692 22764
rect 96740 22708 96796 22764
rect 96844 22708 96900 22764
rect 127356 22708 127412 22764
rect 127460 22708 127516 22764
rect 127564 22708 127620 22764
rect 158076 22708 158132 22764
rect 158180 22708 158236 22764
rect 158284 22708 158340 22764
rect 188796 22708 188852 22764
rect 188900 22708 188956 22764
rect 189004 22708 189060 22764
rect 219516 22708 219572 22764
rect 219620 22708 219676 22764
rect 219724 22708 219780 22764
rect 250236 22708 250292 22764
rect 250340 22708 250396 22764
rect 250444 22708 250500 22764
rect 280956 22708 281012 22764
rect 281060 22708 281116 22764
rect 281164 22708 281220 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 81276 21924 81332 21980
rect 81380 21924 81436 21980
rect 81484 21924 81540 21980
rect 111996 21924 112052 21980
rect 112100 21924 112156 21980
rect 112204 21924 112260 21980
rect 142716 21924 142772 21980
rect 142820 21924 142876 21980
rect 142924 21924 142980 21980
rect 173436 21924 173492 21980
rect 173540 21924 173596 21980
rect 173644 21924 173700 21980
rect 204156 21924 204212 21980
rect 204260 21924 204316 21980
rect 204364 21924 204420 21980
rect 234876 21924 234932 21980
rect 234980 21924 235036 21980
rect 235084 21924 235140 21980
rect 265596 21924 265652 21980
rect 265700 21924 265756 21980
rect 265804 21924 265860 21980
rect 296316 21924 296372 21980
rect 296420 21924 296476 21980
rect 296524 21924 296580 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 96636 21140 96692 21196
rect 96740 21140 96796 21196
rect 96844 21140 96900 21196
rect 127356 21140 127412 21196
rect 127460 21140 127516 21196
rect 127564 21140 127620 21196
rect 158076 21140 158132 21196
rect 158180 21140 158236 21196
rect 158284 21140 158340 21196
rect 188796 21140 188852 21196
rect 188900 21140 188956 21196
rect 189004 21140 189060 21196
rect 219516 21140 219572 21196
rect 219620 21140 219676 21196
rect 219724 21140 219780 21196
rect 250236 21140 250292 21196
rect 250340 21140 250396 21196
rect 250444 21140 250500 21196
rect 280956 21140 281012 21196
rect 281060 21140 281116 21196
rect 281164 21140 281220 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 81276 20356 81332 20412
rect 81380 20356 81436 20412
rect 81484 20356 81540 20412
rect 111996 20356 112052 20412
rect 112100 20356 112156 20412
rect 112204 20356 112260 20412
rect 142716 20356 142772 20412
rect 142820 20356 142876 20412
rect 142924 20356 142980 20412
rect 173436 20356 173492 20412
rect 173540 20356 173596 20412
rect 173644 20356 173700 20412
rect 204156 20356 204212 20412
rect 204260 20356 204316 20412
rect 204364 20356 204420 20412
rect 234876 20356 234932 20412
rect 234980 20356 235036 20412
rect 235084 20356 235140 20412
rect 265596 20356 265652 20412
rect 265700 20356 265756 20412
rect 265804 20356 265860 20412
rect 296316 20356 296372 20412
rect 296420 20356 296476 20412
rect 296524 20356 296580 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 96636 19572 96692 19628
rect 96740 19572 96796 19628
rect 96844 19572 96900 19628
rect 127356 19572 127412 19628
rect 127460 19572 127516 19628
rect 127564 19572 127620 19628
rect 158076 19572 158132 19628
rect 158180 19572 158236 19628
rect 158284 19572 158340 19628
rect 188796 19572 188852 19628
rect 188900 19572 188956 19628
rect 189004 19572 189060 19628
rect 219516 19572 219572 19628
rect 219620 19572 219676 19628
rect 219724 19572 219780 19628
rect 250236 19572 250292 19628
rect 250340 19572 250396 19628
rect 250444 19572 250500 19628
rect 280956 19572 281012 19628
rect 281060 19572 281116 19628
rect 281164 19572 281220 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 81276 18788 81332 18844
rect 81380 18788 81436 18844
rect 81484 18788 81540 18844
rect 111996 18788 112052 18844
rect 112100 18788 112156 18844
rect 112204 18788 112260 18844
rect 142716 18788 142772 18844
rect 142820 18788 142876 18844
rect 142924 18788 142980 18844
rect 173436 18788 173492 18844
rect 173540 18788 173596 18844
rect 173644 18788 173700 18844
rect 204156 18788 204212 18844
rect 204260 18788 204316 18844
rect 204364 18788 204420 18844
rect 234876 18788 234932 18844
rect 234980 18788 235036 18844
rect 235084 18788 235140 18844
rect 265596 18788 265652 18844
rect 265700 18788 265756 18844
rect 265804 18788 265860 18844
rect 296316 18788 296372 18844
rect 296420 18788 296476 18844
rect 296524 18788 296580 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 96636 18004 96692 18060
rect 96740 18004 96796 18060
rect 96844 18004 96900 18060
rect 127356 18004 127412 18060
rect 127460 18004 127516 18060
rect 127564 18004 127620 18060
rect 158076 18004 158132 18060
rect 158180 18004 158236 18060
rect 158284 18004 158340 18060
rect 188796 18004 188852 18060
rect 188900 18004 188956 18060
rect 189004 18004 189060 18060
rect 219516 18004 219572 18060
rect 219620 18004 219676 18060
rect 219724 18004 219780 18060
rect 250236 18004 250292 18060
rect 250340 18004 250396 18060
rect 250444 18004 250500 18060
rect 280956 18004 281012 18060
rect 281060 18004 281116 18060
rect 281164 18004 281220 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 81276 17220 81332 17276
rect 81380 17220 81436 17276
rect 81484 17220 81540 17276
rect 111996 17220 112052 17276
rect 112100 17220 112156 17276
rect 112204 17220 112260 17276
rect 142716 17220 142772 17276
rect 142820 17220 142876 17276
rect 142924 17220 142980 17276
rect 173436 17220 173492 17276
rect 173540 17220 173596 17276
rect 173644 17220 173700 17276
rect 204156 17220 204212 17276
rect 204260 17220 204316 17276
rect 204364 17220 204420 17276
rect 234876 17220 234932 17276
rect 234980 17220 235036 17276
rect 235084 17220 235140 17276
rect 265596 17220 265652 17276
rect 265700 17220 265756 17276
rect 265804 17220 265860 17276
rect 296316 17220 296372 17276
rect 296420 17220 296476 17276
rect 296524 17220 296580 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 96636 16436 96692 16492
rect 96740 16436 96796 16492
rect 96844 16436 96900 16492
rect 127356 16436 127412 16492
rect 127460 16436 127516 16492
rect 127564 16436 127620 16492
rect 158076 16436 158132 16492
rect 158180 16436 158236 16492
rect 158284 16436 158340 16492
rect 188796 16436 188852 16492
rect 188900 16436 188956 16492
rect 189004 16436 189060 16492
rect 219516 16436 219572 16492
rect 219620 16436 219676 16492
rect 219724 16436 219780 16492
rect 250236 16436 250292 16492
rect 250340 16436 250396 16492
rect 250444 16436 250500 16492
rect 280956 16436 281012 16492
rect 281060 16436 281116 16492
rect 281164 16436 281220 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 81276 15652 81332 15708
rect 81380 15652 81436 15708
rect 81484 15652 81540 15708
rect 111996 15652 112052 15708
rect 112100 15652 112156 15708
rect 112204 15652 112260 15708
rect 142716 15652 142772 15708
rect 142820 15652 142876 15708
rect 142924 15652 142980 15708
rect 173436 15652 173492 15708
rect 173540 15652 173596 15708
rect 173644 15652 173700 15708
rect 204156 15652 204212 15708
rect 204260 15652 204316 15708
rect 204364 15652 204420 15708
rect 234876 15652 234932 15708
rect 234980 15652 235036 15708
rect 235084 15652 235140 15708
rect 265596 15652 265652 15708
rect 265700 15652 265756 15708
rect 265804 15652 265860 15708
rect 296316 15652 296372 15708
rect 296420 15652 296476 15708
rect 296524 15652 296580 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 96636 14868 96692 14924
rect 96740 14868 96796 14924
rect 96844 14868 96900 14924
rect 127356 14868 127412 14924
rect 127460 14868 127516 14924
rect 127564 14868 127620 14924
rect 158076 14868 158132 14924
rect 158180 14868 158236 14924
rect 158284 14868 158340 14924
rect 188796 14868 188852 14924
rect 188900 14868 188956 14924
rect 189004 14868 189060 14924
rect 219516 14868 219572 14924
rect 219620 14868 219676 14924
rect 219724 14868 219780 14924
rect 250236 14868 250292 14924
rect 250340 14868 250396 14924
rect 250444 14868 250500 14924
rect 280956 14868 281012 14924
rect 281060 14868 281116 14924
rect 281164 14868 281220 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 81276 14084 81332 14140
rect 81380 14084 81436 14140
rect 81484 14084 81540 14140
rect 111996 14084 112052 14140
rect 112100 14084 112156 14140
rect 112204 14084 112260 14140
rect 142716 14084 142772 14140
rect 142820 14084 142876 14140
rect 142924 14084 142980 14140
rect 173436 14084 173492 14140
rect 173540 14084 173596 14140
rect 173644 14084 173700 14140
rect 204156 14084 204212 14140
rect 204260 14084 204316 14140
rect 204364 14084 204420 14140
rect 234876 14084 234932 14140
rect 234980 14084 235036 14140
rect 235084 14084 235140 14140
rect 265596 14084 265652 14140
rect 265700 14084 265756 14140
rect 265804 14084 265860 14140
rect 296316 14084 296372 14140
rect 296420 14084 296476 14140
rect 296524 14084 296580 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 96636 13300 96692 13356
rect 96740 13300 96796 13356
rect 96844 13300 96900 13356
rect 127356 13300 127412 13356
rect 127460 13300 127516 13356
rect 127564 13300 127620 13356
rect 158076 13300 158132 13356
rect 158180 13300 158236 13356
rect 158284 13300 158340 13356
rect 188796 13300 188852 13356
rect 188900 13300 188956 13356
rect 189004 13300 189060 13356
rect 219516 13300 219572 13356
rect 219620 13300 219676 13356
rect 219724 13300 219780 13356
rect 250236 13300 250292 13356
rect 250340 13300 250396 13356
rect 250444 13300 250500 13356
rect 280956 13300 281012 13356
rect 281060 13300 281116 13356
rect 281164 13300 281220 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 81276 12516 81332 12572
rect 81380 12516 81436 12572
rect 81484 12516 81540 12572
rect 111996 12516 112052 12572
rect 112100 12516 112156 12572
rect 112204 12516 112260 12572
rect 142716 12516 142772 12572
rect 142820 12516 142876 12572
rect 142924 12516 142980 12572
rect 173436 12516 173492 12572
rect 173540 12516 173596 12572
rect 173644 12516 173700 12572
rect 204156 12516 204212 12572
rect 204260 12516 204316 12572
rect 204364 12516 204420 12572
rect 234876 12516 234932 12572
rect 234980 12516 235036 12572
rect 235084 12516 235140 12572
rect 265596 12516 265652 12572
rect 265700 12516 265756 12572
rect 265804 12516 265860 12572
rect 296316 12516 296372 12572
rect 296420 12516 296476 12572
rect 296524 12516 296580 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 96636 11732 96692 11788
rect 96740 11732 96796 11788
rect 96844 11732 96900 11788
rect 127356 11732 127412 11788
rect 127460 11732 127516 11788
rect 127564 11732 127620 11788
rect 158076 11732 158132 11788
rect 158180 11732 158236 11788
rect 158284 11732 158340 11788
rect 188796 11732 188852 11788
rect 188900 11732 188956 11788
rect 189004 11732 189060 11788
rect 219516 11732 219572 11788
rect 219620 11732 219676 11788
rect 219724 11732 219780 11788
rect 250236 11732 250292 11788
rect 250340 11732 250396 11788
rect 250444 11732 250500 11788
rect 280956 11732 281012 11788
rect 281060 11732 281116 11788
rect 281164 11732 281220 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 81276 10948 81332 11004
rect 81380 10948 81436 11004
rect 81484 10948 81540 11004
rect 111996 10948 112052 11004
rect 112100 10948 112156 11004
rect 112204 10948 112260 11004
rect 142716 10948 142772 11004
rect 142820 10948 142876 11004
rect 142924 10948 142980 11004
rect 173436 10948 173492 11004
rect 173540 10948 173596 11004
rect 173644 10948 173700 11004
rect 204156 10948 204212 11004
rect 204260 10948 204316 11004
rect 204364 10948 204420 11004
rect 234876 10948 234932 11004
rect 234980 10948 235036 11004
rect 235084 10948 235140 11004
rect 265596 10948 265652 11004
rect 265700 10948 265756 11004
rect 265804 10948 265860 11004
rect 296316 10948 296372 11004
rect 296420 10948 296476 11004
rect 296524 10948 296580 11004
rect 220780 10444 220836 10500
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 96636 10164 96692 10220
rect 96740 10164 96796 10220
rect 96844 10164 96900 10220
rect 127356 10164 127412 10220
rect 127460 10164 127516 10220
rect 127564 10164 127620 10220
rect 158076 10164 158132 10220
rect 158180 10164 158236 10220
rect 158284 10164 158340 10220
rect 188796 10164 188852 10220
rect 188900 10164 188956 10220
rect 189004 10164 189060 10220
rect 219516 10164 219572 10220
rect 219620 10164 219676 10220
rect 219724 10164 219780 10220
rect 250236 10164 250292 10220
rect 250340 10164 250396 10220
rect 250444 10164 250500 10220
rect 280956 10164 281012 10220
rect 281060 10164 281116 10220
rect 281164 10164 281220 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 81276 9380 81332 9436
rect 81380 9380 81436 9436
rect 81484 9380 81540 9436
rect 111996 9380 112052 9436
rect 112100 9380 112156 9436
rect 112204 9380 112260 9436
rect 142716 9380 142772 9436
rect 142820 9380 142876 9436
rect 142924 9380 142980 9436
rect 173436 9380 173492 9436
rect 173540 9380 173596 9436
rect 173644 9380 173700 9436
rect 204156 9380 204212 9436
rect 204260 9380 204316 9436
rect 204364 9380 204420 9436
rect 234876 9380 234932 9436
rect 234980 9380 235036 9436
rect 235084 9380 235140 9436
rect 265596 9380 265652 9436
rect 265700 9380 265756 9436
rect 265804 9380 265860 9436
rect 296316 9380 296372 9436
rect 296420 9380 296476 9436
rect 296524 9380 296580 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 96636 8596 96692 8652
rect 96740 8596 96796 8652
rect 96844 8596 96900 8652
rect 127356 8596 127412 8652
rect 127460 8596 127516 8652
rect 127564 8596 127620 8652
rect 158076 8596 158132 8652
rect 158180 8596 158236 8652
rect 158284 8596 158340 8652
rect 188796 8596 188852 8652
rect 188900 8596 188956 8652
rect 189004 8596 189060 8652
rect 219516 8596 219572 8652
rect 219620 8596 219676 8652
rect 219724 8596 219780 8652
rect 250236 8596 250292 8652
rect 250340 8596 250396 8652
rect 250444 8596 250500 8652
rect 280956 8596 281012 8652
rect 281060 8596 281116 8652
rect 281164 8596 281220 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 81276 7812 81332 7868
rect 81380 7812 81436 7868
rect 81484 7812 81540 7868
rect 111996 7812 112052 7868
rect 112100 7812 112156 7868
rect 112204 7812 112260 7868
rect 142716 7812 142772 7868
rect 142820 7812 142876 7868
rect 142924 7812 142980 7868
rect 173436 7812 173492 7868
rect 173540 7812 173596 7868
rect 173644 7812 173700 7868
rect 204156 7812 204212 7868
rect 204260 7812 204316 7868
rect 204364 7812 204420 7868
rect 234876 7812 234932 7868
rect 234980 7812 235036 7868
rect 235084 7812 235140 7868
rect 265596 7812 265652 7868
rect 265700 7812 265756 7868
rect 265804 7812 265860 7868
rect 296316 7812 296372 7868
rect 296420 7812 296476 7868
rect 296524 7812 296580 7868
rect 220780 7756 220836 7812
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 96636 7028 96692 7084
rect 96740 7028 96796 7084
rect 96844 7028 96900 7084
rect 127356 7028 127412 7084
rect 127460 7028 127516 7084
rect 127564 7028 127620 7084
rect 158076 7028 158132 7084
rect 158180 7028 158236 7084
rect 158284 7028 158340 7084
rect 188796 7028 188852 7084
rect 188900 7028 188956 7084
rect 189004 7028 189060 7084
rect 219516 7028 219572 7084
rect 219620 7028 219676 7084
rect 219724 7028 219780 7084
rect 250236 7028 250292 7084
rect 250340 7028 250396 7084
rect 250444 7028 250500 7084
rect 280956 7028 281012 7084
rect 281060 7028 281116 7084
rect 281164 7028 281220 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 81276 6244 81332 6300
rect 81380 6244 81436 6300
rect 81484 6244 81540 6300
rect 111996 6244 112052 6300
rect 112100 6244 112156 6300
rect 112204 6244 112260 6300
rect 142716 6244 142772 6300
rect 142820 6244 142876 6300
rect 142924 6244 142980 6300
rect 173436 6244 173492 6300
rect 173540 6244 173596 6300
rect 173644 6244 173700 6300
rect 204156 6244 204212 6300
rect 204260 6244 204316 6300
rect 204364 6244 204420 6300
rect 234876 6244 234932 6300
rect 234980 6244 235036 6300
rect 235084 6244 235140 6300
rect 265596 6244 265652 6300
rect 265700 6244 265756 6300
rect 265804 6244 265860 6300
rect 296316 6244 296372 6300
rect 296420 6244 296476 6300
rect 296524 6244 296580 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 96636 5460 96692 5516
rect 96740 5460 96796 5516
rect 96844 5460 96900 5516
rect 127356 5460 127412 5516
rect 127460 5460 127516 5516
rect 127564 5460 127620 5516
rect 158076 5460 158132 5516
rect 158180 5460 158236 5516
rect 158284 5460 158340 5516
rect 188796 5460 188852 5516
rect 188900 5460 188956 5516
rect 189004 5460 189060 5516
rect 219516 5460 219572 5516
rect 219620 5460 219676 5516
rect 219724 5460 219780 5516
rect 250236 5460 250292 5516
rect 250340 5460 250396 5516
rect 250444 5460 250500 5516
rect 280956 5460 281012 5516
rect 281060 5460 281116 5516
rect 281164 5460 281220 5516
rect 217084 4844 217140 4900
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 81276 4676 81332 4732
rect 81380 4676 81436 4732
rect 81484 4676 81540 4732
rect 111996 4676 112052 4732
rect 112100 4676 112156 4732
rect 112204 4676 112260 4732
rect 142716 4676 142772 4732
rect 142820 4676 142876 4732
rect 142924 4676 142980 4732
rect 173436 4676 173492 4732
rect 173540 4676 173596 4732
rect 173644 4676 173700 4732
rect 204156 4676 204212 4732
rect 204260 4676 204316 4732
rect 204364 4676 204420 4732
rect 234876 4676 234932 4732
rect 234980 4676 235036 4732
rect 235084 4676 235140 4732
rect 265596 4676 265652 4732
rect 265700 4676 265756 4732
rect 265804 4676 265860 4732
rect 296316 4676 296372 4732
rect 296420 4676 296476 4732
rect 296524 4676 296580 4732
rect 217084 4508 217140 4564
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 96636 3892 96692 3948
rect 96740 3892 96796 3948
rect 96844 3892 96900 3948
rect 127356 3892 127412 3948
rect 127460 3892 127516 3948
rect 127564 3892 127620 3948
rect 158076 3892 158132 3948
rect 158180 3892 158236 3948
rect 158284 3892 158340 3948
rect 188796 3892 188852 3948
rect 188900 3892 188956 3948
rect 189004 3892 189060 3948
rect 219516 3892 219572 3948
rect 219620 3892 219676 3948
rect 219724 3892 219780 3948
rect 250236 3892 250292 3948
rect 250340 3892 250396 3948
rect 250444 3892 250500 3948
rect 280956 3892 281012 3948
rect 281060 3892 281116 3948
rect 281164 3892 281220 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 81276 3108 81332 3164
rect 81380 3108 81436 3164
rect 81484 3108 81540 3164
rect 111996 3108 112052 3164
rect 112100 3108 112156 3164
rect 112204 3108 112260 3164
rect 142716 3108 142772 3164
rect 142820 3108 142876 3164
rect 142924 3108 142980 3164
rect 173436 3108 173492 3164
rect 173540 3108 173596 3164
rect 173644 3108 173700 3164
rect 204156 3108 204212 3164
rect 204260 3108 204316 3164
rect 204364 3108 204420 3164
rect 234876 3108 234932 3164
rect 234980 3108 235036 3164
rect 235084 3108 235140 3164
rect 265596 3108 265652 3164
rect 265700 3108 265756 3164
rect 265804 3108 265860 3164
rect 296316 3108 296372 3164
rect 296420 3108 296476 3164
rect 296524 3108 296580 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 55692 66208 56508
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
rect 81248 56476 81568 56508
rect 81248 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81568 56476
rect 81248 54908 81568 56420
rect 81248 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81568 54908
rect 81248 53340 81568 54852
rect 81248 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81568 53340
rect 81248 51772 81568 53284
rect 81248 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81568 51772
rect 81248 50204 81568 51716
rect 81248 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81568 50204
rect 81248 48636 81568 50148
rect 81248 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81568 48636
rect 81248 47068 81568 48580
rect 81248 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81568 47068
rect 81248 45500 81568 47012
rect 81248 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81568 45500
rect 81248 43932 81568 45444
rect 81248 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81568 43932
rect 81248 42364 81568 43876
rect 81248 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81568 42364
rect 81248 40796 81568 42308
rect 81248 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81568 40796
rect 81248 39228 81568 40740
rect 81248 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81568 39228
rect 81248 37660 81568 39172
rect 81248 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81568 37660
rect 81248 36092 81568 37604
rect 81248 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81568 36092
rect 81248 34524 81568 36036
rect 81248 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81568 34524
rect 81248 32956 81568 34468
rect 81248 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81568 32956
rect 81248 31388 81568 32900
rect 81248 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81568 31388
rect 81248 29820 81568 31332
rect 81248 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81568 29820
rect 81248 28252 81568 29764
rect 81248 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81568 28252
rect 81248 26684 81568 28196
rect 81248 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81568 26684
rect 81248 25116 81568 26628
rect 81248 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81568 25116
rect 81248 23548 81568 25060
rect 81248 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81568 23548
rect 81248 21980 81568 23492
rect 81248 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81568 21980
rect 81248 20412 81568 21924
rect 81248 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81568 20412
rect 81248 18844 81568 20356
rect 81248 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81568 18844
rect 81248 17276 81568 18788
rect 81248 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81568 17276
rect 81248 15708 81568 17220
rect 81248 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81568 15708
rect 81248 14140 81568 15652
rect 81248 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81568 14140
rect 81248 12572 81568 14084
rect 81248 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81568 12572
rect 81248 11004 81568 12516
rect 81248 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81568 11004
rect 81248 9436 81568 10948
rect 81248 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81568 9436
rect 81248 7868 81568 9380
rect 81248 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81568 7868
rect 81248 6300 81568 7812
rect 81248 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81568 6300
rect 81248 4732 81568 6244
rect 81248 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81568 4732
rect 81248 3164 81568 4676
rect 81248 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81568 3164
rect 81248 3076 81568 3108
rect 96608 55692 96928 56508
rect 96608 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96928 55692
rect 96608 54124 96928 55636
rect 96608 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96928 54124
rect 96608 52556 96928 54068
rect 96608 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96928 52556
rect 96608 50988 96928 52500
rect 96608 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96928 50988
rect 96608 49420 96928 50932
rect 96608 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96928 49420
rect 96608 47852 96928 49364
rect 96608 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96928 47852
rect 96608 46284 96928 47796
rect 96608 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96928 46284
rect 96608 44716 96928 46228
rect 96608 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96928 44716
rect 96608 43148 96928 44660
rect 96608 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96928 43148
rect 96608 41580 96928 43092
rect 96608 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96928 41580
rect 96608 40012 96928 41524
rect 96608 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96928 40012
rect 96608 38444 96928 39956
rect 96608 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96928 38444
rect 96608 36876 96928 38388
rect 96608 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96928 36876
rect 96608 35308 96928 36820
rect 96608 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96928 35308
rect 96608 33740 96928 35252
rect 96608 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96928 33740
rect 96608 32172 96928 33684
rect 96608 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96928 32172
rect 96608 30604 96928 32116
rect 96608 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96928 30604
rect 96608 29036 96928 30548
rect 96608 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96928 29036
rect 96608 27468 96928 28980
rect 96608 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96928 27468
rect 96608 25900 96928 27412
rect 96608 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96928 25900
rect 96608 24332 96928 25844
rect 96608 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96928 24332
rect 96608 22764 96928 24276
rect 96608 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96928 22764
rect 96608 21196 96928 22708
rect 96608 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96928 21196
rect 96608 19628 96928 21140
rect 96608 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96928 19628
rect 96608 18060 96928 19572
rect 96608 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96928 18060
rect 96608 16492 96928 18004
rect 96608 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96928 16492
rect 96608 14924 96928 16436
rect 96608 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96928 14924
rect 96608 13356 96928 14868
rect 96608 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96928 13356
rect 96608 11788 96928 13300
rect 96608 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96928 11788
rect 96608 10220 96928 11732
rect 96608 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96928 10220
rect 96608 8652 96928 10164
rect 96608 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96928 8652
rect 96608 7084 96928 8596
rect 96608 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96928 7084
rect 96608 5516 96928 7028
rect 96608 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96928 5516
rect 96608 3948 96928 5460
rect 96608 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96928 3948
rect 96608 3076 96928 3892
rect 111968 56476 112288 56508
rect 111968 56420 111996 56476
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 112260 56420 112288 56476
rect 111968 54908 112288 56420
rect 111968 54852 111996 54908
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 112260 54852 112288 54908
rect 111968 53340 112288 54852
rect 111968 53284 111996 53340
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 112260 53284 112288 53340
rect 111968 51772 112288 53284
rect 111968 51716 111996 51772
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 112260 51716 112288 51772
rect 111968 50204 112288 51716
rect 111968 50148 111996 50204
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 112260 50148 112288 50204
rect 111968 48636 112288 50148
rect 111968 48580 111996 48636
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 112260 48580 112288 48636
rect 111968 47068 112288 48580
rect 111968 47012 111996 47068
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 112260 47012 112288 47068
rect 111968 45500 112288 47012
rect 111968 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112288 45500
rect 111968 43932 112288 45444
rect 111968 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112288 43932
rect 111968 42364 112288 43876
rect 111968 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112288 42364
rect 111968 40796 112288 42308
rect 111968 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112288 40796
rect 111968 39228 112288 40740
rect 111968 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112288 39228
rect 111968 37660 112288 39172
rect 111968 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112288 37660
rect 111968 36092 112288 37604
rect 111968 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112288 36092
rect 111968 34524 112288 36036
rect 111968 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112288 34524
rect 111968 32956 112288 34468
rect 111968 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112288 32956
rect 111968 31388 112288 32900
rect 111968 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112288 31388
rect 111968 29820 112288 31332
rect 111968 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112288 29820
rect 111968 28252 112288 29764
rect 111968 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112288 28252
rect 111968 26684 112288 28196
rect 111968 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112288 26684
rect 111968 25116 112288 26628
rect 111968 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112288 25116
rect 111968 23548 112288 25060
rect 111968 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112288 23548
rect 111968 21980 112288 23492
rect 111968 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112288 21980
rect 111968 20412 112288 21924
rect 111968 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112288 20412
rect 111968 18844 112288 20356
rect 111968 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112288 18844
rect 111968 17276 112288 18788
rect 111968 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112288 17276
rect 111968 15708 112288 17220
rect 111968 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112288 15708
rect 111968 14140 112288 15652
rect 111968 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112288 14140
rect 111968 12572 112288 14084
rect 111968 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112288 12572
rect 111968 11004 112288 12516
rect 111968 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112288 11004
rect 111968 9436 112288 10948
rect 111968 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112288 9436
rect 111968 7868 112288 9380
rect 111968 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112288 7868
rect 111968 6300 112288 7812
rect 111968 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112288 6300
rect 111968 4732 112288 6244
rect 111968 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112288 4732
rect 111968 3164 112288 4676
rect 111968 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112288 3164
rect 111968 3076 112288 3108
rect 127328 55692 127648 56508
rect 127328 55636 127356 55692
rect 127412 55636 127460 55692
rect 127516 55636 127564 55692
rect 127620 55636 127648 55692
rect 127328 54124 127648 55636
rect 127328 54068 127356 54124
rect 127412 54068 127460 54124
rect 127516 54068 127564 54124
rect 127620 54068 127648 54124
rect 127328 52556 127648 54068
rect 127328 52500 127356 52556
rect 127412 52500 127460 52556
rect 127516 52500 127564 52556
rect 127620 52500 127648 52556
rect 127328 50988 127648 52500
rect 127328 50932 127356 50988
rect 127412 50932 127460 50988
rect 127516 50932 127564 50988
rect 127620 50932 127648 50988
rect 127328 49420 127648 50932
rect 127328 49364 127356 49420
rect 127412 49364 127460 49420
rect 127516 49364 127564 49420
rect 127620 49364 127648 49420
rect 127328 47852 127648 49364
rect 127328 47796 127356 47852
rect 127412 47796 127460 47852
rect 127516 47796 127564 47852
rect 127620 47796 127648 47852
rect 127328 46284 127648 47796
rect 127328 46228 127356 46284
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127620 46228 127648 46284
rect 127328 44716 127648 46228
rect 127328 44660 127356 44716
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127620 44660 127648 44716
rect 127328 43148 127648 44660
rect 127328 43092 127356 43148
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127620 43092 127648 43148
rect 127328 41580 127648 43092
rect 127328 41524 127356 41580
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127620 41524 127648 41580
rect 127328 40012 127648 41524
rect 127328 39956 127356 40012
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127620 39956 127648 40012
rect 127328 38444 127648 39956
rect 127328 38388 127356 38444
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127620 38388 127648 38444
rect 127328 36876 127648 38388
rect 127328 36820 127356 36876
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127620 36820 127648 36876
rect 127328 35308 127648 36820
rect 127328 35252 127356 35308
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127620 35252 127648 35308
rect 127328 33740 127648 35252
rect 127328 33684 127356 33740
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127620 33684 127648 33740
rect 127328 32172 127648 33684
rect 127328 32116 127356 32172
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127620 32116 127648 32172
rect 127328 30604 127648 32116
rect 127328 30548 127356 30604
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127620 30548 127648 30604
rect 127328 29036 127648 30548
rect 127328 28980 127356 29036
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127620 28980 127648 29036
rect 127328 27468 127648 28980
rect 127328 27412 127356 27468
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127620 27412 127648 27468
rect 127328 25900 127648 27412
rect 127328 25844 127356 25900
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127620 25844 127648 25900
rect 127328 24332 127648 25844
rect 127328 24276 127356 24332
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127620 24276 127648 24332
rect 127328 22764 127648 24276
rect 127328 22708 127356 22764
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127620 22708 127648 22764
rect 127328 21196 127648 22708
rect 127328 21140 127356 21196
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127620 21140 127648 21196
rect 127328 19628 127648 21140
rect 127328 19572 127356 19628
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127620 19572 127648 19628
rect 127328 18060 127648 19572
rect 127328 18004 127356 18060
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127620 18004 127648 18060
rect 127328 16492 127648 18004
rect 127328 16436 127356 16492
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127620 16436 127648 16492
rect 127328 14924 127648 16436
rect 127328 14868 127356 14924
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127620 14868 127648 14924
rect 127328 13356 127648 14868
rect 127328 13300 127356 13356
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127620 13300 127648 13356
rect 127328 11788 127648 13300
rect 127328 11732 127356 11788
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127620 11732 127648 11788
rect 127328 10220 127648 11732
rect 127328 10164 127356 10220
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127620 10164 127648 10220
rect 127328 8652 127648 10164
rect 127328 8596 127356 8652
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127620 8596 127648 8652
rect 127328 7084 127648 8596
rect 127328 7028 127356 7084
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127620 7028 127648 7084
rect 127328 5516 127648 7028
rect 127328 5460 127356 5516
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127620 5460 127648 5516
rect 127328 3948 127648 5460
rect 127328 3892 127356 3948
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127620 3892 127648 3948
rect 127328 3076 127648 3892
rect 142688 56476 143008 56508
rect 142688 56420 142716 56476
rect 142772 56420 142820 56476
rect 142876 56420 142924 56476
rect 142980 56420 143008 56476
rect 142688 54908 143008 56420
rect 142688 54852 142716 54908
rect 142772 54852 142820 54908
rect 142876 54852 142924 54908
rect 142980 54852 143008 54908
rect 142688 53340 143008 54852
rect 142688 53284 142716 53340
rect 142772 53284 142820 53340
rect 142876 53284 142924 53340
rect 142980 53284 143008 53340
rect 142688 51772 143008 53284
rect 142688 51716 142716 51772
rect 142772 51716 142820 51772
rect 142876 51716 142924 51772
rect 142980 51716 143008 51772
rect 142688 50204 143008 51716
rect 142688 50148 142716 50204
rect 142772 50148 142820 50204
rect 142876 50148 142924 50204
rect 142980 50148 143008 50204
rect 142688 48636 143008 50148
rect 142688 48580 142716 48636
rect 142772 48580 142820 48636
rect 142876 48580 142924 48636
rect 142980 48580 143008 48636
rect 142688 47068 143008 48580
rect 142688 47012 142716 47068
rect 142772 47012 142820 47068
rect 142876 47012 142924 47068
rect 142980 47012 143008 47068
rect 142688 45500 143008 47012
rect 142688 45444 142716 45500
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142980 45444 143008 45500
rect 142688 43932 143008 45444
rect 142688 43876 142716 43932
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142980 43876 143008 43932
rect 142688 42364 143008 43876
rect 142688 42308 142716 42364
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142980 42308 143008 42364
rect 142688 40796 143008 42308
rect 142688 40740 142716 40796
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142980 40740 143008 40796
rect 142688 39228 143008 40740
rect 142688 39172 142716 39228
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142980 39172 143008 39228
rect 142688 37660 143008 39172
rect 142688 37604 142716 37660
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142980 37604 143008 37660
rect 142688 36092 143008 37604
rect 142688 36036 142716 36092
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142980 36036 143008 36092
rect 142688 34524 143008 36036
rect 142688 34468 142716 34524
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142980 34468 143008 34524
rect 142688 32956 143008 34468
rect 142688 32900 142716 32956
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142980 32900 143008 32956
rect 142688 31388 143008 32900
rect 142688 31332 142716 31388
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142980 31332 143008 31388
rect 142688 29820 143008 31332
rect 142688 29764 142716 29820
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142980 29764 143008 29820
rect 142688 28252 143008 29764
rect 142688 28196 142716 28252
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142980 28196 143008 28252
rect 142688 26684 143008 28196
rect 142688 26628 142716 26684
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142980 26628 143008 26684
rect 142688 25116 143008 26628
rect 142688 25060 142716 25116
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142980 25060 143008 25116
rect 142688 23548 143008 25060
rect 142688 23492 142716 23548
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142980 23492 143008 23548
rect 142688 21980 143008 23492
rect 142688 21924 142716 21980
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142980 21924 143008 21980
rect 142688 20412 143008 21924
rect 142688 20356 142716 20412
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142980 20356 143008 20412
rect 142688 18844 143008 20356
rect 142688 18788 142716 18844
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142980 18788 143008 18844
rect 142688 17276 143008 18788
rect 142688 17220 142716 17276
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142980 17220 143008 17276
rect 142688 15708 143008 17220
rect 142688 15652 142716 15708
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142980 15652 143008 15708
rect 142688 14140 143008 15652
rect 142688 14084 142716 14140
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142980 14084 143008 14140
rect 142688 12572 143008 14084
rect 142688 12516 142716 12572
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142980 12516 143008 12572
rect 142688 11004 143008 12516
rect 142688 10948 142716 11004
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142980 10948 143008 11004
rect 142688 9436 143008 10948
rect 142688 9380 142716 9436
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142980 9380 143008 9436
rect 142688 7868 143008 9380
rect 142688 7812 142716 7868
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142980 7812 143008 7868
rect 142688 6300 143008 7812
rect 142688 6244 142716 6300
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142980 6244 143008 6300
rect 142688 4732 143008 6244
rect 142688 4676 142716 4732
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142980 4676 143008 4732
rect 142688 3164 143008 4676
rect 142688 3108 142716 3164
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142980 3108 143008 3164
rect 142688 3076 143008 3108
rect 158048 55692 158368 56508
rect 158048 55636 158076 55692
rect 158132 55636 158180 55692
rect 158236 55636 158284 55692
rect 158340 55636 158368 55692
rect 158048 54124 158368 55636
rect 158048 54068 158076 54124
rect 158132 54068 158180 54124
rect 158236 54068 158284 54124
rect 158340 54068 158368 54124
rect 158048 52556 158368 54068
rect 158048 52500 158076 52556
rect 158132 52500 158180 52556
rect 158236 52500 158284 52556
rect 158340 52500 158368 52556
rect 158048 50988 158368 52500
rect 158048 50932 158076 50988
rect 158132 50932 158180 50988
rect 158236 50932 158284 50988
rect 158340 50932 158368 50988
rect 158048 49420 158368 50932
rect 158048 49364 158076 49420
rect 158132 49364 158180 49420
rect 158236 49364 158284 49420
rect 158340 49364 158368 49420
rect 158048 47852 158368 49364
rect 158048 47796 158076 47852
rect 158132 47796 158180 47852
rect 158236 47796 158284 47852
rect 158340 47796 158368 47852
rect 158048 46284 158368 47796
rect 158048 46228 158076 46284
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158340 46228 158368 46284
rect 158048 44716 158368 46228
rect 158048 44660 158076 44716
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158340 44660 158368 44716
rect 158048 43148 158368 44660
rect 158048 43092 158076 43148
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158340 43092 158368 43148
rect 158048 41580 158368 43092
rect 158048 41524 158076 41580
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158340 41524 158368 41580
rect 158048 40012 158368 41524
rect 158048 39956 158076 40012
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158340 39956 158368 40012
rect 158048 38444 158368 39956
rect 158048 38388 158076 38444
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158340 38388 158368 38444
rect 158048 36876 158368 38388
rect 158048 36820 158076 36876
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158340 36820 158368 36876
rect 158048 35308 158368 36820
rect 158048 35252 158076 35308
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158340 35252 158368 35308
rect 158048 33740 158368 35252
rect 158048 33684 158076 33740
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158340 33684 158368 33740
rect 158048 32172 158368 33684
rect 158048 32116 158076 32172
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158340 32116 158368 32172
rect 158048 30604 158368 32116
rect 158048 30548 158076 30604
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158340 30548 158368 30604
rect 158048 29036 158368 30548
rect 158048 28980 158076 29036
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158340 28980 158368 29036
rect 158048 27468 158368 28980
rect 158048 27412 158076 27468
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158340 27412 158368 27468
rect 158048 25900 158368 27412
rect 158048 25844 158076 25900
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158340 25844 158368 25900
rect 158048 24332 158368 25844
rect 158048 24276 158076 24332
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158340 24276 158368 24332
rect 158048 22764 158368 24276
rect 158048 22708 158076 22764
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158340 22708 158368 22764
rect 158048 21196 158368 22708
rect 158048 21140 158076 21196
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158340 21140 158368 21196
rect 158048 19628 158368 21140
rect 158048 19572 158076 19628
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158340 19572 158368 19628
rect 158048 18060 158368 19572
rect 158048 18004 158076 18060
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158340 18004 158368 18060
rect 158048 16492 158368 18004
rect 158048 16436 158076 16492
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158340 16436 158368 16492
rect 158048 14924 158368 16436
rect 158048 14868 158076 14924
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158340 14868 158368 14924
rect 158048 13356 158368 14868
rect 158048 13300 158076 13356
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158340 13300 158368 13356
rect 158048 11788 158368 13300
rect 158048 11732 158076 11788
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158340 11732 158368 11788
rect 158048 10220 158368 11732
rect 158048 10164 158076 10220
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158340 10164 158368 10220
rect 158048 8652 158368 10164
rect 158048 8596 158076 8652
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158340 8596 158368 8652
rect 158048 7084 158368 8596
rect 158048 7028 158076 7084
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158340 7028 158368 7084
rect 158048 5516 158368 7028
rect 158048 5460 158076 5516
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158340 5460 158368 5516
rect 158048 3948 158368 5460
rect 158048 3892 158076 3948
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158340 3892 158368 3948
rect 158048 3076 158368 3892
rect 173408 56476 173728 56508
rect 173408 56420 173436 56476
rect 173492 56420 173540 56476
rect 173596 56420 173644 56476
rect 173700 56420 173728 56476
rect 173408 54908 173728 56420
rect 173408 54852 173436 54908
rect 173492 54852 173540 54908
rect 173596 54852 173644 54908
rect 173700 54852 173728 54908
rect 173408 53340 173728 54852
rect 173408 53284 173436 53340
rect 173492 53284 173540 53340
rect 173596 53284 173644 53340
rect 173700 53284 173728 53340
rect 173408 51772 173728 53284
rect 173408 51716 173436 51772
rect 173492 51716 173540 51772
rect 173596 51716 173644 51772
rect 173700 51716 173728 51772
rect 173408 50204 173728 51716
rect 173408 50148 173436 50204
rect 173492 50148 173540 50204
rect 173596 50148 173644 50204
rect 173700 50148 173728 50204
rect 173408 48636 173728 50148
rect 173408 48580 173436 48636
rect 173492 48580 173540 48636
rect 173596 48580 173644 48636
rect 173700 48580 173728 48636
rect 173408 47068 173728 48580
rect 173408 47012 173436 47068
rect 173492 47012 173540 47068
rect 173596 47012 173644 47068
rect 173700 47012 173728 47068
rect 173408 45500 173728 47012
rect 173408 45444 173436 45500
rect 173492 45444 173540 45500
rect 173596 45444 173644 45500
rect 173700 45444 173728 45500
rect 173408 43932 173728 45444
rect 173408 43876 173436 43932
rect 173492 43876 173540 43932
rect 173596 43876 173644 43932
rect 173700 43876 173728 43932
rect 173408 42364 173728 43876
rect 173408 42308 173436 42364
rect 173492 42308 173540 42364
rect 173596 42308 173644 42364
rect 173700 42308 173728 42364
rect 173408 40796 173728 42308
rect 173408 40740 173436 40796
rect 173492 40740 173540 40796
rect 173596 40740 173644 40796
rect 173700 40740 173728 40796
rect 173408 39228 173728 40740
rect 173408 39172 173436 39228
rect 173492 39172 173540 39228
rect 173596 39172 173644 39228
rect 173700 39172 173728 39228
rect 173408 37660 173728 39172
rect 173408 37604 173436 37660
rect 173492 37604 173540 37660
rect 173596 37604 173644 37660
rect 173700 37604 173728 37660
rect 173408 36092 173728 37604
rect 173408 36036 173436 36092
rect 173492 36036 173540 36092
rect 173596 36036 173644 36092
rect 173700 36036 173728 36092
rect 173408 34524 173728 36036
rect 173408 34468 173436 34524
rect 173492 34468 173540 34524
rect 173596 34468 173644 34524
rect 173700 34468 173728 34524
rect 173408 32956 173728 34468
rect 173408 32900 173436 32956
rect 173492 32900 173540 32956
rect 173596 32900 173644 32956
rect 173700 32900 173728 32956
rect 173408 31388 173728 32900
rect 173408 31332 173436 31388
rect 173492 31332 173540 31388
rect 173596 31332 173644 31388
rect 173700 31332 173728 31388
rect 173408 29820 173728 31332
rect 173408 29764 173436 29820
rect 173492 29764 173540 29820
rect 173596 29764 173644 29820
rect 173700 29764 173728 29820
rect 173408 28252 173728 29764
rect 173408 28196 173436 28252
rect 173492 28196 173540 28252
rect 173596 28196 173644 28252
rect 173700 28196 173728 28252
rect 173408 26684 173728 28196
rect 173408 26628 173436 26684
rect 173492 26628 173540 26684
rect 173596 26628 173644 26684
rect 173700 26628 173728 26684
rect 173408 25116 173728 26628
rect 173408 25060 173436 25116
rect 173492 25060 173540 25116
rect 173596 25060 173644 25116
rect 173700 25060 173728 25116
rect 173408 23548 173728 25060
rect 173408 23492 173436 23548
rect 173492 23492 173540 23548
rect 173596 23492 173644 23548
rect 173700 23492 173728 23548
rect 173408 21980 173728 23492
rect 173408 21924 173436 21980
rect 173492 21924 173540 21980
rect 173596 21924 173644 21980
rect 173700 21924 173728 21980
rect 173408 20412 173728 21924
rect 173408 20356 173436 20412
rect 173492 20356 173540 20412
rect 173596 20356 173644 20412
rect 173700 20356 173728 20412
rect 173408 18844 173728 20356
rect 173408 18788 173436 18844
rect 173492 18788 173540 18844
rect 173596 18788 173644 18844
rect 173700 18788 173728 18844
rect 173408 17276 173728 18788
rect 173408 17220 173436 17276
rect 173492 17220 173540 17276
rect 173596 17220 173644 17276
rect 173700 17220 173728 17276
rect 173408 15708 173728 17220
rect 173408 15652 173436 15708
rect 173492 15652 173540 15708
rect 173596 15652 173644 15708
rect 173700 15652 173728 15708
rect 173408 14140 173728 15652
rect 173408 14084 173436 14140
rect 173492 14084 173540 14140
rect 173596 14084 173644 14140
rect 173700 14084 173728 14140
rect 173408 12572 173728 14084
rect 173408 12516 173436 12572
rect 173492 12516 173540 12572
rect 173596 12516 173644 12572
rect 173700 12516 173728 12572
rect 173408 11004 173728 12516
rect 173408 10948 173436 11004
rect 173492 10948 173540 11004
rect 173596 10948 173644 11004
rect 173700 10948 173728 11004
rect 173408 9436 173728 10948
rect 173408 9380 173436 9436
rect 173492 9380 173540 9436
rect 173596 9380 173644 9436
rect 173700 9380 173728 9436
rect 173408 7868 173728 9380
rect 173408 7812 173436 7868
rect 173492 7812 173540 7868
rect 173596 7812 173644 7868
rect 173700 7812 173728 7868
rect 173408 6300 173728 7812
rect 173408 6244 173436 6300
rect 173492 6244 173540 6300
rect 173596 6244 173644 6300
rect 173700 6244 173728 6300
rect 173408 4732 173728 6244
rect 173408 4676 173436 4732
rect 173492 4676 173540 4732
rect 173596 4676 173644 4732
rect 173700 4676 173728 4732
rect 173408 3164 173728 4676
rect 173408 3108 173436 3164
rect 173492 3108 173540 3164
rect 173596 3108 173644 3164
rect 173700 3108 173728 3164
rect 173408 3076 173728 3108
rect 188768 55692 189088 56508
rect 188768 55636 188796 55692
rect 188852 55636 188900 55692
rect 188956 55636 189004 55692
rect 189060 55636 189088 55692
rect 188768 54124 189088 55636
rect 188768 54068 188796 54124
rect 188852 54068 188900 54124
rect 188956 54068 189004 54124
rect 189060 54068 189088 54124
rect 188768 52556 189088 54068
rect 188768 52500 188796 52556
rect 188852 52500 188900 52556
rect 188956 52500 189004 52556
rect 189060 52500 189088 52556
rect 188768 50988 189088 52500
rect 188768 50932 188796 50988
rect 188852 50932 188900 50988
rect 188956 50932 189004 50988
rect 189060 50932 189088 50988
rect 188768 49420 189088 50932
rect 188768 49364 188796 49420
rect 188852 49364 188900 49420
rect 188956 49364 189004 49420
rect 189060 49364 189088 49420
rect 188768 47852 189088 49364
rect 188768 47796 188796 47852
rect 188852 47796 188900 47852
rect 188956 47796 189004 47852
rect 189060 47796 189088 47852
rect 188768 46284 189088 47796
rect 188768 46228 188796 46284
rect 188852 46228 188900 46284
rect 188956 46228 189004 46284
rect 189060 46228 189088 46284
rect 188768 44716 189088 46228
rect 188768 44660 188796 44716
rect 188852 44660 188900 44716
rect 188956 44660 189004 44716
rect 189060 44660 189088 44716
rect 188768 43148 189088 44660
rect 188768 43092 188796 43148
rect 188852 43092 188900 43148
rect 188956 43092 189004 43148
rect 189060 43092 189088 43148
rect 188768 41580 189088 43092
rect 188768 41524 188796 41580
rect 188852 41524 188900 41580
rect 188956 41524 189004 41580
rect 189060 41524 189088 41580
rect 188768 40012 189088 41524
rect 188768 39956 188796 40012
rect 188852 39956 188900 40012
rect 188956 39956 189004 40012
rect 189060 39956 189088 40012
rect 188768 38444 189088 39956
rect 188768 38388 188796 38444
rect 188852 38388 188900 38444
rect 188956 38388 189004 38444
rect 189060 38388 189088 38444
rect 188768 36876 189088 38388
rect 188768 36820 188796 36876
rect 188852 36820 188900 36876
rect 188956 36820 189004 36876
rect 189060 36820 189088 36876
rect 188768 35308 189088 36820
rect 188768 35252 188796 35308
rect 188852 35252 188900 35308
rect 188956 35252 189004 35308
rect 189060 35252 189088 35308
rect 188768 33740 189088 35252
rect 188768 33684 188796 33740
rect 188852 33684 188900 33740
rect 188956 33684 189004 33740
rect 189060 33684 189088 33740
rect 188768 32172 189088 33684
rect 188768 32116 188796 32172
rect 188852 32116 188900 32172
rect 188956 32116 189004 32172
rect 189060 32116 189088 32172
rect 188768 30604 189088 32116
rect 188768 30548 188796 30604
rect 188852 30548 188900 30604
rect 188956 30548 189004 30604
rect 189060 30548 189088 30604
rect 188768 29036 189088 30548
rect 188768 28980 188796 29036
rect 188852 28980 188900 29036
rect 188956 28980 189004 29036
rect 189060 28980 189088 29036
rect 188768 27468 189088 28980
rect 188768 27412 188796 27468
rect 188852 27412 188900 27468
rect 188956 27412 189004 27468
rect 189060 27412 189088 27468
rect 188768 25900 189088 27412
rect 188768 25844 188796 25900
rect 188852 25844 188900 25900
rect 188956 25844 189004 25900
rect 189060 25844 189088 25900
rect 188768 24332 189088 25844
rect 188768 24276 188796 24332
rect 188852 24276 188900 24332
rect 188956 24276 189004 24332
rect 189060 24276 189088 24332
rect 188768 22764 189088 24276
rect 188768 22708 188796 22764
rect 188852 22708 188900 22764
rect 188956 22708 189004 22764
rect 189060 22708 189088 22764
rect 188768 21196 189088 22708
rect 188768 21140 188796 21196
rect 188852 21140 188900 21196
rect 188956 21140 189004 21196
rect 189060 21140 189088 21196
rect 188768 19628 189088 21140
rect 188768 19572 188796 19628
rect 188852 19572 188900 19628
rect 188956 19572 189004 19628
rect 189060 19572 189088 19628
rect 188768 18060 189088 19572
rect 188768 18004 188796 18060
rect 188852 18004 188900 18060
rect 188956 18004 189004 18060
rect 189060 18004 189088 18060
rect 188768 16492 189088 18004
rect 188768 16436 188796 16492
rect 188852 16436 188900 16492
rect 188956 16436 189004 16492
rect 189060 16436 189088 16492
rect 188768 14924 189088 16436
rect 188768 14868 188796 14924
rect 188852 14868 188900 14924
rect 188956 14868 189004 14924
rect 189060 14868 189088 14924
rect 188768 13356 189088 14868
rect 188768 13300 188796 13356
rect 188852 13300 188900 13356
rect 188956 13300 189004 13356
rect 189060 13300 189088 13356
rect 188768 11788 189088 13300
rect 188768 11732 188796 11788
rect 188852 11732 188900 11788
rect 188956 11732 189004 11788
rect 189060 11732 189088 11788
rect 188768 10220 189088 11732
rect 188768 10164 188796 10220
rect 188852 10164 188900 10220
rect 188956 10164 189004 10220
rect 189060 10164 189088 10220
rect 188768 8652 189088 10164
rect 188768 8596 188796 8652
rect 188852 8596 188900 8652
rect 188956 8596 189004 8652
rect 189060 8596 189088 8652
rect 188768 7084 189088 8596
rect 188768 7028 188796 7084
rect 188852 7028 188900 7084
rect 188956 7028 189004 7084
rect 189060 7028 189088 7084
rect 188768 5516 189088 7028
rect 188768 5460 188796 5516
rect 188852 5460 188900 5516
rect 188956 5460 189004 5516
rect 189060 5460 189088 5516
rect 188768 3948 189088 5460
rect 188768 3892 188796 3948
rect 188852 3892 188900 3948
rect 188956 3892 189004 3948
rect 189060 3892 189088 3948
rect 188768 3076 189088 3892
rect 204128 56476 204448 56508
rect 204128 56420 204156 56476
rect 204212 56420 204260 56476
rect 204316 56420 204364 56476
rect 204420 56420 204448 56476
rect 204128 54908 204448 56420
rect 204128 54852 204156 54908
rect 204212 54852 204260 54908
rect 204316 54852 204364 54908
rect 204420 54852 204448 54908
rect 204128 53340 204448 54852
rect 204128 53284 204156 53340
rect 204212 53284 204260 53340
rect 204316 53284 204364 53340
rect 204420 53284 204448 53340
rect 204128 51772 204448 53284
rect 204128 51716 204156 51772
rect 204212 51716 204260 51772
rect 204316 51716 204364 51772
rect 204420 51716 204448 51772
rect 204128 50204 204448 51716
rect 204128 50148 204156 50204
rect 204212 50148 204260 50204
rect 204316 50148 204364 50204
rect 204420 50148 204448 50204
rect 204128 48636 204448 50148
rect 204128 48580 204156 48636
rect 204212 48580 204260 48636
rect 204316 48580 204364 48636
rect 204420 48580 204448 48636
rect 204128 47068 204448 48580
rect 204128 47012 204156 47068
rect 204212 47012 204260 47068
rect 204316 47012 204364 47068
rect 204420 47012 204448 47068
rect 204128 45500 204448 47012
rect 204128 45444 204156 45500
rect 204212 45444 204260 45500
rect 204316 45444 204364 45500
rect 204420 45444 204448 45500
rect 204128 43932 204448 45444
rect 204128 43876 204156 43932
rect 204212 43876 204260 43932
rect 204316 43876 204364 43932
rect 204420 43876 204448 43932
rect 204128 42364 204448 43876
rect 204128 42308 204156 42364
rect 204212 42308 204260 42364
rect 204316 42308 204364 42364
rect 204420 42308 204448 42364
rect 204128 40796 204448 42308
rect 204128 40740 204156 40796
rect 204212 40740 204260 40796
rect 204316 40740 204364 40796
rect 204420 40740 204448 40796
rect 204128 39228 204448 40740
rect 204128 39172 204156 39228
rect 204212 39172 204260 39228
rect 204316 39172 204364 39228
rect 204420 39172 204448 39228
rect 204128 37660 204448 39172
rect 204128 37604 204156 37660
rect 204212 37604 204260 37660
rect 204316 37604 204364 37660
rect 204420 37604 204448 37660
rect 204128 36092 204448 37604
rect 204128 36036 204156 36092
rect 204212 36036 204260 36092
rect 204316 36036 204364 36092
rect 204420 36036 204448 36092
rect 204128 34524 204448 36036
rect 204128 34468 204156 34524
rect 204212 34468 204260 34524
rect 204316 34468 204364 34524
rect 204420 34468 204448 34524
rect 204128 32956 204448 34468
rect 204128 32900 204156 32956
rect 204212 32900 204260 32956
rect 204316 32900 204364 32956
rect 204420 32900 204448 32956
rect 204128 31388 204448 32900
rect 204128 31332 204156 31388
rect 204212 31332 204260 31388
rect 204316 31332 204364 31388
rect 204420 31332 204448 31388
rect 204128 29820 204448 31332
rect 204128 29764 204156 29820
rect 204212 29764 204260 29820
rect 204316 29764 204364 29820
rect 204420 29764 204448 29820
rect 204128 28252 204448 29764
rect 204128 28196 204156 28252
rect 204212 28196 204260 28252
rect 204316 28196 204364 28252
rect 204420 28196 204448 28252
rect 204128 26684 204448 28196
rect 204128 26628 204156 26684
rect 204212 26628 204260 26684
rect 204316 26628 204364 26684
rect 204420 26628 204448 26684
rect 204128 25116 204448 26628
rect 204128 25060 204156 25116
rect 204212 25060 204260 25116
rect 204316 25060 204364 25116
rect 204420 25060 204448 25116
rect 204128 23548 204448 25060
rect 204128 23492 204156 23548
rect 204212 23492 204260 23548
rect 204316 23492 204364 23548
rect 204420 23492 204448 23548
rect 204128 21980 204448 23492
rect 204128 21924 204156 21980
rect 204212 21924 204260 21980
rect 204316 21924 204364 21980
rect 204420 21924 204448 21980
rect 204128 20412 204448 21924
rect 204128 20356 204156 20412
rect 204212 20356 204260 20412
rect 204316 20356 204364 20412
rect 204420 20356 204448 20412
rect 204128 18844 204448 20356
rect 204128 18788 204156 18844
rect 204212 18788 204260 18844
rect 204316 18788 204364 18844
rect 204420 18788 204448 18844
rect 204128 17276 204448 18788
rect 204128 17220 204156 17276
rect 204212 17220 204260 17276
rect 204316 17220 204364 17276
rect 204420 17220 204448 17276
rect 204128 15708 204448 17220
rect 204128 15652 204156 15708
rect 204212 15652 204260 15708
rect 204316 15652 204364 15708
rect 204420 15652 204448 15708
rect 204128 14140 204448 15652
rect 204128 14084 204156 14140
rect 204212 14084 204260 14140
rect 204316 14084 204364 14140
rect 204420 14084 204448 14140
rect 204128 12572 204448 14084
rect 204128 12516 204156 12572
rect 204212 12516 204260 12572
rect 204316 12516 204364 12572
rect 204420 12516 204448 12572
rect 204128 11004 204448 12516
rect 204128 10948 204156 11004
rect 204212 10948 204260 11004
rect 204316 10948 204364 11004
rect 204420 10948 204448 11004
rect 204128 9436 204448 10948
rect 204128 9380 204156 9436
rect 204212 9380 204260 9436
rect 204316 9380 204364 9436
rect 204420 9380 204448 9436
rect 204128 7868 204448 9380
rect 204128 7812 204156 7868
rect 204212 7812 204260 7868
rect 204316 7812 204364 7868
rect 204420 7812 204448 7868
rect 204128 6300 204448 7812
rect 204128 6244 204156 6300
rect 204212 6244 204260 6300
rect 204316 6244 204364 6300
rect 204420 6244 204448 6300
rect 204128 4732 204448 6244
rect 219488 55692 219808 56508
rect 219488 55636 219516 55692
rect 219572 55636 219620 55692
rect 219676 55636 219724 55692
rect 219780 55636 219808 55692
rect 219488 54124 219808 55636
rect 219488 54068 219516 54124
rect 219572 54068 219620 54124
rect 219676 54068 219724 54124
rect 219780 54068 219808 54124
rect 219488 52556 219808 54068
rect 219488 52500 219516 52556
rect 219572 52500 219620 52556
rect 219676 52500 219724 52556
rect 219780 52500 219808 52556
rect 219488 50988 219808 52500
rect 219488 50932 219516 50988
rect 219572 50932 219620 50988
rect 219676 50932 219724 50988
rect 219780 50932 219808 50988
rect 219488 49420 219808 50932
rect 219488 49364 219516 49420
rect 219572 49364 219620 49420
rect 219676 49364 219724 49420
rect 219780 49364 219808 49420
rect 219488 47852 219808 49364
rect 219488 47796 219516 47852
rect 219572 47796 219620 47852
rect 219676 47796 219724 47852
rect 219780 47796 219808 47852
rect 219488 46284 219808 47796
rect 219488 46228 219516 46284
rect 219572 46228 219620 46284
rect 219676 46228 219724 46284
rect 219780 46228 219808 46284
rect 219488 44716 219808 46228
rect 219488 44660 219516 44716
rect 219572 44660 219620 44716
rect 219676 44660 219724 44716
rect 219780 44660 219808 44716
rect 219488 43148 219808 44660
rect 219488 43092 219516 43148
rect 219572 43092 219620 43148
rect 219676 43092 219724 43148
rect 219780 43092 219808 43148
rect 219488 41580 219808 43092
rect 219488 41524 219516 41580
rect 219572 41524 219620 41580
rect 219676 41524 219724 41580
rect 219780 41524 219808 41580
rect 219488 40012 219808 41524
rect 219488 39956 219516 40012
rect 219572 39956 219620 40012
rect 219676 39956 219724 40012
rect 219780 39956 219808 40012
rect 219488 38444 219808 39956
rect 219488 38388 219516 38444
rect 219572 38388 219620 38444
rect 219676 38388 219724 38444
rect 219780 38388 219808 38444
rect 219488 36876 219808 38388
rect 219488 36820 219516 36876
rect 219572 36820 219620 36876
rect 219676 36820 219724 36876
rect 219780 36820 219808 36876
rect 219488 35308 219808 36820
rect 219488 35252 219516 35308
rect 219572 35252 219620 35308
rect 219676 35252 219724 35308
rect 219780 35252 219808 35308
rect 219488 33740 219808 35252
rect 219488 33684 219516 33740
rect 219572 33684 219620 33740
rect 219676 33684 219724 33740
rect 219780 33684 219808 33740
rect 219488 32172 219808 33684
rect 219488 32116 219516 32172
rect 219572 32116 219620 32172
rect 219676 32116 219724 32172
rect 219780 32116 219808 32172
rect 219488 30604 219808 32116
rect 219488 30548 219516 30604
rect 219572 30548 219620 30604
rect 219676 30548 219724 30604
rect 219780 30548 219808 30604
rect 219488 29036 219808 30548
rect 219488 28980 219516 29036
rect 219572 28980 219620 29036
rect 219676 28980 219724 29036
rect 219780 28980 219808 29036
rect 219488 27468 219808 28980
rect 219488 27412 219516 27468
rect 219572 27412 219620 27468
rect 219676 27412 219724 27468
rect 219780 27412 219808 27468
rect 219488 25900 219808 27412
rect 219488 25844 219516 25900
rect 219572 25844 219620 25900
rect 219676 25844 219724 25900
rect 219780 25844 219808 25900
rect 219488 24332 219808 25844
rect 219488 24276 219516 24332
rect 219572 24276 219620 24332
rect 219676 24276 219724 24332
rect 219780 24276 219808 24332
rect 219488 22764 219808 24276
rect 219488 22708 219516 22764
rect 219572 22708 219620 22764
rect 219676 22708 219724 22764
rect 219780 22708 219808 22764
rect 219488 21196 219808 22708
rect 219488 21140 219516 21196
rect 219572 21140 219620 21196
rect 219676 21140 219724 21196
rect 219780 21140 219808 21196
rect 219488 19628 219808 21140
rect 219488 19572 219516 19628
rect 219572 19572 219620 19628
rect 219676 19572 219724 19628
rect 219780 19572 219808 19628
rect 219488 18060 219808 19572
rect 219488 18004 219516 18060
rect 219572 18004 219620 18060
rect 219676 18004 219724 18060
rect 219780 18004 219808 18060
rect 219488 16492 219808 18004
rect 219488 16436 219516 16492
rect 219572 16436 219620 16492
rect 219676 16436 219724 16492
rect 219780 16436 219808 16492
rect 219488 14924 219808 16436
rect 219488 14868 219516 14924
rect 219572 14868 219620 14924
rect 219676 14868 219724 14924
rect 219780 14868 219808 14924
rect 219488 13356 219808 14868
rect 219488 13300 219516 13356
rect 219572 13300 219620 13356
rect 219676 13300 219724 13356
rect 219780 13300 219808 13356
rect 219488 11788 219808 13300
rect 219488 11732 219516 11788
rect 219572 11732 219620 11788
rect 219676 11732 219724 11788
rect 219780 11732 219808 11788
rect 219488 10220 219808 11732
rect 234848 56476 235168 56508
rect 234848 56420 234876 56476
rect 234932 56420 234980 56476
rect 235036 56420 235084 56476
rect 235140 56420 235168 56476
rect 234848 54908 235168 56420
rect 234848 54852 234876 54908
rect 234932 54852 234980 54908
rect 235036 54852 235084 54908
rect 235140 54852 235168 54908
rect 234848 53340 235168 54852
rect 234848 53284 234876 53340
rect 234932 53284 234980 53340
rect 235036 53284 235084 53340
rect 235140 53284 235168 53340
rect 234848 51772 235168 53284
rect 234848 51716 234876 51772
rect 234932 51716 234980 51772
rect 235036 51716 235084 51772
rect 235140 51716 235168 51772
rect 234848 50204 235168 51716
rect 234848 50148 234876 50204
rect 234932 50148 234980 50204
rect 235036 50148 235084 50204
rect 235140 50148 235168 50204
rect 234848 48636 235168 50148
rect 234848 48580 234876 48636
rect 234932 48580 234980 48636
rect 235036 48580 235084 48636
rect 235140 48580 235168 48636
rect 234848 47068 235168 48580
rect 234848 47012 234876 47068
rect 234932 47012 234980 47068
rect 235036 47012 235084 47068
rect 235140 47012 235168 47068
rect 234848 45500 235168 47012
rect 234848 45444 234876 45500
rect 234932 45444 234980 45500
rect 235036 45444 235084 45500
rect 235140 45444 235168 45500
rect 234848 43932 235168 45444
rect 234848 43876 234876 43932
rect 234932 43876 234980 43932
rect 235036 43876 235084 43932
rect 235140 43876 235168 43932
rect 234848 42364 235168 43876
rect 234848 42308 234876 42364
rect 234932 42308 234980 42364
rect 235036 42308 235084 42364
rect 235140 42308 235168 42364
rect 234848 40796 235168 42308
rect 234848 40740 234876 40796
rect 234932 40740 234980 40796
rect 235036 40740 235084 40796
rect 235140 40740 235168 40796
rect 234848 39228 235168 40740
rect 234848 39172 234876 39228
rect 234932 39172 234980 39228
rect 235036 39172 235084 39228
rect 235140 39172 235168 39228
rect 234848 37660 235168 39172
rect 234848 37604 234876 37660
rect 234932 37604 234980 37660
rect 235036 37604 235084 37660
rect 235140 37604 235168 37660
rect 234848 36092 235168 37604
rect 234848 36036 234876 36092
rect 234932 36036 234980 36092
rect 235036 36036 235084 36092
rect 235140 36036 235168 36092
rect 234848 34524 235168 36036
rect 234848 34468 234876 34524
rect 234932 34468 234980 34524
rect 235036 34468 235084 34524
rect 235140 34468 235168 34524
rect 234848 32956 235168 34468
rect 234848 32900 234876 32956
rect 234932 32900 234980 32956
rect 235036 32900 235084 32956
rect 235140 32900 235168 32956
rect 234848 31388 235168 32900
rect 234848 31332 234876 31388
rect 234932 31332 234980 31388
rect 235036 31332 235084 31388
rect 235140 31332 235168 31388
rect 234848 29820 235168 31332
rect 234848 29764 234876 29820
rect 234932 29764 234980 29820
rect 235036 29764 235084 29820
rect 235140 29764 235168 29820
rect 234848 28252 235168 29764
rect 234848 28196 234876 28252
rect 234932 28196 234980 28252
rect 235036 28196 235084 28252
rect 235140 28196 235168 28252
rect 234848 26684 235168 28196
rect 234848 26628 234876 26684
rect 234932 26628 234980 26684
rect 235036 26628 235084 26684
rect 235140 26628 235168 26684
rect 234848 25116 235168 26628
rect 234848 25060 234876 25116
rect 234932 25060 234980 25116
rect 235036 25060 235084 25116
rect 235140 25060 235168 25116
rect 234848 23548 235168 25060
rect 234848 23492 234876 23548
rect 234932 23492 234980 23548
rect 235036 23492 235084 23548
rect 235140 23492 235168 23548
rect 234848 21980 235168 23492
rect 234848 21924 234876 21980
rect 234932 21924 234980 21980
rect 235036 21924 235084 21980
rect 235140 21924 235168 21980
rect 234848 20412 235168 21924
rect 234848 20356 234876 20412
rect 234932 20356 234980 20412
rect 235036 20356 235084 20412
rect 235140 20356 235168 20412
rect 234848 18844 235168 20356
rect 234848 18788 234876 18844
rect 234932 18788 234980 18844
rect 235036 18788 235084 18844
rect 235140 18788 235168 18844
rect 234848 17276 235168 18788
rect 234848 17220 234876 17276
rect 234932 17220 234980 17276
rect 235036 17220 235084 17276
rect 235140 17220 235168 17276
rect 234848 15708 235168 17220
rect 234848 15652 234876 15708
rect 234932 15652 234980 15708
rect 235036 15652 235084 15708
rect 235140 15652 235168 15708
rect 234848 14140 235168 15652
rect 234848 14084 234876 14140
rect 234932 14084 234980 14140
rect 235036 14084 235084 14140
rect 235140 14084 235168 14140
rect 234848 12572 235168 14084
rect 234848 12516 234876 12572
rect 234932 12516 234980 12572
rect 235036 12516 235084 12572
rect 235140 12516 235168 12572
rect 234848 11004 235168 12516
rect 234848 10948 234876 11004
rect 234932 10948 234980 11004
rect 235036 10948 235084 11004
rect 235140 10948 235168 11004
rect 219488 10164 219516 10220
rect 219572 10164 219620 10220
rect 219676 10164 219724 10220
rect 219780 10164 219808 10220
rect 219488 8652 219808 10164
rect 219488 8596 219516 8652
rect 219572 8596 219620 8652
rect 219676 8596 219724 8652
rect 219780 8596 219808 8652
rect 219488 7084 219808 8596
rect 220780 10500 220836 10510
rect 220780 7812 220836 10444
rect 220780 7746 220836 7756
rect 234848 9436 235168 10948
rect 234848 9380 234876 9436
rect 234932 9380 234980 9436
rect 235036 9380 235084 9436
rect 235140 9380 235168 9436
rect 234848 7868 235168 9380
rect 234848 7812 234876 7868
rect 234932 7812 234980 7868
rect 235036 7812 235084 7868
rect 235140 7812 235168 7868
rect 219488 7028 219516 7084
rect 219572 7028 219620 7084
rect 219676 7028 219724 7084
rect 219780 7028 219808 7084
rect 219488 5516 219808 7028
rect 219488 5460 219516 5516
rect 219572 5460 219620 5516
rect 219676 5460 219724 5516
rect 219780 5460 219808 5516
rect 204128 4676 204156 4732
rect 204212 4676 204260 4732
rect 204316 4676 204364 4732
rect 204420 4676 204448 4732
rect 204128 3164 204448 4676
rect 217084 4900 217140 4910
rect 217084 4564 217140 4844
rect 217084 4498 217140 4508
rect 204128 3108 204156 3164
rect 204212 3108 204260 3164
rect 204316 3108 204364 3164
rect 204420 3108 204448 3164
rect 204128 3076 204448 3108
rect 219488 3948 219808 5460
rect 219488 3892 219516 3948
rect 219572 3892 219620 3948
rect 219676 3892 219724 3948
rect 219780 3892 219808 3948
rect 219488 3076 219808 3892
rect 234848 6300 235168 7812
rect 234848 6244 234876 6300
rect 234932 6244 234980 6300
rect 235036 6244 235084 6300
rect 235140 6244 235168 6300
rect 234848 4732 235168 6244
rect 234848 4676 234876 4732
rect 234932 4676 234980 4732
rect 235036 4676 235084 4732
rect 235140 4676 235168 4732
rect 234848 3164 235168 4676
rect 234848 3108 234876 3164
rect 234932 3108 234980 3164
rect 235036 3108 235084 3164
rect 235140 3108 235168 3164
rect 234848 3076 235168 3108
rect 250208 55692 250528 56508
rect 250208 55636 250236 55692
rect 250292 55636 250340 55692
rect 250396 55636 250444 55692
rect 250500 55636 250528 55692
rect 250208 54124 250528 55636
rect 250208 54068 250236 54124
rect 250292 54068 250340 54124
rect 250396 54068 250444 54124
rect 250500 54068 250528 54124
rect 250208 52556 250528 54068
rect 250208 52500 250236 52556
rect 250292 52500 250340 52556
rect 250396 52500 250444 52556
rect 250500 52500 250528 52556
rect 250208 50988 250528 52500
rect 250208 50932 250236 50988
rect 250292 50932 250340 50988
rect 250396 50932 250444 50988
rect 250500 50932 250528 50988
rect 250208 49420 250528 50932
rect 250208 49364 250236 49420
rect 250292 49364 250340 49420
rect 250396 49364 250444 49420
rect 250500 49364 250528 49420
rect 250208 47852 250528 49364
rect 250208 47796 250236 47852
rect 250292 47796 250340 47852
rect 250396 47796 250444 47852
rect 250500 47796 250528 47852
rect 250208 46284 250528 47796
rect 250208 46228 250236 46284
rect 250292 46228 250340 46284
rect 250396 46228 250444 46284
rect 250500 46228 250528 46284
rect 250208 44716 250528 46228
rect 250208 44660 250236 44716
rect 250292 44660 250340 44716
rect 250396 44660 250444 44716
rect 250500 44660 250528 44716
rect 250208 43148 250528 44660
rect 250208 43092 250236 43148
rect 250292 43092 250340 43148
rect 250396 43092 250444 43148
rect 250500 43092 250528 43148
rect 250208 41580 250528 43092
rect 250208 41524 250236 41580
rect 250292 41524 250340 41580
rect 250396 41524 250444 41580
rect 250500 41524 250528 41580
rect 250208 40012 250528 41524
rect 250208 39956 250236 40012
rect 250292 39956 250340 40012
rect 250396 39956 250444 40012
rect 250500 39956 250528 40012
rect 250208 38444 250528 39956
rect 250208 38388 250236 38444
rect 250292 38388 250340 38444
rect 250396 38388 250444 38444
rect 250500 38388 250528 38444
rect 250208 36876 250528 38388
rect 250208 36820 250236 36876
rect 250292 36820 250340 36876
rect 250396 36820 250444 36876
rect 250500 36820 250528 36876
rect 250208 35308 250528 36820
rect 250208 35252 250236 35308
rect 250292 35252 250340 35308
rect 250396 35252 250444 35308
rect 250500 35252 250528 35308
rect 250208 33740 250528 35252
rect 250208 33684 250236 33740
rect 250292 33684 250340 33740
rect 250396 33684 250444 33740
rect 250500 33684 250528 33740
rect 250208 32172 250528 33684
rect 250208 32116 250236 32172
rect 250292 32116 250340 32172
rect 250396 32116 250444 32172
rect 250500 32116 250528 32172
rect 250208 30604 250528 32116
rect 250208 30548 250236 30604
rect 250292 30548 250340 30604
rect 250396 30548 250444 30604
rect 250500 30548 250528 30604
rect 250208 29036 250528 30548
rect 250208 28980 250236 29036
rect 250292 28980 250340 29036
rect 250396 28980 250444 29036
rect 250500 28980 250528 29036
rect 250208 27468 250528 28980
rect 250208 27412 250236 27468
rect 250292 27412 250340 27468
rect 250396 27412 250444 27468
rect 250500 27412 250528 27468
rect 250208 25900 250528 27412
rect 250208 25844 250236 25900
rect 250292 25844 250340 25900
rect 250396 25844 250444 25900
rect 250500 25844 250528 25900
rect 250208 24332 250528 25844
rect 250208 24276 250236 24332
rect 250292 24276 250340 24332
rect 250396 24276 250444 24332
rect 250500 24276 250528 24332
rect 250208 22764 250528 24276
rect 250208 22708 250236 22764
rect 250292 22708 250340 22764
rect 250396 22708 250444 22764
rect 250500 22708 250528 22764
rect 250208 21196 250528 22708
rect 250208 21140 250236 21196
rect 250292 21140 250340 21196
rect 250396 21140 250444 21196
rect 250500 21140 250528 21196
rect 250208 19628 250528 21140
rect 250208 19572 250236 19628
rect 250292 19572 250340 19628
rect 250396 19572 250444 19628
rect 250500 19572 250528 19628
rect 250208 18060 250528 19572
rect 250208 18004 250236 18060
rect 250292 18004 250340 18060
rect 250396 18004 250444 18060
rect 250500 18004 250528 18060
rect 250208 16492 250528 18004
rect 250208 16436 250236 16492
rect 250292 16436 250340 16492
rect 250396 16436 250444 16492
rect 250500 16436 250528 16492
rect 250208 14924 250528 16436
rect 250208 14868 250236 14924
rect 250292 14868 250340 14924
rect 250396 14868 250444 14924
rect 250500 14868 250528 14924
rect 250208 13356 250528 14868
rect 250208 13300 250236 13356
rect 250292 13300 250340 13356
rect 250396 13300 250444 13356
rect 250500 13300 250528 13356
rect 250208 11788 250528 13300
rect 250208 11732 250236 11788
rect 250292 11732 250340 11788
rect 250396 11732 250444 11788
rect 250500 11732 250528 11788
rect 250208 10220 250528 11732
rect 250208 10164 250236 10220
rect 250292 10164 250340 10220
rect 250396 10164 250444 10220
rect 250500 10164 250528 10220
rect 250208 8652 250528 10164
rect 250208 8596 250236 8652
rect 250292 8596 250340 8652
rect 250396 8596 250444 8652
rect 250500 8596 250528 8652
rect 250208 7084 250528 8596
rect 250208 7028 250236 7084
rect 250292 7028 250340 7084
rect 250396 7028 250444 7084
rect 250500 7028 250528 7084
rect 250208 5516 250528 7028
rect 250208 5460 250236 5516
rect 250292 5460 250340 5516
rect 250396 5460 250444 5516
rect 250500 5460 250528 5516
rect 250208 3948 250528 5460
rect 250208 3892 250236 3948
rect 250292 3892 250340 3948
rect 250396 3892 250444 3948
rect 250500 3892 250528 3948
rect 250208 3076 250528 3892
rect 265568 56476 265888 56508
rect 265568 56420 265596 56476
rect 265652 56420 265700 56476
rect 265756 56420 265804 56476
rect 265860 56420 265888 56476
rect 265568 54908 265888 56420
rect 265568 54852 265596 54908
rect 265652 54852 265700 54908
rect 265756 54852 265804 54908
rect 265860 54852 265888 54908
rect 265568 53340 265888 54852
rect 265568 53284 265596 53340
rect 265652 53284 265700 53340
rect 265756 53284 265804 53340
rect 265860 53284 265888 53340
rect 265568 51772 265888 53284
rect 265568 51716 265596 51772
rect 265652 51716 265700 51772
rect 265756 51716 265804 51772
rect 265860 51716 265888 51772
rect 265568 50204 265888 51716
rect 265568 50148 265596 50204
rect 265652 50148 265700 50204
rect 265756 50148 265804 50204
rect 265860 50148 265888 50204
rect 265568 48636 265888 50148
rect 265568 48580 265596 48636
rect 265652 48580 265700 48636
rect 265756 48580 265804 48636
rect 265860 48580 265888 48636
rect 265568 47068 265888 48580
rect 265568 47012 265596 47068
rect 265652 47012 265700 47068
rect 265756 47012 265804 47068
rect 265860 47012 265888 47068
rect 265568 45500 265888 47012
rect 265568 45444 265596 45500
rect 265652 45444 265700 45500
rect 265756 45444 265804 45500
rect 265860 45444 265888 45500
rect 265568 43932 265888 45444
rect 265568 43876 265596 43932
rect 265652 43876 265700 43932
rect 265756 43876 265804 43932
rect 265860 43876 265888 43932
rect 265568 42364 265888 43876
rect 265568 42308 265596 42364
rect 265652 42308 265700 42364
rect 265756 42308 265804 42364
rect 265860 42308 265888 42364
rect 265568 40796 265888 42308
rect 265568 40740 265596 40796
rect 265652 40740 265700 40796
rect 265756 40740 265804 40796
rect 265860 40740 265888 40796
rect 265568 39228 265888 40740
rect 265568 39172 265596 39228
rect 265652 39172 265700 39228
rect 265756 39172 265804 39228
rect 265860 39172 265888 39228
rect 265568 37660 265888 39172
rect 265568 37604 265596 37660
rect 265652 37604 265700 37660
rect 265756 37604 265804 37660
rect 265860 37604 265888 37660
rect 265568 36092 265888 37604
rect 265568 36036 265596 36092
rect 265652 36036 265700 36092
rect 265756 36036 265804 36092
rect 265860 36036 265888 36092
rect 265568 34524 265888 36036
rect 265568 34468 265596 34524
rect 265652 34468 265700 34524
rect 265756 34468 265804 34524
rect 265860 34468 265888 34524
rect 265568 32956 265888 34468
rect 265568 32900 265596 32956
rect 265652 32900 265700 32956
rect 265756 32900 265804 32956
rect 265860 32900 265888 32956
rect 265568 31388 265888 32900
rect 265568 31332 265596 31388
rect 265652 31332 265700 31388
rect 265756 31332 265804 31388
rect 265860 31332 265888 31388
rect 265568 29820 265888 31332
rect 265568 29764 265596 29820
rect 265652 29764 265700 29820
rect 265756 29764 265804 29820
rect 265860 29764 265888 29820
rect 265568 28252 265888 29764
rect 265568 28196 265596 28252
rect 265652 28196 265700 28252
rect 265756 28196 265804 28252
rect 265860 28196 265888 28252
rect 265568 26684 265888 28196
rect 265568 26628 265596 26684
rect 265652 26628 265700 26684
rect 265756 26628 265804 26684
rect 265860 26628 265888 26684
rect 265568 25116 265888 26628
rect 265568 25060 265596 25116
rect 265652 25060 265700 25116
rect 265756 25060 265804 25116
rect 265860 25060 265888 25116
rect 265568 23548 265888 25060
rect 265568 23492 265596 23548
rect 265652 23492 265700 23548
rect 265756 23492 265804 23548
rect 265860 23492 265888 23548
rect 265568 21980 265888 23492
rect 265568 21924 265596 21980
rect 265652 21924 265700 21980
rect 265756 21924 265804 21980
rect 265860 21924 265888 21980
rect 265568 20412 265888 21924
rect 265568 20356 265596 20412
rect 265652 20356 265700 20412
rect 265756 20356 265804 20412
rect 265860 20356 265888 20412
rect 265568 18844 265888 20356
rect 265568 18788 265596 18844
rect 265652 18788 265700 18844
rect 265756 18788 265804 18844
rect 265860 18788 265888 18844
rect 265568 17276 265888 18788
rect 265568 17220 265596 17276
rect 265652 17220 265700 17276
rect 265756 17220 265804 17276
rect 265860 17220 265888 17276
rect 265568 15708 265888 17220
rect 265568 15652 265596 15708
rect 265652 15652 265700 15708
rect 265756 15652 265804 15708
rect 265860 15652 265888 15708
rect 265568 14140 265888 15652
rect 265568 14084 265596 14140
rect 265652 14084 265700 14140
rect 265756 14084 265804 14140
rect 265860 14084 265888 14140
rect 265568 12572 265888 14084
rect 265568 12516 265596 12572
rect 265652 12516 265700 12572
rect 265756 12516 265804 12572
rect 265860 12516 265888 12572
rect 265568 11004 265888 12516
rect 265568 10948 265596 11004
rect 265652 10948 265700 11004
rect 265756 10948 265804 11004
rect 265860 10948 265888 11004
rect 265568 9436 265888 10948
rect 265568 9380 265596 9436
rect 265652 9380 265700 9436
rect 265756 9380 265804 9436
rect 265860 9380 265888 9436
rect 265568 7868 265888 9380
rect 265568 7812 265596 7868
rect 265652 7812 265700 7868
rect 265756 7812 265804 7868
rect 265860 7812 265888 7868
rect 265568 6300 265888 7812
rect 265568 6244 265596 6300
rect 265652 6244 265700 6300
rect 265756 6244 265804 6300
rect 265860 6244 265888 6300
rect 265568 4732 265888 6244
rect 265568 4676 265596 4732
rect 265652 4676 265700 4732
rect 265756 4676 265804 4732
rect 265860 4676 265888 4732
rect 265568 3164 265888 4676
rect 265568 3108 265596 3164
rect 265652 3108 265700 3164
rect 265756 3108 265804 3164
rect 265860 3108 265888 3164
rect 265568 3076 265888 3108
rect 280928 55692 281248 56508
rect 280928 55636 280956 55692
rect 281012 55636 281060 55692
rect 281116 55636 281164 55692
rect 281220 55636 281248 55692
rect 280928 54124 281248 55636
rect 280928 54068 280956 54124
rect 281012 54068 281060 54124
rect 281116 54068 281164 54124
rect 281220 54068 281248 54124
rect 280928 52556 281248 54068
rect 280928 52500 280956 52556
rect 281012 52500 281060 52556
rect 281116 52500 281164 52556
rect 281220 52500 281248 52556
rect 280928 50988 281248 52500
rect 280928 50932 280956 50988
rect 281012 50932 281060 50988
rect 281116 50932 281164 50988
rect 281220 50932 281248 50988
rect 280928 49420 281248 50932
rect 280928 49364 280956 49420
rect 281012 49364 281060 49420
rect 281116 49364 281164 49420
rect 281220 49364 281248 49420
rect 280928 47852 281248 49364
rect 280928 47796 280956 47852
rect 281012 47796 281060 47852
rect 281116 47796 281164 47852
rect 281220 47796 281248 47852
rect 280928 46284 281248 47796
rect 280928 46228 280956 46284
rect 281012 46228 281060 46284
rect 281116 46228 281164 46284
rect 281220 46228 281248 46284
rect 280928 44716 281248 46228
rect 280928 44660 280956 44716
rect 281012 44660 281060 44716
rect 281116 44660 281164 44716
rect 281220 44660 281248 44716
rect 280928 43148 281248 44660
rect 280928 43092 280956 43148
rect 281012 43092 281060 43148
rect 281116 43092 281164 43148
rect 281220 43092 281248 43148
rect 280928 41580 281248 43092
rect 280928 41524 280956 41580
rect 281012 41524 281060 41580
rect 281116 41524 281164 41580
rect 281220 41524 281248 41580
rect 280928 40012 281248 41524
rect 280928 39956 280956 40012
rect 281012 39956 281060 40012
rect 281116 39956 281164 40012
rect 281220 39956 281248 40012
rect 280928 38444 281248 39956
rect 280928 38388 280956 38444
rect 281012 38388 281060 38444
rect 281116 38388 281164 38444
rect 281220 38388 281248 38444
rect 280928 36876 281248 38388
rect 280928 36820 280956 36876
rect 281012 36820 281060 36876
rect 281116 36820 281164 36876
rect 281220 36820 281248 36876
rect 280928 35308 281248 36820
rect 280928 35252 280956 35308
rect 281012 35252 281060 35308
rect 281116 35252 281164 35308
rect 281220 35252 281248 35308
rect 280928 33740 281248 35252
rect 280928 33684 280956 33740
rect 281012 33684 281060 33740
rect 281116 33684 281164 33740
rect 281220 33684 281248 33740
rect 280928 32172 281248 33684
rect 280928 32116 280956 32172
rect 281012 32116 281060 32172
rect 281116 32116 281164 32172
rect 281220 32116 281248 32172
rect 280928 30604 281248 32116
rect 280928 30548 280956 30604
rect 281012 30548 281060 30604
rect 281116 30548 281164 30604
rect 281220 30548 281248 30604
rect 280928 29036 281248 30548
rect 280928 28980 280956 29036
rect 281012 28980 281060 29036
rect 281116 28980 281164 29036
rect 281220 28980 281248 29036
rect 280928 27468 281248 28980
rect 280928 27412 280956 27468
rect 281012 27412 281060 27468
rect 281116 27412 281164 27468
rect 281220 27412 281248 27468
rect 280928 25900 281248 27412
rect 280928 25844 280956 25900
rect 281012 25844 281060 25900
rect 281116 25844 281164 25900
rect 281220 25844 281248 25900
rect 280928 24332 281248 25844
rect 280928 24276 280956 24332
rect 281012 24276 281060 24332
rect 281116 24276 281164 24332
rect 281220 24276 281248 24332
rect 280928 22764 281248 24276
rect 280928 22708 280956 22764
rect 281012 22708 281060 22764
rect 281116 22708 281164 22764
rect 281220 22708 281248 22764
rect 280928 21196 281248 22708
rect 280928 21140 280956 21196
rect 281012 21140 281060 21196
rect 281116 21140 281164 21196
rect 281220 21140 281248 21196
rect 280928 19628 281248 21140
rect 280928 19572 280956 19628
rect 281012 19572 281060 19628
rect 281116 19572 281164 19628
rect 281220 19572 281248 19628
rect 280928 18060 281248 19572
rect 280928 18004 280956 18060
rect 281012 18004 281060 18060
rect 281116 18004 281164 18060
rect 281220 18004 281248 18060
rect 280928 16492 281248 18004
rect 280928 16436 280956 16492
rect 281012 16436 281060 16492
rect 281116 16436 281164 16492
rect 281220 16436 281248 16492
rect 280928 14924 281248 16436
rect 280928 14868 280956 14924
rect 281012 14868 281060 14924
rect 281116 14868 281164 14924
rect 281220 14868 281248 14924
rect 280928 13356 281248 14868
rect 280928 13300 280956 13356
rect 281012 13300 281060 13356
rect 281116 13300 281164 13356
rect 281220 13300 281248 13356
rect 280928 11788 281248 13300
rect 280928 11732 280956 11788
rect 281012 11732 281060 11788
rect 281116 11732 281164 11788
rect 281220 11732 281248 11788
rect 280928 10220 281248 11732
rect 280928 10164 280956 10220
rect 281012 10164 281060 10220
rect 281116 10164 281164 10220
rect 281220 10164 281248 10220
rect 280928 8652 281248 10164
rect 280928 8596 280956 8652
rect 281012 8596 281060 8652
rect 281116 8596 281164 8652
rect 281220 8596 281248 8652
rect 280928 7084 281248 8596
rect 280928 7028 280956 7084
rect 281012 7028 281060 7084
rect 281116 7028 281164 7084
rect 281220 7028 281248 7084
rect 280928 5516 281248 7028
rect 280928 5460 280956 5516
rect 281012 5460 281060 5516
rect 281116 5460 281164 5516
rect 281220 5460 281248 5516
rect 280928 3948 281248 5460
rect 280928 3892 280956 3948
rect 281012 3892 281060 3948
rect 281116 3892 281164 3948
rect 281220 3892 281248 3948
rect 280928 3076 281248 3892
rect 296288 56476 296608 56508
rect 296288 56420 296316 56476
rect 296372 56420 296420 56476
rect 296476 56420 296524 56476
rect 296580 56420 296608 56476
rect 296288 54908 296608 56420
rect 296288 54852 296316 54908
rect 296372 54852 296420 54908
rect 296476 54852 296524 54908
rect 296580 54852 296608 54908
rect 296288 53340 296608 54852
rect 296288 53284 296316 53340
rect 296372 53284 296420 53340
rect 296476 53284 296524 53340
rect 296580 53284 296608 53340
rect 296288 51772 296608 53284
rect 296288 51716 296316 51772
rect 296372 51716 296420 51772
rect 296476 51716 296524 51772
rect 296580 51716 296608 51772
rect 296288 50204 296608 51716
rect 296288 50148 296316 50204
rect 296372 50148 296420 50204
rect 296476 50148 296524 50204
rect 296580 50148 296608 50204
rect 296288 48636 296608 50148
rect 296288 48580 296316 48636
rect 296372 48580 296420 48636
rect 296476 48580 296524 48636
rect 296580 48580 296608 48636
rect 296288 47068 296608 48580
rect 296288 47012 296316 47068
rect 296372 47012 296420 47068
rect 296476 47012 296524 47068
rect 296580 47012 296608 47068
rect 296288 45500 296608 47012
rect 296288 45444 296316 45500
rect 296372 45444 296420 45500
rect 296476 45444 296524 45500
rect 296580 45444 296608 45500
rect 296288 43932 296608 45444
rect 296288 43876 296316 43932
rect 296372 43876 296420 43932
rect 296476 43876 296524 43932
rect 296580 43876 296608 43932
rect 296288 42364 296608 43876
rect 296288 42308 296316 42364
rect 296372 42308 296420 42364
rect 296476 42308 296524 42364
rect 296580 42308 296608 42364
rect 296288 40796 296608 42308
rect 296288 40740 296316 40796
rect 296372 40740 296420 40796
rect 296476 40740 296524 40796
rect 296580 40740 296608 40796
rect 296288 39228 296608 40740
rect 296288 39172 296316 39228
rect 296372 39172 296420 39228
rect 296476 39172 296524 39228
rect 296580 39172 296608 39228
rect 296288 37660 296608 39172
rect 296288 37604 296316 37660
rect 296372 37604 296420 37660
rect 296476 37604 296524 37660
rect 296580 37604 296608 37660
rect 296288 36092 296608 37604
rect 296288 36036 296316 36092
rect 296372 36036 296420 36092
rect 296476 36036 296524 36092
rect 296580 36036 296608 36092
rect 296288 34524 296608 36036
rect 296288 34468 296316 34524
rect 296372 34468 296420 34524
rect 296476 34468 296524 34524
rect 296580 34468 296608 34524
rect 296288 32956 296608 34468
rect 296288 32900 296316 32956
rect 296372 32900 296420 32956
rect 296476 32900 296524 32956
rect 296580 32900 296608 32956
rect 296288 31388 296608 32900
rect 296288 31332 296316 31388
rect 296372 31332 296420 31388
rect 296476 31332 296524 31388
rect 296580 31332 296608 31388
rect 296288 29820 296608 31332
rect 296288 29764 296316 29820
rect 296372 29764 296420 29820
rect 296476 29764 296524 29820
rect 296580 29764 296608 29820
rect 296288 28252 296608 29764
rect 296288 28196 296316 28252
rect 296372 28196 296420 28252
rect 296476 28196 296524 28252
rect 296580 28196 296608 28252
rect 296288 26684 296608 28196
rect 296288 26628 296316 26684
rect 296372 26628 296420 26684
rect 296476 26628 296524 26684
rect 296580 26628 296608 26684
rect 296288 25116 296608 26628
rect 296288 25060 296316 25116
rect 296372 25060 296420 25116
rect 296476 25060 296524 25116
rect 296580 25060 296608 25116
rect 296288 23548 296608 25060
rect 296288 23492 296316 23548
rect 296372 23492 296420 23548
rect 296476 23492 296524 23548
rect 296580 23492 296608 23548
rect 296288 21980 296608 23492
rect 296288 21924 296316 21980
rect 296372 21924 296420 21980
rect 296476 21924 296524 21980
rect 296580 21924 296608 21980
rect 296288 20412 296608 21924
rect 296288 20356 296316 20412
rect 296372 20356 296420 20412
rect 296476 20356 296524 20412
rect 296580 20356 296608 20412
rect 296288 18844 296608 20356
rect 296288 18788 296316 18844
rect 296372 18788 296420 18844
rect 296476 18788 296524 18844
rect 296580 18788 296608 18844
rect 296288 17276 296608 18788
rect 296288 17220 296316 17276
rect 296372 17220 296420 17276
rect 296476 17220 296524 17276
rect 296580 17220 296608 17276
rect 296288 15708 296608 17220
rect 296288 15652 296316 15708
rect 296372 15652 296420 15708
rect 296476 15652 296524 15708
rect 296580 15652 296608 15708
rect 296288 14140 296608 15652
rect 296288 14084 296316 14140
rect 296372 14084 296420 14140
rect 296476 14084 296524 14140
rect 296580 14084 296608 14140
rect 296288 12572 296608 14084
rect 296288 12516 296316 12572
rect 296372 12516 296420 12572
rect 296476 12516 296524 12572
rect 296580 12516 296608 12572
rect 296288 11004 296608 12516
rect 296288 10948 296316 11004
rect 296372 10948 296420 11004
rect 296476 10948 296524 11004
rect 296580 10948 296608 11004
rect 296288 9436 296608 10948
rect 296288 9380 296316 9436
rect 296372 9380 296420 9436
rect 296476 9380 296524 9436
rect 296580 9380 296608 9436
rect 296288 7868 296608 9380
rect 296288 7812 296316 7868
rect 296372 7812 296420 7868
rect 296476 7812 296524 7868
rect 296580 7812 296608 7868
rect 296288 6300 296608 7812
rect 296288 6244 296316 6300
rect 296372 6244 296420 6300
rect 296476 6244 296524 6300
rect 296580 6244 296608 6300
rect 296288 4732 296608 6244
rect 296288 4676 296316 4732
rect 296372 4676 296420 4732
rect 296476 4676 296524 4732
rect 296580 4676 296608 4732
rect 296288 3164 296608 4676
rect 296288 3108 296316 3164
rect 296372 3108 296420 3164
rect 296476 3108 296524 3164
rect 296580 3108 296608 3164
rect 296288 3076 296608 3108
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _106_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 218624 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _107_
timestamp 1698175906
transform 1 0 217280 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _108_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 222096 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _109_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 219632 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _110_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 195776 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _111_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 193424 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _112_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 201264 0 1 4704
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _113_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 201600 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _114_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 220080 0 1 3136
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _115_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 223440 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _116_
timestamp 1698175906
transform -1 0 221648 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _117_
timestamp 1698175906
transform -1 0 222320 0 -1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _118_
timestamp 1698175906
transform -1 0 195552 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _119_
timestamp 1698175906
transform 1 0 191520 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _120_
timestamp 1698175906
transform -1 0 202832 0 -1 6272
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _121_
timestamp 1698175906
transform 1 0 202832 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _122_
timestamp 1698175906
transform 1 0 220864 0 1 3136
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _123_
timestamp 1698175906
transform -1 0 224336 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _124_
timestamp 1698175906
transform -1 0 220864 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _125_
timestamp 1698175906
transform -1 0 222096 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _126_
timestamp 1698175906
transform -1 0 195776 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1698175906
transform 1 0 192528 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _128_
timestamp 1698175906
transform 1 0 196000 0 1 6272
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _129_
timestamp 1698175906
transform -1 0 204400 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _130_
timestamp 1698175906
transform -1 0 217728 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _131_
timestamp 1698175906
transform -1 0 219296 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _132_
timestamp 1698175906
transform -1 0 218624 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _133_
timestamp 1698175906
transform 1 0 217168 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _134_
timestamp 1698175906
transform -1 0 195776 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _135_
timestamp 1698175906
transform 1 0 184240 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _136_
timestamp 1698175906
transform 1 0 201488 0 1 6272
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _137_
timestamp 1698175906
transform -1 0 206416 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _138_
timestamp 1698175906
transform 1 0 216048 0 -1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _139_
timestamp 1698175906
transform -1 0 218064 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _140_
timestamp 1698175906
transform -1 0 217392 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _141_
timestamp 1698175906
transform -1 0 216944 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _142_
timestamp 1698175906
transform -1 0 188496 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _143_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 185808 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 186704 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _145_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 191072 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _146_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 188832 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _147_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 200256 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _148_
timestamp 1698175906
transform 1 0 205632 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _149_
timestamp 1698175906
transform 1 0 201152 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _150_
timestamp 1698175906
transform 1 0 204400 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 198688 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _152_
timestamp 1698175906
transform -1 0 207536 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _153_
timestamp 1698175906
transform 1 0 205744 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _154_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 187712 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _155_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 186144 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _156_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 206080 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _157_
timestamp 1698175906
transform 1 0 204288 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _158_
timestamp 1698175906
transform 1 0 206416 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _159_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 199808 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform 1 0 200592 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _161_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 209104 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _162_
timestamp 1698175906
transform 1 0 188944 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _163_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 208992 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _164_
timestamp 1698175906
transform 1 0 201264 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _165_
timestamp 1698175906
transform -1 0 190848 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _166_
timestamp 1698175906
transform 1 0 186592 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _167_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 199360 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _168_
timestamp 1698175906
transform -1 0 210560 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _169_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 211904 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _170_
timestamp 1698175906
transform 1 0 209664 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _171_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 204512 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _172_
timestamp 1698175906
transform -1 0 214816 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _173_
timestamp 1698175906
transform -1 0 212576 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _174_
timestamp 1698175906
transform -1 0 203392 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _175_
timestamp 1698175906
transform 1 0 201488 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _176_
timestamp 1698175906
transform -1 0 189504 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _177_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 186816 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _178_
timestamp 1698175906
transform -1 0 214144 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _179_
timestamp 1698175906
transform -1 0 212800 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _180_
timestamp 1698175906
transform 1 0 209440 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _181_
timestamp 1698175906
transform -1 0 200592 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _182_
timestamp 1698175906
transform -1 0 191296 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _183_
timestamp 1698175906
transform 1 0 188496 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _184_
timestamp 1698175906
transform 1 0 182112 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _185_
timestamp 1698175906
transform -1 0 194992 0 -1 4704
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _186_
timestamp 1698175906
transform 1 0 200592 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _187_
timestamp 1698175906
transform -1 0 214144 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _188_
timestamp 1698175906
transform -1 0 207648 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _189_
timestamp 1698175906
transform -1 0 209664 0 1 3136
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _190_
timestamp 1698175906
transform 1 0 214480 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _191_
timestamp 1698175906
transform -1 0 216496 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _192_
timestamp 1698175906
transform -1 0 211568 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _193_
timestamp 1698175906
transform 1 0 209328 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _194_
timestamp 1698175906
transform -1 0 186592 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _195_
timestamp 1698175906
transform 1 0 182560 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _196_
timestamp 1698175906
transform -1 0 192528 0 1 4704
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _197_
timestamp 1698175906
transform 1 0 205632 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _198_
timestamp 1698175906
transform -1 0 211792 0 1 3136
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _199_
timestamp 1698175906
transform -1 0 215600 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _200_
timestamp 1698175906
transform -1 0 211904 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _201_
timestamp 1698175906
transform -1 0 211792 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _202_
timestamp 1698175906
transform -1 0 186592 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _203_
timestamp 1698175906
transform 1 0 182112 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _204_
timestamp 1698175906
transform -1 0 192528 0 1 6272
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _205_
timestamp 1698175906
transform -1 0 205296 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _206_
timestamp 1698175906
transform 1 0 204736 0 1 3136
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _207_
timestamp 1698175906
transform 1 0 210560 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _208_
timestamp 1698175906
transform 1 0 211904 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _209_
timestamp 1698175906
transform 1 0 214032 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _210_
timestamp 1698175906
transform -1 0 215712 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _211_
timestamp 1698175906
transform 1 0 207648 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _212_
timestamp 1698175906
transform -1 0 212576 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _213_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 213024 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _214_
timestamp 1698175906
transform -1 0 185584 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _215_
timestamp 1698175906
transform 1 0 190624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _216_
timestamp 1698175906
transform -1 0 194768 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _217_
timestamp 1698175906
transform -1 0 198688 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _218_
timestamp 1698175906
transform 1 0 196224 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _219_
timestamp 1698175906
transform 1 0 195888 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _220_
timestamp 1698175906
transform -1 0 202832 0 -1 4704
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _221_
timestamp 1698175906
transform -1 0 203728 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _222_
timestamp 1698175906
transform -1 0 204288 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _223_
timestamp 1698175906
transform 1 0 201376 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _224_
timestamp 1698175906
transform 1 0 216272 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _225_
timestamp 1698175906
transform 1 0 219520 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _226_
timestamp 1698175906
transform 1 0 218064 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _227_
timestamp 1698175906
transform -1 0 223440 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 186256 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 190176 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 182336 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform -1 0 132720 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 134848 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 140336 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform -1 0 148400 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform -1 0 154112 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 156464 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 162288 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform -1 0 169904 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform -1 0 175280 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 179312 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 183120 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform -1 0 191408 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform -1 0 194880 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  _252_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 130480 0 1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _253_
timestamp 1698175906
transform -1 0 135968 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _254_
timestamp 1698175906
transform -1 0 141232 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _255_
timestamp 1698175906
transform -1 0 146160 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _256_
timestamp 1698175906
transform -1 0 151760 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _257_
timestamp 1698175906
transform -1 0 157360 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _258_
timestamp 1698175906
transform -1 0 162512 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _259_
timestamp 1698175906
transform -1 0 168112 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _260_
timestamp 1698175906
transform -1 0 172928 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _261_
timestamp 1698175906
transform -1 0 12096 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _262_
timestamp 1698175906
transform 1 0 71232 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _263_
timestamp 1698175906
transform 1 0 74928 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _264_
timestamp 1698175906
transform 1 0 78512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _265_
timestamp 1698175906
transform 1 0 82992 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _266_
timestamp 1698175906
transform 1 0 86576 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _267_
timestamp 1698175906
transform 1 0 89152 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _268_
timestamp 1698175906
transform 1 0 93744 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _269_
timestamp 1698175906
transform 1 0 96320 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__A4 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 222320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__A1
timestamp 1698175906
transform -1 0 219632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__B2
timestamp 1698175906
transform 1 0 196000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__I
timestamp 1698175906
transform 1 0 193872 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__B2
timestamp 1698175906
transform -1 0 201376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__C1
timestamp 1698175906
transform 1 0 203952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__A4
timestamp 1698175906
transform -1 0 200928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__A2
timestamp 1698175906
transform -1 0 223664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__A4
timestamp 1698175906
transform -1 0 222096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__A1
timestamp 1698175906
transform -1 0 222096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__B2
timestamp 1698175906
transform 1 0 197568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I
timestamp 1698175906
transform -1 0 191744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__B2
timestamp 1698175906
transform 1 0 204848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__C1
timestamp 1698175906
transform 1 0 203616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__A4
timestamp 1698175906
transform 1 0 206640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__A2
timestamp 1698175906
transform -1 0 224784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__A4
timestamp 1698175906
transform 1 0 220864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__A1
timestamp 1698175906
transform 1 0 220640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__B2
timestamp 1698175906
transform -1 0 196000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1698175906
transform 1 0 194992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__B2
timestamp 1698175906
transform -1 0 199248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__C1
timestamp 1698175906
transform 1 0 202272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__A4
timestamp 1698175906
transform 1 0 204512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__A2
timestamp 1698175906
transform 1 0 219296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__A4
timestamp 1698175906
transform 1 0 219520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__B2
timestamp 1698175906
transform 1 0 196000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__I
timestamp 1698175906
transform 1 0 184016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__B1
timestamp 1698175906
transform 1 0 206976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__B2
timestamp 1698175906
transform 1 0 207424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__C1
timestamp 1698175906
transform 1 0 207872 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__137__A4
timestamp 1698175906
transform 1 0 207536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__A2
timestamp 1698175906
transform 1 0 217056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__A3
timestamp 1698175906
transform 1 0 215824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__A2
timestamp 1698175906
transform -1 0 219184 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__A4
timestamp 1698175906
transform 1 0 217392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__A2
timestamp 1698175906
transform -1 0 189504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__B1
timestamp 1698175906
transform -1 0 190512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__B2
timestamp 1698175906
transform 1 0 191072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__A1
timestamp 1698175906
transform 1 0 187488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__A1
timestamp 1698175906
transform -1 0 187936 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__146__I
timestamp 1698175906
transform 1 0 188832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__I
timestamp 1698175906
transform 1 0 200032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__I
timestamp 1698175906
transform 1 0 200928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__I
timestamp 1698175906
transform 1 0 198464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I
timestamp 1698175906
transform 1 0 187936 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__I
timestamp 1698175906
transform 1 0 199584 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__I
timestamp 1698175906
transform 1 0 190736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__A4
timestamp 1698175906
transform -1 0 208768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__A1
timestamp 1698175906
transform -1 0 199136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__A2
timestamp 1698175906
transform 1 0 199136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__I
timestamp 1698175906
transform 1 0 209440 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A2
timestamp 1698175906
transform 1 0 208880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__A2
timestamp 1698175906
transform 1 0 209440 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__I
timestamp 1698175906
transform 1 0 189280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__A4
timestamp 1698175906
transform 1 0 209216 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__A2
timestamp 1698175906
transform -1 0 199696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__I
timestamp 1698175906
transform -1 0 181664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__B2
timestamp 1698175906
transform -1 0 195888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__C1
timestamp 1698175906
transform -1 0 196896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__A4
timestamp 1698175906
transform 1 0 207984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__A2
timestamp 1698175906
transform -1 0 216944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__A4
timestamp 1698175906
transform 1 0 212800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__B2
timestamp 1698175906
transform -1 0 186816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__I
timestamp 1698175906
transform 1 0 182784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__B2
timestamp 1698175906
transform 1 0 195440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__C1
timestamp 1698175906
transform 1 0 194320 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__A4
timestamp 1698175906
transform 1 0 206304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__A2
timestamp 1698175906
transform 1 0 215936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__A4
timestamp 1698175906
transform 1 0 211904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__B2
timestamp 1698175906
transform -1 0 186816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1698175906
transform -1 0 182112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__B2
timestamp 1698175906
transform 1 0 192752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__C1
timestamp 1698175906
transform 1 0 193200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__A4
timestamp 1698175906
transform 1 0 210560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__A2
timestamp 1698175906
transform -1 0 215936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__A4
timestamp 1698175906
transform -1 0 213472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__B2
timestamp 1698175906
transform 1 0 187040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__I
timestamp 1698175906
transform -1 0 190624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__I
timestamp 1698175906
transform -1 0 195440 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__I
timestamp 1698175906
transform -1 0 198240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__B2
timestamp 1698175906
transform -1 0 208096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__C1
timestamp 1698175906
transform -1 0 208320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__A4
timestamp 1698175906
transform -1 0 200480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__I
timestamp 1698175906
transform 1 0 217952 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__A2
timestamp 1698175906
transform 1 0 223664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 185808 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__D
timestamp 1698175906
transform -1 0 186256 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 189728 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__D
timestamp 1698175906
transform -1 0 189504 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 182112 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__D
timestamp 1698175906
transform 1 0 181440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 132944 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 138320 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 143808 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 148624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 150080 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 156240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 161840 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 170352 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 175504 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 182784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 182896 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 187936 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 191408 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__I
timestamp 1698175906
transform -1 0 12544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__I
timestamp 1698175906
transform -1 0 71232 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__I
timestamp 1698175906
transform -1 0 74928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__I
timestamp 1698175906
transform 1 0 78288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__I
timestamp 1698175906
transform -1 0 82992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__I
timestamp 1698175906
transform -1 0 86576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__I
timestamp 1698175906
transform 1 0 88704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__I
timestamp 1698175906
transform 1 0 93520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__I
timestamp 1698175906
transform -1 0 96320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698175906
transform -1 0 162064 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_0__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 153216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_1__f_wb_clk_i_I
timestamp 1698175906
transform -1 0 177744 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698175906
transform -1 0 123200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698175906
transform -1 0 127008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698175906
transform -1 0 130816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698175906
transform -1 0 133840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698175906
transform -1 0 137424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698175906
transform -1 0 141008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698175906
transform -1 0 144592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698175906
transform -1 0 148176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698175906
transform -1 0 151760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698175906
transform -1 0 155344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698175906
transform -1 0 158928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698175906
transform -1 0 162512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698175906
transform -1 0 166096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698175906
transform -1 0 169680 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698175906
transform -1 0 172704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698175906
transform -1 0 176512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698175906
transform -1 0 180320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698175906
transform -1 0 183456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698175906
transform -1 0 187936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698175906
transform -1 0 190176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698175906
transform 1 0 197120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698175906
transform 1 0 199808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698175906
transform -1 0 205744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698175906
transform 1 0 208432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698175906
transform 1 0 212016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698175906
transform -1 0 212688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698175906
transform -1 0 215488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698175906
transform -1 0 219408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698175906
transform -1 0 223440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698175906
transform -1 0 227024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698175906
transform -1 0 230608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698175906
transform -1 0 233632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698175906
transform -1 0 237440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698175906
transform -1 0 241248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698175906
transform -1 0 245056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698175906
transform -1 0 248864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698175906
transform -1 0 252672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698175906
transform -1 0 255696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698175906
transform -1 0 259280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698175906
transform -1 0 262864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698175906
transform -1 0 266448 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698175906
transform -1 0 270032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698175906
transform -1 0 273616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698175906
transform -1 0 277200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698175906
transform -1 0 280784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698175906
transform -1 0 284368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698175906
transform -1 0 287952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698175906
transform -1 0 291536 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698175906
transform -1 0 211792 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698175906
transform -1 0 217168 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698175906
transform -1 0 222208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698175906
transform -1 0 227920 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698175906
transform -1 0 233632 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698175906
transform -1 0 238672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698175906
transform -1 0 244048 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698175906
transform -1 0 248864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698175906
transform -1 0 254800 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698175906
transform 1 0 260064 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698175906
transform -1 0 265552 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698175906
transform 1 0 271488 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698175906
transform -1 0 276304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698175906
transform 1 0 283584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1698175906
transform -1 0 286944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1698175906
transform -1 0 292432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1698175906
transform -1 0 18256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1698175906
transform -1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1698175906
transform -1 0 29008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1698175906
transform -1 0 34384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1698175906
transform -1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1698175906
transform -1 0 45136 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1698175906
transform -1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1698175906
transform -1 0 55888 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1698175906
transform -1 0 61264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1698175906
transform -1 0 109648 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1698175906
transform -1 0 115584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1698175906
transform -1 0 168896 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1698175906
transform -1 0 174160 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1698175906
transform -1 0 179536 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1698175906
transform -1 0 184912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1698175906
transform 1 0 192192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1698175906
transform -1 0 195552 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1698175906
transform -1 0 120400 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1698175906
transform -1 0 125776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1698175906
transform -1 0 130816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1698175906
transform -1 0 136528 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1698175906
transform -1 0 142240 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1698175906
transform -1 0 147280 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1698175906
transform -1 0 152656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1698175906
transform -1 0 157472 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1698175906
transform -1 0 163408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1698175906
transform -1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output92_I
timestamp 1698175906
transform -1 0 43904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output93_I
timestamp 1698175906
transform -1 0 47712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output94_I
timestamp 1698175906
transform 1 0 50736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output95_I
timestamp 1698175906
transform 1 0 54320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output96_I
timestamp 1698175906
transform -1 0 58352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output97_I
timestamp 1698175906
transform -1 0 62048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output98_I
timestamp 1698175906
transform -1 0 65856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output99_I
timestamp 1698175906
transform -1 0 69664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output100_I
timestamp 1698175906
transform -1 0 73472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output110_I
timestamp 1698175906
transform -1 0 104832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output111_I
timestamp 1698175906
transform -1 0 108640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output112_I
timestamp 1698175906
transform -1 0 111888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output113_I
timestamp 1698175906
transform -1 0 115472 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output114_I
timestamp 1698175906
transform -1 0 119280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output115_I
timestamp 1698175906
transform 1 0 122528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output116_I
timestamp 1698175906
transform -1 0 203840 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output117_I
timestamp 1698175906
transform -1 0 206976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output118_I
timestamp 1698175906
transform -1 0 70560 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output119_I
timestamp 1698175906
transform 1 0 75152 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output120_I
timestamp 1698175906
transform -1 0 81088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output121_I
timestamp 1698175906
transform -1 0 85792 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output122_I
timestamp 1698175906
transform -1 0 92512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output123_I
timestamp 1698175906
transform -1 0 97216 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output124_I
timestamp 1698175906
transform 1 0 102704 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output125_I
timestamp 1698175906
transform -1 0 107744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 162288 0 1 53312
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1698175906
transform -1 0 152992 0 1 54880
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1698175906
transform 1 0 177968 0 1 53312
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_100 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_104 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_120 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_124
timestamp 1698175906
transform 1 0 15232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_126 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_131
timestamp 1698175906
transform 1 0 16016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698175906
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_154
timestamp 1698175906
transform 1 0 18592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_158
timestamp 1698175906
transform 1 0 19040 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_163
timestamp 1698175906
transform 1 0 19600 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_167
timestamp 1698175906
transform 1 0 20048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_188
timestamp 1698175906
transform 1 0 22400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_190
timestamp 1698175906
transform 1 0 22624 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_195 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23184 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_222
timestamp 1698175906
transform 1 0 26208 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_227
timestamp 1698175906
transform 1 0 26768 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_235
timestamp 1698175906
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_248
timestamp 1698175906
transform 1 0 29120 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_252
timestamp 1698175906
transform 1 0 29568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_254
timestamp 1698175906
transform 1 0 29792 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_259
timestamp 1698175906
transform 1 0 30352 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_267
timestamp 1698175906
transform 1 0 31248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698175906
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_282
timestamp 1698175906
transform 1 0 32928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_286
timestamp 1698175906
transform 1 0 33376 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_291
timestamp 1698175906
transform 1 0 33936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_299
timestamp 1698175906
transform 1 0 34832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303
timestamp 1698175906
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698175906
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_316
timestamp 1698175906
transform 1 0 36736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_318
timestamp 1698175906
transform 1 0 36960 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_323
timestamp 1698175906
transform 1 0 37520 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698175906
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698175906
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_380
timestamp 1698175906
transform 1 0 43904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_410
timestamp 1698175906
transform 1 0 47264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_414
timestamp 1698175906
transform 1 0 47712 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_441
timestamp 1698175906
transform 1 0 50736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_444
timestamp 1698175906
transform 1 0 51072 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_446
timestamp 1698175906
transform 1 0 51296 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_473
timestamp 1698175906
transform 1 0 54320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_475
timestamp 1698175906
transform 1 0 54544 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_478
timestamp 1698175906
transform 1 0 54880 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_505
timestamp 1698175906
transform 1 0 57904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_509
timestamp 1698175906
transform 1 0 58352 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_538
timestamp 1698175906
transform 1 0 61600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_542
timestamp 1698175906
transform 1 0 62048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_572
timestamp 1698175906
transform 1 0 65408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_576
timestamp 1698175906
transform 1 0 65856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_606
timestamp 1698175906
transform 1 0 69216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_610
timestamp 1698175906
transform 1 0 69664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_640
timestamp 1698175906
transform 1 0 73024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_644
timestamp 1698175906
transform 1 0 73472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_674
timestamp 1698175906
transform 1 0 76832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_678
timestamp 1698175906
transform 1 0 77280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_682
timestamp 1698175906
transform 1 0 77728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_686
timestamp 1698175906
transform 1 0 78176 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_695
timestamp 1698175906
transform 1 0 79184 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_711
timestamp 1698175906
transform 1 0 80976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_713
timestamp 1698175906
transform 1 0 81200 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_716
timestamp 1698175906
transform 1 0 81536 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_724
timestamp 1698175906
transform 1 0 82432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_726
timestamp 1698175906
transform 1 0 82656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_729
timestamp 1698175906
transform 1 0 82992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_745
timestamp 1698175906
transform 1 0 84784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_747
timestamp 1698175906
transform 1 0 85008 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_750
timestamp 1698175906
transform 1 0 85344 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_758
timestamp 1698175906
transform 1 0 86240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_761
timestamp 1698175906
transform 1 0 86576 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_777
timestamp 1698175906
transform 1 0 88368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_779
timestamp 1698175906
transform 1 0 88592 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_790
timestamp 1698175906
transform 1 0 89824 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_806
timestamp 1698175906
transform 1 0 91616 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_814
timestamp 1698175906
transform 1 0 92512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_818
timestamp 1698175906
transform 1 0 92960 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_822
timestamp 1698175906
transform 1 0 93408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_852
timestamp 1698175906
transform 1 0 96768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_856
timestamp 1698175906
transform 1 0 97216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_886
timestamp 1698175906
transform 1 0 100576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_890
timestamp 1698175906
transform 1 0 101024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_920
timestamp 1698175906
transform 1 0 104384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_924
timestamp 1698175906
transform 1 0 104832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_954
timestamp 1698175906
transform 1 0 108192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_958
timestamp 1698175906
transform 1 0 108640 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_985
timestamp 1698175906
transform 1 0 111664 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_988
timestamp 1698175906
transform 1 0 112000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_990
timestamp 1698175906
transform 1 0 112224 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1017
timestamp 1698175906
transform 1 0 115248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1019
timestamp 1698175906
transform 1 0 115472 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1022
timestamp 1698175906
transform 1 0 115808 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1049
timestamp 1698175906
transform 1 0 118832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1053
timestamp 1698175906
transform 1 0 119280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1082
timestamp 1698175906
transform 1 0 122528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1096
timestamp 1698175906
transform 1 0 124096 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1112
timestamp 1698175906
transform 1 0 125888 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1130
timestamp 1698175906
transform 1 0 127904 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1146
timestamp 1698175906
transform 1 0 129696 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1164
timestamp 1698175906
transform 1 0 131712 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1180
timestamp 1698175906
transform 1 0 133504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1189
timestamp 1698175906
transform 1 0 134512 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1192
timestamp 1698175906
transform 1 0 134848 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1208
timestamp 1698175906
transform 1 0 136640 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1212
timestamp 1698175906
transform 1 0 137088 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1221
timestamp 1698175906
transform 1 0 138096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1223
timestamp 1698175906
transform 1 0 138320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1226
timestamp 1698175906
transform 1 0 138656 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1242
timestamp 1698175906
transform 1 0 140448 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1244
timestamp 1698175906
transform 1 0 140672 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1253
timestamp 1698175906
transform 1 0 141680 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1257
timestamp 1698175906
transform 1 0 142128 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1260
timestamp 1698175906
transform 1 0 142464 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1276
timestamp 1698175906
transform 1 0 144256 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1285
timestamp 1698175906
transform 1 0 145264 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1289
timestamp 1698175906
transform 1 0 145712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1291
timestamp 1698175906
transform 1 0 145936 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1294
timestamp 1698175906
transform 1 0 146272 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1302
timestamp 1698175906
transform 1 0 147168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1306
timestamp 1698175906
transform 1 0 147616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1308
timestamp 1698175906
transform 1 0 147840 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1317
timestamp 1698175906
transform 1 0 148848 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1325
timestamp 1698175906
transform 1 0 149744 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1328
timestamp 1698175906
transform 1 0 150080 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1336
timestamp 1698175906
transform 1 0 150976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1340
timestamp 1698175906
transform 1 0 151424 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1349
timestamp 1698175906
transform 1 0 152432 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1357
timestamp 1698175906
transform 1 0 153328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1359
timestamp 1698175906
transform 1 0 153552 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1362
timestamp 1698175906
transform 1 0 153888 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1370
timestamp 1698175906
transform 1 0 154784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1372
timestamp 1698175906
transform 1 0 155008 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1381
timestamp 1698175906
transform 1 0 156016 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1389
timestamp 1698175906
transform 1 0 156912 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1393
timestamp 1698175906
transform 1 0 157360 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1396
timestamp 1698175906
transform 1 0 157696 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1404
timestamp 1698175906
transform 1 0 158592 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1413
timestamp 1698175906
transform 1 0 159600 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1421
timestamp 1698175906
transform 1 0 160496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1425
timestamp 1698175906
transform 1 0 160944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1427
timestamp 1698175906
transform 1 0 161168 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1430
timestamp 1698175906
transform 1 0 161504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1434
timestamp 1698175906
transform 1 0 161952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1436
timestamp 1698175906
transform 1 0 162176 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1445
timestamp 1698175906
transform 1 0 163184 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1461
timestamp 1698175906
transform 1 0 164976 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1464
timestamp 1698175906
transform 1 0 165312 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1468
timestamp 1698175906
transform 1 0 165760 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1477
timestamp 1698175906
transform 1 0 166768 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1493
timestamp 1698175906
transform 1 0 168560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1495
timestamp 1698175906
transform 1 0 168784 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1498
timestamp 1698175906
transform 1 0 169120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1500
timestamp 1698175906
transform 1 0 169344 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1509
timestamp 1698175906
transform 1 0 170352 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1525
timestamp 1698175906
transform 1 0 172144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1527
timestamp 1698175906
transform 1 0 172368 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1532
timestamp 1698175906
transform 1 0 172928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1534
timestamp 1698175906
transform 1 0 173152 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1541
timestamp 1698175906
transform 1 0 173936 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1557
timestamp 1698175906
transform 1 0 175728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1561
timestamp 1698175906
transform 1 0 176176 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1566
timestamp 1698175906
transform 1 0 176736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1573
timestamp 1698175906
transform 1 0 177520 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1589
timestamp 1698175906
transform 1 0 179312 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1593
timestamp 1698175906
transform 1 0 179760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1595
timestamp 1698175906
transform 1 0 179984 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1606
timestamp 1698175906
transform 1 0 181216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1610
timestamp 1698175906
transform 1 0 181664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1618
timestamp 1698175906
transform 1 0 182560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1622
timestamp 1698175906
transform 1 0 183008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1650
timestamp 1698175906
transform 1 0 186144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1656
timestamp 1698175906
transform 1 0 186816 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1674
timestamp 1698175906
transform 1 0 188832 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1682
timestamp 1698175906
transform 1 0 189728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1686
timestamp 1698175906
transform 1 0 190176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1742
timestamp 1698175906
transform 1 0 196448 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1746
timestamp 1698175906
transform 1 0 196896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1750
timestamp 1698175906
transform 1 0 197344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1754
timestamp 1698175906
transform 1 0 197792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1758
timestamp 1698175906
transform 1 0 198240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1765
timestamp 1698175906
transform 1 0 199024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1767
timestamp 1698175906
transform 1 0 199248 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1770
timestamp 1698175906
transform 1 0 199584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1774
timestamp 1698175906
transform 1 0 200032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1778
timestamp 1698175906
transform 1 0 200480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1782
timestamp 1698175906
transform 1 0 200928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1812
timestamp 1698175906
transform 1 0 204288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1831
timestamp 1698175906
transform 1 0 206416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1835
timestamp 1698175906
transform 1 0 206864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1844
timestamp 1698175906
transform 1 0 207872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1848
timestamp 1698175906
transform 1 0 208320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1852
timestamp 1698175906
transform 1 0 208768 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1866
timestamp 1698175906
transform 1 0 210336 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1879
timestamp 1698175906
transform 1 0 211792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1883
timestamp 1698175906
transform 1 0 212240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1893
timestamp 1698175906
transform 1 0 213360 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1901
timestamp 1698175906
transform 1 0 214256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1903
timestamp 1698175906
transform 1 0 214480 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1906
timestamp 1698175906
transform 1 0 214816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1912
timestamp 1698175906
transform 1 0 215488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1916
timestamp 1698175906
transform 1 0 215936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1918
timestamp 1698175906
transform 1 0 216160 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1925
timestamp 1698175906
transform 1 0 216944 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1933
timestamp 1698175906
transform 1 0 217840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1937
timestamp 1698175906
transform 1 0 218288 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1940
timestamp 1698175906
transform 1 0 218624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1944
timestamp 1698175906
transform 1 0 219072 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1967
timestamp 1698175906
transform 1 0 221648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1971
timestamp 1698175906
transform 1 0 222096 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1974
timestamp 1698175906
transform 1 0 222432 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1978
timestamp 1698175906
transform 1 0 222880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1980
timestamp 1698175906
transform 1 0 223104 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1989
timestamp 1698175906
transform 1 0 224112 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2005
timestamp 1698175906
transform 1 0 225904 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2008
timestamp 1698175906
transform 1 0 226240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2012
timestamp 1698175906
transform 1 0 226688 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2021
timestamp 1698175906
transform 1 0 227696 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2037
timestamp 1698175906
transform 1 0 229488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2039
timestamp 1698175906
transform 1 0 229712 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2042
timestamp 1698175906
transform 1 0 230048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2044
timestamp 1698175906
transform 1 0 230272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2053
timestamp 1698175906
transform 1 0 231280 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2069
timestamp 1698175906
transform 1 0 233072 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2071
timestamp 1698175906
transform 1 0 233296 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2076
timestamp 1698175906
transform 1 0 233856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2078
timestamp 1698175906
transform 1 0 234080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2085
timestamp 1698175906
transform 1 0 234864 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2101
timestamp 1698175906
transform 1 0 236656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2105
timestamp 1698175906
transform 1 0 237104 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2110
timestamp 1698175906
transform 1 0 237664 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2117
timestamp 1698175906
transform 1 0 238448 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2133
timestamp 1698175906
transform 1 0 240240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2137
timestamp 1698175906
transform 1 0 240688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2139
timestamp 1698175906
transform 1 0 240912 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2150
timestamp 1698175906
transform 1 0 242144 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2166
timestamp 1698175906
transform 1 0 243936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2184
timestamp 1698175906
transform 1 0 245952 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2200
timestamp 1698175906
transform 1 0 247744 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2218
timestamp 1698175906
transform 1 0 249760 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2234
timestamp 1698175906
transform 1 0 251552 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2252
timestamp 1698175906
transform 1 0 253568 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2268
timestamp 1698175906
transform 1 0 255360 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2277
timestamp 1698175906
transform 1 0 256368 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2280
timestamp 1698175906
transform 1 0 256704 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2296
timestamp 1698175906
transform 1 0 258496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2300
timestamp 1698175906
transform 1 0 258944 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2309
timestamp 1698175906
transform 1 0 259952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2311
timestamp 1698175906
transform 1 0 260176 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2314
timestamp 1698175906
transform 1 0 260512 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2330
timestamp 1698175906
transform 1 0 262304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2332
timestamp 1698175906
transform 1 0 262528 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2341
timestamp 1698175906
transform 1 0 263536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2345
timestamp 1698175906
transform 1 0 263984 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2348
timestamp 1698175906
transform 1 0 264320 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2364
timestamp 1698175906
transform 1 0 266112 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2375
timestamp 1698175906
transform 1 0 267344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2379
timestamp 1698175906
transform 1 0 267792 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2382
timestamp 1698175906
transform 1 0 268128 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2390
timestamp 1698175906
transform 1 0 269024 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2394
timestamp 1698175906
transform 1 0 269472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2396
timestamp 1698175906
transform 1 0 269696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2407
timestamp 1698175906
transform 1 0 270928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2411
timestamp 1698175906
transform 1 0 271376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2413
timestamp 1698175906
transform 1 0 271600 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2416
timestamp 1698175906
transform 1 0 271936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2424
timestamp 1698175906
transform 1 0 272832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2428
timestamp 1698175906
transform 1 0 273280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2439
timestamp 1698175906
transform 1 0 274512 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2447
timestamp 1698175906
transform 1 0 275408 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2450
timestamp 1698175906
transform 1 0 275744 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2458
timestamp 1698175906
transform 1 0 276640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2460
timestamp 1698175906
transform 1 0 276864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2471
timestamp 1698175906
transform 1 0 278096 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2479
timestamp 1698175906
transform 1 0 278992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2481
timestamp 1698175906
transform 1 0 279216 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2484
timestamp 1698175906
transform 1 0 279552 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2492
timestamp 1698175906
transform 1 0 280448 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2503
timestamp 1698175906
transform 1 0 281680 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2511
timestamp 1698175906
transform 1 0 282576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2515
timestamp 1698175906
transform 1 0 283024 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2518
timestamp 1698175906
transform 1 0 283360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2522
timestamp 1698175906
transform 1 0 283808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2524
timestamp 1698175906
transform 1 0 284032 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2535
timestamp 1698175906
transform 1 0 285264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2543
timestamp 1698175906
transform 1 0 286160 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2547
timestamp 1698175906
transform 1 0 286608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2549
timestamp 1698175906
transform 1 0 286832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_2552
timestamp 1698175906
transform 1 0 287168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2556
timestamp 1698175906
transform 1 0 287616 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2567
timestamp 1698175906
transform 1 0 288848 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2583
timestamp 1698175906
transform 1 0 290640 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2586
timestamp 1698175906
transform 1 0 290976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2588
timestamp 1698175906
transform 1 0 291200 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2599
timestamp 1698175906
transform 1 0 292432 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2615
timestamp 1698175906
transform 1 0 294224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2617
timestamp 1698175906
transform 1 0 294448 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2620
timestamp 1698175906
transform 1 0 294784 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_88
timestamp 1698175906
transform 1 0 11200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_96
timestamp 1698175906
transform 1 0 12096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_100
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_132
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698175906
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698175906
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_422
timestamp 1698175906
transform 1 0 48608 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_438
timestamp 1698175906
transform 1 0 50400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_440
timestamp 1698175906
transform 1 0 50624 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_443
timestamp 1698175906
transform 1 0 50960 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_459
timestamp 1698175906
transform 1 0 52752 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_467
timestamp 1698175906
transform 1 0 53648 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_471
timestamp 1698175906
transform 1 0 54096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_475
timestamp 1698175906
transform 1 0 54544 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_483
timestamp 1698175906
transform 1 0 55440 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_487
timestamp 1698175906
transform 1 0 55888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1698175906
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_492
timestamp 1698175906
transform 1 0 56448 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_556
timestamp 1698175906
transform 1 0 63616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_562
timestamp 1698175906
transform 1 0 64288 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_594
timestamp 1698175906
transform 1 0 67872 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_610
timestamp 1698175906
transform 1 0 69664 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_618
timestamp 1698175906
transform 1 0 70560 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_632
timestamp 1698175906
transform 1 0 72128 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_648
timestamp 1698175906
transform 1 0 73920 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_652
timestamp 1698175906
transform 1 0 74368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_654
timestamp 1698175906
transform 1 0 74592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_663
timestamp 1698175906
transform 1 0 75600 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_697
timestamp 1698175906
transform 1 0 79408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_699
timestamp 1698175906
transform 1 0 79632 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_702
timestamp 1698175906
transform 1 0 79968 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_767
timestamp 1698175906
transform 1 0 87248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_769
timestamp 1698175906
transform 1 0 87472 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_798
timestamp 1698175906
transform 1 0 90720 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_831
timestamp 1698175906
transform 1 0 94416 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_839
timestamp 1698175906
transform 1 0 95312 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_842
timestamp 1698175906
transform 1 0 95648 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_854
timestamp 1698175906
transform 1 0 96992 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_886
timestamp 1698175906
transform 1 0 100576 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_902
timestamp 1698175906
transform 1 0 102368 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_912
timestamp 1698175906
transform 1 0 103488 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_976
timestamp 1698175906
transform 1 0 110656 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_982
timestamp 1698175906
transform 1 0 111328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_984
timestamp 1698175906
transform 1 0 111552 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_987
timestamp 1698175906
transform 1 0 111888 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1003
timestamp 1698175906
transform 1 0 113680 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1011
timestamp 1698175906
transform 1 0 114576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1015
timestamp 1698175906
transform 1 0 115024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_1019
timestamp 1698175906
transform 1 0 115472 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1035
timestamp 1698175906
transform 1 0 117264 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1043
timestamp 1698175906
transform 1 0 118160 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1047
timestamp 1698175906
transform 1 0 118608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1049
timestamp 1698175906
transform 1 0 118832 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_1052
timestamp 1698175906
transform 1 0 119168 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1068
timestamp 1698175906
transform 1 0 120960 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1076
timestamp 1698175906
transform 1 0 121856 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1080
timestamp 1698175906
transform 1 0 122304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_1084
timestamp 1698175906
transform 1 0 122752 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1116
timestamp 1698175906
transform 1 0 126336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1122
timestamp 1698175906
transform 1 0 127008 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1186
timestamp 1698175906
transform 1 0 134176 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1192
timestamp 1698175906
transform 1 0 134848 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1256
timestamp 1698175906
transform 1 0 142016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1262
timestamp 1698175906
transform 1 0 142688 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1326
timestamp 1698175906
transform 1 0 149856 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1332
timestamp 1698175906
transform 1 0 150528 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1396
timestamp 1698175906
transform 1 0 157696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1402
timestamp 1698175906
transform 1 0 158368 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1466
timestamp 1698175906
transform 1 0 165536 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1472
timestamp 1698175906
transform 1 0 166208 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1536
timestamp 1698175906
transform 1 0 173376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1542
timestamp 1698175906
transform 1 0 174048 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1606
timestamp 1698175906
transform 1 0 181216 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1612
timestamp 1698175906
transform 1 0 181888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1670
timestamp 1698175906
transform 1 0 188384 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1729
timestamp 1698175906
transform 1 0 194992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1733
timestamp 1698175906
transform 1 0 195440 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1737
timestamp 1698175906
transform 1 0 195888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1739
timestamp 1698175906
transform 1 0 196112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1815
timestamp 1698175906
transform 1 0 204624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1819
timestamp 1698175906
transform 1 0 205072 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1887
timestamp 1698175906
transform 1 0 212688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1889
timestamp 1698175906
transform 1 0 212912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1892
timestamp 1698175906
transform 1 0 213248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1900
timestamp 1698175906
transform 1 0 214144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1904
timestamp 1698175906
transform 1 0 214592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1914
timestamp 1698175906
transform 1 0 215712 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1918
timestamp 1698175906
transform 1 0 216160 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1932
timestamp 1698175906
transform 1 0 217728 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1936
timestamp 1698175906
transform 1 0 218176 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1944
timestamp 1698175906
transform 1 0 219072 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1955
timestamp 1698175906
transform 1 0 220304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1957
timestamp 1698175906
transform 1 0 220528 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1973
timestamp 1698175906
transform 1 0 222320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1983
timestamp 1698175906
transform 1 0 223440 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_1987
timestamp 1698175906
transform 1 0 223888 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_2019
timestamp 1698175906
transform 1 0 227472 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_2027
timestamp 1698175906
transform 1 0 228368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_2029
timestamp 1698175906
transform 1 0 228592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2032
timestamp 1698175906
transform 1 0 228928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2096
timestamp 1698175906
transform 1 0 236096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2102
timestamp 1698175906
transform 1 0 236768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2166
timestamp 1698175906
transform 1 0 243936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2172
timestamp 1698175906
transform 1 0 244608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2236
timestamp 1698175906
transform 1 0 251776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2242
timestamp 1698175906
transform 1 0 252448 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2306
timestamp 1698175906
transform 1 0 259616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2312
timestamp 1698175906
transform 1 0 260288 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2376
timestamp 1698175906
transform 1 0 267456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2382
timestamp 1698175906
transform 1 0 268128 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2446
timestamp 1698175906
transform 1 0 275296 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2452
timestamp 1698175906
transform 1 0 275968 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2516
timestamp 1698175906
transform 1 0 283136 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2522
timestamp 1698175906
transform 1 0 283808 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2586
timestamp 1698175906
transform 1 0 290976 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_2592
timestamp 1698175906
transform 1 0 291648 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_2624
timestamp 1698175906
transform 1 0 295232 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_2640
timestamp 1698175906
transform 1 0 297024 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2648
timestamp 1698175906
transform 1 0 297920 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698175906
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698175906
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698175906
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_457
timestamp 1698175906
transform 1 0 52528 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_521
timestamp 1698175906
transform 1 0 59696 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_527
timestamp 1698175906
transform 1 0 60368 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_591
timestamp 1698175906
transform 1 0 67536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_597
timestamp 1698175906
transform 1 0 68208 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_661
timestamp 1698175906
transform 1 0 75376 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_667
timestamp 1698175906
transform 1 0 76048 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_731
timestamp 1698175906
transform 1 0 83216 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_737
timestamp 1698175906
transform 1 0 83888 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_801
timestamp 1698175906
transform 1 0 91056 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_807
timestamp 1698175906
transform 1 0 91728 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_825
timestamp 1698175906
transform 1 0 93744 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_857
timestamp 1698175906
transform 1 0 97328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_873
timestamp 1698175906
transform 1 0 99120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_877
timestamp 1698175906
transform 1 0 99568 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_941
timestamp 1698175906
transform 1 0 106736 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_947
timestamp 1698175906
transform 1 0 107408 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1011
timestamp 1698175906
transform 1 0 114576 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1017
timestamp 1698175906
transform 1 0 115248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1081
timestamp 1698175906
transform 1 0 122416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1087
timestamp 1698175906
transform 1 0 123088 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1151
timestamp 1698175906
transform 1 0 130256 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1157
timestamp 1698175906
transform 1 0 130928 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1221
timestamp 1698175906
transform 1 0 138096 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1227
timestamp 1698175906
transform 1 0 138768 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1291
timestamp 1698175906
transform 1 0 145936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1297
timestamp 1698175906
transform 1 0 146608 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1361
timestamp 1698175906
transform 1 0 153776 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1367
timestamp 1698175906
transform 1 0 154448 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1431
timestamp 1698175906
transform 1 0 161616 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1437
timestamp 1698175906
transform 1 0 162288 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1501
timestamp 1698175906
transform 1 0 169456 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1507
timestamp 1698175906
transform 1 0 170128 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1571
timestamp 1698175906
transform 1 0 177296 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_1577
timestamp 1698175906
transform 1 0 177968 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1609
timestamp 1698175906
transform 1 0 181552 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1656
timestamp 1698175906
transform 1 0 186816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1727
timestamp 1698175906
transform 1 0 194768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1731
timestamp 1698175906
transform 1 0 195216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1735
timestamp 1698175906
transform 1 0 195664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1737
timestamp 1698175906
transform 1 0 195888 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1787
timestamp 1698175906
transform 1 0 201488 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1821
timestamp 1698175906
transform 1 0 205296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1823
timestamp 1698175906
transform 1 0 205520 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1842
timestamp 1698175906
transform 1 0 207648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1846
timestamp 1698175906
transform 1 0 208096 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1874
timestamp 1698175906
transform 1 0 211232 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1876
timestamp 1698175906
transform 1 0 211456 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1890
timestamp 1698175906
transform 1 0 213024 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1898
timestamp 1698175906
transform 1 0 213920 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1921
timestamp 1698175906
transform 1 0 216496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1946
timestamp 1698175906
transform 1 0 219296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1948
timestamp 1698175906
transform 1 0 219520 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1971
timestamp 1698175906
transform 1 0 222096 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1991
timestamp 1698175906
transform 1 0 224336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1997
timestamp 1698175906
transform 1 0 225008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_2061
timestamp 1698175906
transform 1 0 232176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_2067
timestamp 1698175906
transform 1 0 232848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_2131
timestamp 1698175906
transform 1 0 240016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_2137
timestamp 1698175906
transform 1 0 240688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_2201
timestamp 1698175906
transform 1 0 247856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_2207
timestamp 1698175906
transform 1 0 248528 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_2271
timestamp 1698175906
transform 1 0 255696 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_2277
timestamp 1698175906
transform 1 0 256368 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_2341
timestamp 1698175906
transform 1 0 263536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_2347
timestamp 1698175906
transform 1 0 264208 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_2411
timestamp 1698175906
transform 1 0 271376 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_2417
timestamp 1698175906
transform 1 0 272048 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_2481
timestamp 1698175906
transform 1 0 279216 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_2487
timestamp 1698175906
transform 1 0 279888 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_2551
timestamp 1698175906
transform 1 0 287056 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_2557
timestamp 1698175906
transform 1 0 287728 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_2621
timestamp 1698175906
transform 1 0 294896 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_2627
timestamp 1698175906
transform 1 0 295568 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_2643
timestamp 1698175906
transform 1 0 297360 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_2651
timestamp 1698175906
transform 1 0 298256 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698175906
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698175906
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698175906
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698175906
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_492
timestamp 1698175906
transform 1 0 56448 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_556
timestamp 1698175906
transform 1 0 63616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_562
timestamp 1698175906
transform 1 0 64288 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_626
timestamp 1698175906
transform 1 0 71456 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_632
timestamp 1698175906
transform 1 0 72128 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_696
timestamp 1698175906
transform 1 0 79296 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_702
timestamp 1698175906
transform 1 0 79968 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_766
timestamp 1698175906
transform 1 0 87136 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_772
timestamp 1698175906
transform 1 0 87808 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_836
timestamp 1698175906
transform 1 0 94976 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_842
timestamp 1698175906
transform 1 0 95648 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_906
timestamp 1698175906
transform 1 0 102816 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_912
timestamp 1698175906
transform 1 0 103488 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_976
timestamp 1698175906
transform 1 0 110656 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_982
timestamp 1698175906
transform 1 0 111328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1046
timestamp 1698175906
transform 1 0 118496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1052
timestamp 1698175906
transform 1 0 119168 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1116
timestamp 1698175906
transform 1 0 126336 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1122
timestamp 1698175906
transform 1 0 127008 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1186
timestamp 1698175906
transform 1 0 134176 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1192
timestamp 1698175906
transform 1 0 134848 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1256
timestamp 1698175906
transform 1 0 142016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1262
timestamp 1698175906
transform 1 0 142688 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1326
timestamp 1698175906
transform 1 0 149856 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1332
timestamp 1698175906
transform 1 0 150528 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1396
timestamp 1698175906
transform 1 0 157696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1402
timestamp 1698175906
transform 1 0 158368 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1466
timestamp 1698175906
transform 1 0 165536 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1472
timestamp 1698175906
transform 1 0 166208 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1536
timestamp 1698175906
transform 1 0 173376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1542
timestamp 1698175906
transform 1 0 174048 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1606
timestamp 1698175906
transform 1 0 181216 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_1612
timestamp 1698175906
transform 1 0 181888 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1620
timestamp 1698175906
transform 1 0 182784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1664
timestamp 1698175906
transform 1 0 187712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1668
timestamp 1698175906
transform 1 0 188160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1696
timestamp 1698175906
transform 1 0 191296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1702
timestamp 1698175906
transform 1 0 191968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1736
timestamp 1698175906
transform 1 0 195776 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1747
timestamp 1698175906
transform 1 0 197008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1749
timestamp 1698175906
transform 1 0 197232 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1807
timestamp 1698175906
transform 1 0 203728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1811
timestamp 1698175906
transform 1 0 204176 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1839
timestamp 1698175906
transform 1 0 207312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1843
timestamp 1698175906
transform 1 0 207760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1847
timestamp 1698175906
transform 1 0 208208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1851
timestamp 1698175906
transform 1 0 208656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1855
timestamp 1698175906
transform 1 0 209104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1857
timestamp 1698175906
transform 1 0 209328 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_1879
timestamp 1698175906
transform 1 0 211792 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1887
timestamp 1698175906
transform 1 0 212688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1889
timestamp 1698175906
transform 1 0 212912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_1892
timestamp 1698175906
transform 1 0 213248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1900
timestamp 1698175906
transform 1 0 214144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1902
timestamp 1698175906
transform 1 0 214368 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1909
timestamp 1698175906
transform 1 0 215152 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1913
timestamp 1698175906
transform 1 0 215600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1924
timestamp 1698175906
transform 1 0 216832 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_1928
timestamp 1698175906
transform 1 0 217280 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1944
timestamp 1698175906
transform 1 0 219072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1946
timestamp 1698175906
transform 1 0 219296 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_1949
timestamp 1698175906
transform 1 0 219632 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1957
timestamp 1698175906
transform 1 0 220528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1959
timestamp 1698175906
transform 1 0 220752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_1962
timestamp 1698175906
transform 1 0 221088 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1978
timestamp 1698175906
transform 1 0 222880 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1982
timestamp 1698175906
transform 1 0 223328 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_1985
timestamp 1698175906
transform 1 0 223664 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_2017
timestamp 1698175906
transform 1 0 227248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2025
timestamp 1698175906
transform 1 0 228144 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_2029
timestamp 1698175906
transform 1 0 228592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2032
timestamp 1698175906
transform 1 0 228928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2096
timestamp 1698175906
transform 1 0 236096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2102
timestamp 1698175906
transform 1 0 236768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2166
timestamp 1698175906
transform 1 0 243936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2172
timestamp 1698175906
transform 1 0 244608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2236
timestamp 1698175906
transform 1 0 251776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2242
timestamp 1698175906
transform 1 0 252448 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2306
timestamp 1698175906
transform 1 0 259616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2312
timestamp 1698175906
transform 1 0 260288 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2376
timestamp 1698175906
transform 1 0 267456 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2382
timestamp 1698175906
transform 1 0 268128 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2446
timestamp 1698175906
transform 1 0 275296 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2452
timestamp 1698175906
transform 1 0 275968 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2516
timestamp 1698175906
transform 1 0 283136 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2522
timestamp 1698175906
transform 1 0 283808 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2586
timestamp 1698175906
transform 1 0 290976 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_2592
timestamp 1698175906
transform 1 0 291648 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_2624
timestamp 1698175906
transform 1 0 295232 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_2640
timestamp 1698175906
transform 1 0 297024 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2648
timestamp 1698175906
transform 1 0 297920 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698175906
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698175906
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698175906
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_457
timestamp 1698175906
transform 1 0 52528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_521
timestamp 1698175906
transform 1 0 59696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_527
timestamp 1698175906
transform 1 0 60368 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_591
timestamp 1698175906
transform 1 0 67536 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_597
timestamp 1698175906
transform 1 0 68208 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_661
timestamp 1698175906
transform 1 0 75376 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_667
timestamp 1698175906
transform 1 0 76048 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_731
timestamp 1698175906
transform 1 0 83216 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_737
timestamp 1698175906
transform 1 0 83888 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_801
timestamp 1698175906
transform 1 0 91056 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_807
timestamp 1698175906
transform 1 0 91728 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_871
timestamp 1698175906
transform 1 0 98896 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_877
timestamp 1698175906
transform 1 0 99568 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_941
timestamp 1698175906
transform 1 0 106736 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_947
timestamp 1698175906
transform 1 0 107408 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1011
timestamp 1698175906
transform 1 0 114576 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1017
timestamp 1698175906
transform 1 0 115248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1081
timestamp 1698175906
transform 1 0 122416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1087
timestamp 1698175906
transform 1 0 123088 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1151
timestamp 1698175906
transform 1 0 130256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1157
timestamp 1698175906
transform 1 0 130928 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1221
timestamp 1698175906
transform 1 0 138096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1227
timestamp 1698175906
transform 1 0 138768 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1291
timestamp 1698175906
transform 1 0 145936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1297
timestamp 1698175906
transform 1 0 146608 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1361
timestamp 1698175906
transform 1 0 153776 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1367
timestamp 1698175906
transform 1 0 154448 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1431
timestamp 1698175906
transform 1 0 161616 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1437
timestamp 1698175906
transform 1 0 162288 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1501
timestamp 1698175906
transform 1 0 169456 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1507
timestamp 1698175906
transform 1 0 170128 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1571
timestamp 1698175906
transform 1 0 177296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_1577
timestamp 1698175906
transform 1 0 177968 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_1609
timestamp 1698175906
transform 1 0 181552 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1625
timestamp 1698175906
transform 1 0 183344 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1629
timestamp 1698175906
transform 1 0 183792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_1637
timestamp 1698175906
transform 1 0 184688 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1647
timestamp 1698175906
transform 1 0 185808 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1651
timestamp 1698175906
transform 1 0 186256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1653
timestamp 1698175906
transform 1 0 186480 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1656
timestamp 1698175906
transform 1 0 186816 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1707
timestamp 1698175906
transform 1 0 192528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1711
timestamp 1698175906
transform 1 0 192976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1717
timestamp 1698175906
transform 1 0 193648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1721
timestamp 1698175906
transform 1 0 194096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_1725
timestamp 1698175906
transform 1 0 194544 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1733
timestamp 1698175906
transform 1 0 195440 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1735
timestamp 1698175906
transform 1 0 195664 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1834
timestamp 1698175906
transform 1 0 206752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1838
timestamp 1698175906
transform 1 0 207200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1842
timestamp 1698175906
transform 1 0 207648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_1846
timestamp 1698175906
transform 1 0 208096 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1854
timestamp 1698175906
transform 1 0 208992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_1857
timestamp 1698175906
transform 1 0 209328 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1889
timestamp 1698175906
transform 1 0 212912 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1893
timestamp 1698175906
transform 1 0 213360 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_1900
timestamp 1698175906
transform 1 0 214144 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_1916
timestamp 1698175906
transform 1 0 215936 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1924
timestamp 1698175906
transform 1 0 216832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1941
timestamp 1698175906
transform 1 0 218736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_1945
timestamp 1698175906
transform 1 0 219184 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_1977
timestamp 1698175906
transform 1 0 222768 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1993
timestamp 1698175906
transform 1 0 224560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1997
timestamp 1698175906
transform 1 0 225008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2061
timestamp 1698175906
transform 1 0 232176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_2067
timestamp 1698175906
transform 1 0 232848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2131
timestamp 1698175906
transform 1 0 240016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_2137
timestamp 1698175906
transform 1 0 240688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2201
timestamp 1698175906
transform 1 0 247856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_2207
timestamp 1698175906
transform 1 0 248528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2271
timestamp 1698175906
transform 1 0 255696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_2277
timestamp 1698175906
transform 1 0 256368 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2341
timestamp 1698175906
transform 1 0 263536 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_2347
timestamp 1698175906
transform 1 0 264208 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2411
timestamp 1698175906
transform 1 0 271376 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_2417
timestamp 1698175906
transform 1 0 272048 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2481
timestamp 1698175906
transform 1 0 279216 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_2487
timestamp 1698175906
transform 1 0 279888 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2551
timestamp 1698175906
transform 1 0 287056 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_2557
timestamp 1698175906
transform 1 0 287728 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2621
timestamp 1698175906
transform 1 0 294896 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_2627
timestamp 1698175906
transform 1 0 295568 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_2643
timestamp 1698175906
transform 1 0 297360 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_2651
timestamp 1698175906
transform 1 0 298256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698175906
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698175906
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698175906
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698175906
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_492
timestamp 1698175906
transform 1 0 56448 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_556
timestamp 1698175906
transform 1 0 63616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_562
timestamp 1698175906
transform 1 0 64288 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_626
timestamp 1698175906
transform 1 0 71456 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_632
timestamp 1698175906
transform 1 0 72128 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_696
timestamp 1698175906
transform 1 0 79296 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_702
timestamp 1698175906
transform 1 0 79968 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_766
timestamp 1698175906
transform 1 0 87136 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_772
timestamp 1698175906
transform 1 0 87808 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_836
timestamp 1698175906
transform 1 0 94976 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_842
timestamp 1698175906
transform 1 0 95648 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_906
timestamp 1698175906
transform 1 0 102816 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_912
timestamp 1698175906
transform 1 0 103488 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_976
timestamp 1698175906
transform 1 0 110656 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_982
timestamp 1698175906
transform 1 0 111328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1046
timestamp 1698175906
transform 1 0 118496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1052
timestamp 1698175906
transform 1 0 119168 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1116
timestamp 1698175906
transform 1 0 126336 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1122
timestamp 1698175906
transform 1 0 127008 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1186
timestamp 1698175906
transform 1 0 134176 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1192
timestamp 1698175906
transform 1 0 134848 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1256
timestamp 1698175906
transform 1 0 142016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1262
timestamp 1698175906
transform 1 0 142688 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1326
timestamp 1698175906
transform 1 0 149856 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1332
timestamp 1698175906
transform 1 0 150528 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1396
timestamp 1698175906
transform 1 0 157696 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1402
timestamp 1698175906
transform 1 0 158368 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1466
timestamp 1698175906
transform 1 0 165536 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1472
timestamp 1698175906
transform 1 0 166208 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1536
timestamp 1698175906
transform 1 0 173376 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1542
timestamp 1698175906
transform 1 0 174048 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1606
timestamp 1698175906
transform 1 0 181216 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_1612
timestamp 1698175906
transform 1 0 181888 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_1628
timestamp 1698175906
transform 1 0 183680 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1636
timestamp 1698175906
transform 1 0 184576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_1638
timestamp 1698175906
transform 1 0 184800 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1692
timestamp 1698175906
transform 1 0 190848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1696
timestamp 1698175906
transform 1 0 191296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1700
timestamp 1698175906
transform 1 0 191744 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1736
timestamp 1698175906
transform 1 0 195776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_1740
timestamp 1698175906
transform 1 0 196224 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1748
timestamp 1698175906
transform 1 0 197120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1762
timestamp 1698175906
transform 1 0 198688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_1764
timestamp 1698175906
transform 1 0 198912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1767
timestamp 1698175906
transform 1 0 199248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1811
timestamp 1698175906
transform 1 0 204176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_1813
timestamp 1698175906
transform 1 0 204400 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1828
timestamp 1698175906
transform 1 0 206080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_1832
timestamp 1698175906
transform 1 0 206528 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_1841
timestamp 1698175906
transform 1 0 207536 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_1857
timestamp 1698175906
transform 1 0 209328 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1886
timestamp 1698175906
transform 1 0 212576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1892
timestamp 1698175906
transform 1 0 213248 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1896
timestamp 1698175906
transform 1 0 213696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_1906
timestamp 1698175906
transform 1 0 214816 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_1925
timestamp 1698175906
transform 1 0 216944 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1957
timestamp 1698175906
transform 1 0 220528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_1959
timestamp 1698175906
transform 1 0 220752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1962
timestamp 1698175906
transform 1 0 221088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2026
timestamp 1698175906
transform 1 0 228256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2032
timestamp 1698175906
transform 1 0 228928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2096
timestamp 1698175906
transform 1 0 236096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2102
timestamp 1698175906
transform 1 0 236768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2166
timestamp 1698175906
transform 1 0 243936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2172
timestamp 1698175906
transform 1 0 244608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2236
timestamp 1698175906
transform 1 0 251776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2242
timestamp 1698175906
transform 1 0 252448 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2306
timestamp 1698175906
transform 1 0 259616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2312
timestamp 1698175906
transform 1 0 260288 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2376
timestamp 1698175906
transform 1 0 267456 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2382
timestamp 1698175906
transform 1 0 268128 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2446
timestamp 1698175906
transform 1 0 275296 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2452
timestamp 1698175906
transform 1 0 275968 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2516
timestamp 1698175906
transform 1 0 283136 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2522
timestamp 1698175906
transform 1 0 283808 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2586
timestamp 1698175906
transform 1 0 290976 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_2592
timestamp 1698175906
transform 1 0 291648 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_2624
timestamp 1698175906
transform 1 0 295232 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_2640
timestamp 1698175906
transform 1 0 297024 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2648
timestamp 1698175906
transform 1 0 297920 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698175906
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698175906
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698175906
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_457
timestamp 1698175906
transform 1 0 52528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_521
timestamp 1698175906
transform 1 0 59696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_527
timestamp 1698175906
transform 1 0 60368 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_591
timestamp 1698175906
transform 1 0 67536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_597
timestamp 1698175906
transform 1 0 68208 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_661
timestamp 1698175906
transform 1 0 75376 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_667
timestamp 1698175906
transform 1 0 76048 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_731
timestamp 1698175906
transform 1 0 83216 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_737
timestamp 1698175906
transform 1 0 83888 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_801
timestamp 1698175906
transform 1 0 91056 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_807
timestamp 1698175906
transform 1 0 91728 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_871
timestamp 1698175906
transform 1 0 98896 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_877
timestamp 1698175906
transform 1 0 99568 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_941
timestamp 1698175906
transform 1 0 106736 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_947
timestamp 1698175906
transform 1 0 107408 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1011
timestamp 1698175906
transform 1 0 114576 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1017
timestamp 1698175906
transform 1 0 115248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1081
timestamp 1698175906
transform 1 0 122416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1087
timestamp 1698175906
transform 1 0 123088 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1151
timestamp 1698175906
transform 1 0 130256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1157
timestamp 1698175906
transform 1 0 130928 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1221
timestamp 1698175906
transform 1 0 138096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1227
timestamp 1698175906
transform 1 0 138768 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1291
timestamp 1698175906
transform 1 0 145936 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1297
timestamp 1698175906
transform 1 0 146608 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1361
timestamp 1698175906
transform 1 0 153776 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1367
timestamp 1698175906
transform 1 0 154448 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1431
timestamp 1698175906
transform 1 0 161616 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1437
timestamp 1698175906
transform 1 0 162288 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1501
timestamp 1698175906
transform 1 0 169456 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1507
timestamp 1698175906
transform 1 0 170128 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1571
timestamp 1698175906
transform 1 0 177296 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1577
timestamp 1698175906
transform 1 0 177968 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1641
timestamp 1698175906
transform 1 0 185136 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1647
timestamp 1698175906
transform 1 0 185808 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1655
timestamp 1698175906
transform 1 0 186704 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1659
timestamp 1698175906
transform 1 0 187152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1674
timestamp 1698175906
transform 1 0 188832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1685
timestamp 1698175906
transform 1 0 190064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1689
timestamp 1698175906
transform 1 0 190512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_1693
timestamp 1698175906
transform 1 0 190960 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1709
timestamp 1698175906
transform 1 0 192752 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1713
timestamp 1698175906
transform 1 0 193200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_1717
timestamp 1698175906
transform 1 0 193648 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1749
timestamp 1698175906
transform 1 0 197232 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1757
timestamp 1698175906
transform 1 0 198128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1761
timestamp 1698175906
transform 1 0 198576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1763
timestamp 1698175906
transform 1 0 198800 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1766
timestamp 1698175906
transform 1 0 199136 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1776
timestamp 1698175906
transform 1 0 200256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1778
timestamp 1698175906
transform 1 0 200480 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1821
timestamp 1698175906
transform 1 0 205296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1851
timestamp 1698175906
transform 1 0 208656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1857
timestamp 1698175906
transform 1 0 209328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1859
timestamp 1698175906
transform 1 0 209552 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1886
timestamp 1698175906
transform 1 0 212576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1890
timestamp 1698175906
transform 1 0 213024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_1894
timestamp 1698175906
transform 1 0 213472 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1910
timestamp 1698175906
transform 1 0 215264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1918
timestamp 1698175906
transform 1 0 216160 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1922
timestamp 1698175906
transform 1 0 216608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1924
timestamp 1698175906
transform 1 0 216832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1927
timestamp 1698175906
transform 1 0 217168 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_1934
timestamp 1698175906
transform 1 0 217952 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1950
timestamp 1698175906
transform 1 0 219744 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1967
timestamp 1698175906
transform 1 0 221648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_1971
timestamp 1698175906
transform 1 0 222096 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1987
timestamp 1698175906
transform 1 0 223888 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1997
timestamp 1698175906
transform 1 0 225008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2061
timestamp 1698175906
transform 1 0 232176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_2067
timestamp 1698175906
transform 1 0 232848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2131
timestamp 1698175906
transform 1 0 240016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_2137
timestamp 1698175906
transform 1 0 240688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2201
timestamp 1698175906
transform 1 0 247856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_2207
timestamp 1698175906
transform 1 0 248528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2271
timestamp 1698175906
transform 1 0 255696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_2277
timestamp 1698175906
transform 1 0 256368 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2341
timestamp 1698175906
transform 1 0 263536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_2347
timestamp 1698175906
transform 1 0 264208 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2411
timestamp 1698175906
transform 1 0 271376 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_2417
timestamp 1698175906
transform 1 0 272048 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2481
timestamp 1698175906
transform 1 0 279216 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_2487
timestamp 1698175906
transform 1 0 279888 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2551
timestamp 1698175906
transform 1 0 287056 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_2557
timestamp 1698175906
transform 1 0 287728 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2621
timestamp 1698175906
transform 1 0 294896 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_2627
timestamp 1698175906
transform 1 0 295568 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_2643
timestamp 1698175906
transform 1 0 297360 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_2651
timestamp 1698175906
transform 1 0 298256 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698175906
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698175906
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698175906
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698175906
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_492
timestamp 1698175906
transform 1 0 56448 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_556
timestamp 1698175906
transform 1 0 63616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_562
timestamp 1698175906
transform 1 0 64288 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_626
timestamp 1698175906
transform 1 0 71456 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_632
timestamp 1698175906
transform 1 0 72128 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_696
timestamp 1698175906
transform 1 0 79296 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_702
timestamp 1698175906
transform 1 0 79968 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_766
timestamp 1698175906
transform 1 0 87136 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_772
timestamp 1698175906
transform 1 0 87808 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_836
timestamp 1698175906
transform 1 0 94976 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_842
timestamp 1698175906
transform 1 0 95648 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_906
timestamp 1698175906
transform 1 0 102816 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_912
timestamp 1698175906
transform 1 0 103488 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_976
timestamp 1698175906
transform 1 0 110656 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_982
timestamp 1698175906
transform 1 0 111328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1046
timestamp 1698175906
transform 1 0 118496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1052
timestamp 1698175906
transform 1 0 119168 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1116
timestamp 1698175906
transform 1 0 126336 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1122
timestamp 1698175906
transform 1 0 127008 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1186
timestamp 1698175906
transform 1 0 134176 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1192
timestamp 1698175906
transform 1 0 134848 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1256
timestamp 1698175906
transform 1 0 142016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1262
timestamp 1698175906
transform 1 0 142688 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1326
timestamp 1698175906
transform 1 0 149856 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1332
timestamp 1698175906
transform 1 0 150528 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1396
timestamp 1698175906
transform 1 0 157696 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1402
timestamp 1698175906
transform 1 0 158368 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1466
timestamp 1698175906
transform 1 0 165536 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1472
timestamp 1698175906
transform 1 0 166208 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1536
timestamp 1698175906
transform 1 0 173376 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1542
timestamp 1698175906
transform 1 0 174048 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1606
timestamp 1698175906
transform 1 0 181216 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_1612
timestamp 1698175906
transform 1 0 181888 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_1644
timestamp 1698175906
transform 1 0 185472 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_1660
timestamp 1698175906
transform 1 0 187264 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1668
timestamp 1698175906
transform 1 0 188160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1672
timestamp 1698175906
transform 1 0 188608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1676
timestamp 1698175906
transform 1 0 189056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_1682
timestamp 1698175906
transform 1 0 189728 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1698
timestamp 1698175906
transform 1 0 191520 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1702
timestamp 1698175906
transform 1 0 191968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1736
timestamp 1698175906
transform 1 0 195776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_1740
timestamp 1698175906
transform 1 0 196224 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1748
timestamp 1698175906
transform 1 0 197120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_1752
timestamp 1698175906
transform 1 0 197568 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1792
timestamp 1698175906
transform 1 0 202048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1796
timestamp 1698175906
transform 1 0 202496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1804
timestamp 1698175906
transform 1 0 203392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_1808
timestamp 1698175906
transform 1 0 203840 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1816
timestamp 1698175906
transform 1 0 204736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1822
timestamp 1698175906
transform 1 0 205408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_1832
timestamp 1698175906
transform 1 0 206528 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1840
timestamp 1698175906
transform 1 0 207424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_1848
timestamp 1698175906
transform 1 0 208320 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_1900
timestamp 1698175906
transform 1 0 214144 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1916
timestamp 1698175906
transform 1 0 215936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1929
timestamp 1698175906
transform 1 0 217392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1946
timestamp 1698175906
transform 1 0 219296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_1950
timestamp 1698175906
transform 1 0 219744 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1971
timestamp 1698175906
transform 1 0 222096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_1975
timestamp 1698175906
transform 1 0 222544 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2007
timestamp 1698175906
transform 1 0 226128 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2023
timestamp 1698175906
transform 1 0 227920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_2027
timestamp 1698175906
transform 1 0 228368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_2029
timestamp 1698175906
transform 1 0 228592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2032
timestamp 1698175906
transform 1 0 228928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2096
timestamp 1698175906
transform 1 0 236096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2102
timestamp 1698175906
transform 1 0 236768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2166
timestamp 1698175906
transform 1 0 243936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2172
timestamp 1698175906
transform 1 0 244608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2236
timestamp 1698175906
transform 1 0 251776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2242
timestamp 1698175906
transform 1 0 252448 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2306
timestamp 1698175906
transform 1 0 259616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2312
timestamp 1698175906
transform 1 0 260288 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2376
timestamp 1698175906
transform 1 0 267456 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2382
timestamp 1698175906
transform 1 0 268128 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2446
timestamp 1698175906
transform 1 0 275296 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2452
timestamp 1698175906
transform 1 0 275968 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2516
timestamp 1698175906
transform 1 0 283136 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2522
timestamp 1698175906
transform 1 0 283808 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2586
timestamp 1698175906
transform 1 0 290976 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2592
timestamp 1698175906
transform 1 0 291648 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2624
timestamp 1698175906
transform 1 0 295232 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_2640
timestamp 1698175906
transform 1 0 297024 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2648
timestamp 1698175906
transform 1 0 297920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698175906
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698175906
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698175906
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_457
timestamp 1698175906
transform 1 0 52528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_521
timestamp 1698175906
transform 1 0 59696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_527
timestamp 1698175906
transform 1 0 60368 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_591
timestamp 1698175906
transform 1 0 67536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_597
timestamp 1698175906
transform 1 0 68208 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_661
timestamp 1698175906
transform 1 0 75376 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_667
timestamp 1698175906
transform 1 0 76048 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_731
timestamp 1698175906
transform 1 0 83216 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_737
timestamp 1698175906
transform 1 0 83888 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_801
timestamp 1698175906
transform 1 0 91056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_807
timestamp 1698175906
transform 1 0 91728 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_871
timestamp 1698175906
transform 1 0 98896 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_877
timestamp 1698175906
transform 1 0 99568 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_941
timestamp 1698175906
transform 1 0 106736 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_947
timestamp 1698175906
transform 1 0 107408 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1011
timestamp 1698175906
transform 1 0 114576 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1017
timestamp 1698175906
transform 1 0 115248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1081
timestamp 1698175906
transform 1 0 122416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1087
timestamp 1698175906
transform 1 0 123088 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1151
timestamp 1698175906
transform 1 0 130256 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1157
timestamp 1698175906
transform 1 0 130928 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1221
timestamp 1698175906
transform 1 0 138096 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1227
timestamp 1698175906
transform 1 0 138768 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1291
timestamp 1698175906
transform 1 0 145936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1297
timestamp 1698175906
transform 1 0 146608 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1361
timestamp 1698175906
transform 1 0 153776 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1367
timestamp 1698175906
transform 1 0 154448 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1431
timestamp 1698175906
transform 1 0 161616 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1437
timestamp 1698175906
transform 1 0 162288 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1501
timestamp 1698175906
transform 1 0 169456 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1507
timestamp 1698175906
transform 1 0 170128 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1571
timestamp 1698175906
transform 1 0 177296 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1577
timestamp 1698175906
transform 1 0 177968 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1641
timestamp 1698175906
transform 1 0 185136 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1647
timestamp 1698175906
transform 1 0 185808 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1711
timestamp 1698175906
transform 1 0 192976 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_1717
timestamp 1698175906
transform 1 0 193648 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_1749
timestamp 1698175906
transform 1 0 197232 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1765
timestamp 1698175906
transform 1 0 199024 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1768
timestamp 1698175906
transform 1 0 199360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1772
timestamp 1698175906
transform 1 0 199808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1776
timestamp 1698175906
transform 1 0 200256 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1780
timestamp 1698175906
transform 1 0 200704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1784
timestamp 1698175906
transform 1 0 201152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1787
timestamp 1698175906
transform 1 0 201488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1851
timestamp 1698175906
transform 1 0 208656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_1857
timestamp 1698175906
transform 1 0 209328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1865
timestamp 1698175906
transform 1 0 210224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1869
timestamp 1698175906
transform 1 0 210672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_1888
timestamp 1698175906
transform 1 0 212800 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1920
timestamp 1698175906
transform 1 0 216384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1924
timestamp 1698175906
transform 1 0 216832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1927
timestamp 1698175906
transform 1 0 217168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_1931
timestamp 1698175906
transform 1 0 217616 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_1947
timestamp 1698175906
transform 1 0 219408 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1955
timestamp 1698175906
transform 1 0 220304 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1959
timestamp 1698175906
transform 1 0 220752 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_1962
timestamp 1698175906
transform 1 0 221088 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1994
timestamp 1698175906
transform 1 0 224672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1997
timestamp 1698175906
transform 1 0 225008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2061
timestamp 1698175906
transform 1 0 232176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_2067
timestamp 1698175906
transform 1 0 232848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2131
timestamp 1698175906
transform 1 0 240016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_2137
timestamp 1698175906
transform 1 0 240688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2201
timestamp 1698175906
transform 1 0 247856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_2207
timestamp 1698175906
transform 1 0 248528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2271
timestamp 1698175906
transform 1 0 255696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_2277
timestamp 1698175906
transform 1 0 256368 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2341
timestamp 1698175906
transform 1 0 263536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_2347
timestamp 1698175906
transform 1 0 264208 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2411
timestamp 1698175906
transform 1 0 271376 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_2417
timestamp 1698175906
transform 1 0 272048 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2481
timestamp 1698175906
transform 1 0 279216 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_2487
timestamp 1698175906
transform 1 0 279888 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2551
timestamp 1698175906
transform 1 0 287056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_2557
timestamp 1698175906
transform 1 0 287728 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2621
timestamp 1698175906
transform 1 0 294896 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_2627
timestamp 1698175906
transform 1 0 295568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_2643
timestamp 1698175906
transform 1 0 297360 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_2651
timestamp 1698175906
transform 1 0 298256 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698175906
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698175906
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698175906
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698175906
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_492
timestamp 1698175906
transform 1 0 56448 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_556
timestamp 1698175906
transform 1 0 63616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_562
timestamp 1698175906
transform 1 0 64288 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_626
timestamp 1698175906
transform 1 0 71456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_632
timestamp 1698175906
transform 1 0 72128 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_696
timestamp 1698175906
transform 1 0 79296 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_702
timestamp 1698175906
transform 1 0 79968 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_766
timestamp 1698175906
transform 1 0 87136 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_772
timestamp 1698175906
transform 1 0 87808 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_836
timestamp 1698175906
transform 1 0 94976 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_842
timestamp 1698175906
transform 1 0 95648 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_906
timestamp 1698175906
transform 1 0 102816 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_912
timestamp 1698175906
transform 1 0 103488 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_976
timestamp 1698175906
transform 1 0 110656 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_982
timestamp 1698175906
transform 1 0 111328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1046
timestamp 1698175906
transform 1 0 118496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1052
timestamp 1698175906
transform 1 0 119168 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1116
timestamp 1698175906
transform 1 0 126336 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1122
timestamp 1698175906
transform 1 0 127008 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1186
timestamp 1698175906
transform 1 0 134176 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1192
timestamp 1698175906
transform 1 0 134848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1256
timestamp 1698175906
transform 1 0 142016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1262
timestamp 1698175906
transform 1 0 142688 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1326
timestamp 1698175906
transform 1 0 149856 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1332
timestamp 1698175906
transform 1 0 150528 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1396
timestamp 1698175906
transform 1 0 157696 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1402
timestamp 1698175906
transform 1 0 158368 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1466
timestamp 1698175906
transform 1 0 165536 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1472
timestamp 1698175906
transform 1 0 166208 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1536
timestamp 1698175906
transform 1 0 173376 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1542
timestamp 1698175906
transform 1 0 174048 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1606
timestamp 1698175906
transform 1 0 181216 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1612
timestamp 1698175906
transform 1 0 181888 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1676
timestamp 1698175906
transform 1 0 189056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1682
timestamp 1698175906
transform 1 0 189728 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1746
timestamp 1698175906
transform 1 0 196896 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1752
timestamp 1698175906
transform 1 0 197568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1816
timestamp 1698175906
transform 1 0 204736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_1822
timestamp 1698175906
transform 1 0 205408 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_1854
timestamp 1698175906
transform 1 0 208992 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_1870
timestamp 1698175906
transform 1 0 210784 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1878
timestamp 1698175906
transform 1 0 211680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_1882
timestamp 1698175906
transform 1 0 212128 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1892
timestamp 1698175906
transform 1 0 213248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1956
timestamp 1698175906
transform 1 0 220416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1962
timestamp 1698175906
transform 1 0 221088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2026
timestamp 1698175906
transform 1 0 228256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2032
timestamp 1698175906
transform 1 0 228928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2096
timestamp 1698175906
transform 1 0 236096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2102
timestamp 1698175906
transform 1 0 236768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2166
timestamp 1698175906
transform 1 0 243936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2172
timestamp 1698175906
transform 1 0 244608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2236
timestamp 1698175906
transform 1 0 251776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2242
timestamp 1698175906
transform 1 0 252448 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2306
timestamp 1698175906
transform 1 0 259616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2312
timestamp 1698175906
transform 1 0 260288 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2376
timestamp 1698175906
transform 1 0 267456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2382
timestamp 1698175906
transform 1 0 268128 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2446
timestamp 1698175906
transform 1 0 275296 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2452
timestamp 1698175906
transform 1 0 275968 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2516
timestamp 1698175906
transform 1 0 283136 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2522
timestamp 1698175906
transform 1 0 283808 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2586
timestamp 1698175906
transform 1 0 290976 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2592
timestamp 1698175906
transform 1 0 291648 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_2624
timestamp 1698175906
transform 1 0 295232 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_2640
timestamp 1698175906
transform 1 0 297024 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2648
timestamp 1698175906
transform 1 0 297920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698175906
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_387
timestamp 1698175906
transform 1 0 44688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698175906
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_457
timestamp 1698175906
transform 1 0 52528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_521
timestamp 1698175906
transform 1 0 59696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_527
timestamp 1698175906
transform 1 0 60368 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_591
timestamp 1698175906
transform 1 0 67536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_597
timestamp 1698175906
transform 1 0 68208 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_661
timestamp 1698175906
transform 1 0 75376 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_667
timestamp 1698175906
transform 1 0 76048 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_731
timestamp 1698175906
transform 1 0 83216 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_737
timestamp 1698175906
transform 1 0 83888 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_801
timestamp 1698175906
transform 1 0 91056 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_807
timestamp 1698175906
transform 1 0 91728 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_871
timestamp 1698175906
transform 1 0 98896 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_877
timestamp 1698175906
transform 1 0 99568 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_941
timestamp 1698175906
transform 1 0 106736 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_947
timestamp 1698175906
transform 1 0 107408 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1011
timestamp 1698175906
transform 1 0 114576 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1017
timestamp 1698175906
transform 1 0 115248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1081
timestamp 1698175906
transform 1 0 122416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1087
timestamp 1698175906
transform 1 0 123088 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1151
timestamp 1698175906
transform 1 0 130256 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1157
timestamp 1698175906
transform 1 0 130928 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1221
timestamp 1698175906
transform 1 0 138096 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1227
timestamp 1698175906
transform 1 0 138768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1291
timestamp 1698175906
transform 1 0 145936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1297
timestamp 1698175906
transform 1 0 146608 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1361
timestamp 1698175906
transform 1 0 153776 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1367
timestamp 1698175906
transform 1 0 154448 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1431
timestamp 1698175906
transform 1 0 161616 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1437
timestamp 1698175906
transform 1 0 162288 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1501
timestamp 1698175906
transform 1 0 169456 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1507
timestamp 1698175906
transform 1 0 170128 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1571
timestamp 1698175906
transform 1 0 177296 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1577
timestamp 1698175906
transform 1 0 177968 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1641
timestamp 1698175906
transform 1 0 185136 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1647
timestamp 1698175906
transform 1 0 185808 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1711
timestamp 1698175906
transform 1 0 192976 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1717
timestamp 1698175906
transform 1 0 193648 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1781
timestamp 1698175906
transform 1 0 200816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1787
timestamp 1698175906
transform 1 0 201488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1851
timestamp 1698175906
transform 1 0 208656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1857
timestamp 1698175906
transform 1 0 209328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1921
timestamp 1698175906
transform 1 0 216496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1927
timestamp 1698175906
transform 1 0 217168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1991
timestamp 1698175906
transform 1 0 224336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1997
timestamp 1698175906
transform 1 0 225008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2061
timestamp 1698175906
transform 1 0 232176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_2067
timestamp 1698175906
transform 1 0 232848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2131
timestamp 1698175906
transform 1 0 240016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_2137
timestamp 1698175906
transform 1 0 240688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2201
timestamp 1698175906
transform 1 0 247856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_2207
timestamp 1698175906
transform 1 0 248528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2271
timestamp 1698175906
transform 1 0 255696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_2277
timestamp 1698175906
transform 1 0 256368 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2341
timestamp 1698175906
transform 1 0 263536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_2347
timestamp 1698175906
transform 1 0 264208 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2411
timestamp 1698175906
transform 1 0 271376 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_2417
timestamp 1698175906
transform 1 0 272048 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2481
timestamp 1698175906
transform 1 0 279216 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_2487
timestamp 1698175906
transform 1 0 279888 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2551
timestamp 1698175906
transform 1 0 287056 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_2557
timestamp 1698175906
transform 1 0 287728 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2621
timestamp 1698175906
transform 1 0 294896 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2627
timestamp 1698175906
transform 1 0 295568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_2643
timestamp 1698175906
transform 1 0 297360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_2651
timestamp 1698175906
transform 1 0 298256 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698175906
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698175906
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698175906
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698175906
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_492
timestamp 1698175906
transform 1 0 56448 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_556
timestamp 1698175906
transform 1 0 63616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_562
timestamp 1698175906
transform 1 0 64288 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_626
timestamp 1698175906
transform 1 0 71456 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_632
timestamp 1698175906
transform 1 0 72128 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_696
timestamp 1698175906
transform 1 0 79296 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_702
timestamp 1698175906
transform 1 0 79968 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_766
timestamp 1698175906
transform 1 0 87136 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_772
timestamp 1698175906
transform 1 0 87808 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_836
timestamp 1698175906
transform 1 0 94976 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_842
timestamp 1698175906
transform 1 0 95648 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_906
timestamp 1698175906
transform 1 0 102816 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_912
timestamp 1698175906
transform 1 0 103488 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_976
timestamp 1698175906
transform 1 0 110656 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_982
timestamp 1698175906
transform 1 0 111328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1046
timestamp 1698175906
transform 1 0 118496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1052
timestamp 1698175906
transform 1 0 119168 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1116
timestamp 1698175906
transform 1 0 126336 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1122
timestamp 1698175906
transform 1 0 127008 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1186
timestamp 1698175906
transform 1 0 134176 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1192
timestamp 1698175906
transform 1 0 134848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1256
timestamp 1698175906
transform 1 0 142016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1262
timestamp 1698175906
transform 1 0 142688 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1326
timestamp 1698175906
transform 1 0 149856 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1332
timestamp 1698175906
transform 1 0 150528 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1396
timestamp 1698175906
transform 1 0 157696 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1402
timestamp 1698175906
transform 1 0 158368 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1466
timestamp 1698175906
transform 1 0 165536 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1472
timestamp 1698175906
transform 1 0 166208 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1536
timestamp 1698175906
transform 1 0 173376 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1542
timestamp 1698175906
transform 1 0 174048 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1606
timestamp 1698175906
transform 1 0 181216 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1612
timestamp 1698175906
transform 1 0 181888 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1676
timestamp 1698175906
transform 1 0 189056 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1682
timestamp 1698175906
transform 1 0 189728 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1746
timestamp 1698175906
transform 1 0 196896 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1752
timestamp 1698175906
transform 1 0 197568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1816
timestamp 1698175906
transform 1 0 204736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1822
timestamp 1698175906
transform 1 0 205408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1886
timestamp 1698175906
transform 1 0 212576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1892
timestamp 1698175906
transform 1 0 213248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1956
timestamp 1698175906
transform 1 0 220416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1962
timestamp 1698175906
transform 1 0 221088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2026
timestamp 1698175906
transform 1 0 228256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2032
timestamp 1698175906
transform 1 0 228928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2096
timestamp 1698175906
transform 1 0 236096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2102
timestamp 1698175906
transform 1 0 236768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2166
timestamp 1698175906
transform 1 0 243936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2172
timestamp 1698175906
transform 1 0 244608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2236
timestamp 1698175906
transform 1 0 251776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2242
timestamp 1698175906
transform 1 0 252448 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2306
timestamp 1698175906
transform 1 0 259616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2312
timestamp 1698175906
transform 1 0 260288 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2376
timestamp 1698175906
transform 1 0 267456 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2382
timestamp 1698175906
transform 1 0 268128 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2446
timestamp 1698175906
transform 1 0 275296 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2452
timestamp 1698175906
transform 1 0 275968 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2516
timestamp 1698175906
transform 1 0 283136 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2522
timestamp 1698175906
transform 1 0 283808 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2586
timestamp 1698175906
transform 1 0 290976 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_2592
timestamp 1698175906
transform 1 0 291648 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2624
timestamp 1698175906
transform 1 0 295232 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_2640
timestamp 1698175906
transform 1 0 297024 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2648
timestamp 1698175906
transform 1 0 297920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698175906
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698175906
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698175906
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_457
timestamp 1698175906
transform 1 0 52528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_521
timestamp 1698175906
transform 1 0 59696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_527
timestamp 1698175906
transform 1 0 60368 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_591
timestamp 1698175906
transform 1 0 67536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_597
timestamp 1698175906
transform 1 0 68208 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_661
timestamp 1698175906
transform 1 0 75376 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_667
timestamp 1698175906
transform 1 0 76048 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_731
timestamp 1698175906
transform 1 0 83216 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_737
timestamp 1698175906
transform 1 0 83888 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_801
timestamp 1698175906
transform 1 0 91056 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_807
timestamp 1698175906
transform 1 0 91728 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_871
timestamp 1698175906
transform 1 0 98896 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_877
timestamp 1698175906
transform 1 0 99568 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_941
timestamp 1698175906
transform 1 0 106736 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_947
timestamp 1698175906
transform 1 0 107408 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1011
timestamp 1698175906
transform 1 0 114576 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1017
timestamp 1698175906
transform 1 0 115248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1081
timestamp 1698175906
transform 1 0 122416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1087
timestamp 1698175906
transform 1 0 123088 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1151
timestamp 1698175906
transform 1 0 130256 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1157
timestamp 1698175906
transform 1 0 130928 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1221
timestamp 1698175906
transform 1 0 138096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1227
timestamp 1698175906
transform 1 0 138768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1291
timestamp 1698175906
transform 1 0 145936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1297
timestamp 1698175906
transform 1 0 146608 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1361
timestamp 1698175906
transform 1 0 153776 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1367
timestamp 1698175906
transform 1 0 154448 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1431
timestamp 1698175906
transform 1 0 161616 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1437
timestamp 1698175906
transform 1 0 162288 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1501
timestamp 1698175906
transform 1 0 169456 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1507
timestamp 1698175906
transform 1 0 170128 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1571
timestamp 1698175906
transform 1 0 177296 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1577
timestamp 1698175906
transform 1 0 177968 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1641
timestamp 1698175906
transform 1 0 185136 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1647
timestamp 1698175906
transform 1 0 185808 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1711
timestamp 1698175906
transform 1 0 192976 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1717
timestamp 1698175906
transform 1 0 193648 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1781
timestamp 1698175906
transform 1 0 200816 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1787
timestamp 1698175906
transform 1 0 201488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1851
timestamp 1698175906
transform 1 0 208656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1857
timestamp 1698175906
transform 1 0 209328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1921
timestamp 1698175906
transform 1 0 216496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1927
timestamp 1698175906
transform 1 0 217168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1991
timestamp 1698175906
transform 1 0 224336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1997
timestamp 1698175906
transform 1 0 225008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2061
timestamp 1698175906
transform 1 0 232176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_2067
timestamp 1698175906
transform 1 0 232848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2131
timestamp 1698175906
transform 1 0 240016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_2137
timestamp 1698175906
transform 1 0 240688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2201
timestamp 1698175906
transform 1 0 247856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_2207
timestamp 1698175906
transform 1 0 248528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2271
timestamp 1698175906
transform 1 0 255696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_2277
timestamp 1698175906
transform 1 0 256368 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2341
timestamp 1698175906
transform 1 0 263536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_2347
timestamp 1698175906
transform 1 0 264208 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2411
timestamp 1698175906
transform 1 0 271376 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_2417
timestamp 1698175906
transform 1 0 272048 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2481
timestamp 1698175906
transform 1 0 279216 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_2487
timestamp 1698175906
transform 1 0 279888 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2551
timestamp 1698175906
transform 1 0 287056 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_2557
timestamp 1698175906
transform 1 0 287728 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2621
timestamp 1698175906
transform 1 0 294896 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2627
timestamp 1698175906
transform 1 0 295568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_2643
timestamp 1698175906
transform 1 0 297360 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_2651
timestamp 1698175906
transform 1 0 298256 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698175906
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698175906
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698175906
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698175906
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_492
timestamp 1698175906
transform 1 0 56448 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_556
timestamp 1698175906
transform 1 0 63616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_562
timestamp 1698175906
transform 1 0 64288 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_626
timestamp 1698175906
transform 1 0 71456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_632
timestamp 1698175906
transform 1 0 72128 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_696
timestamp 1698175906
transform 1 0 79296 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_702
timestamp 1698175906
transform 1 0 79968 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_766
timestamp 1698175906
transform 1 0 87136 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_772
timestamp 1698175906
transform 1 0 87808 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_836
timestamp 1698175906
transform 1 0 94976 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_842
timestamp 1698175906
transform 1 0 95648 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_906
timestamp 1698175906
transform 1 0 102816 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_912
timestamp 1698175906
transform 1 0 103488 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_976
timestamp 1698175906
transform 1 0 110656 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_982
timestamp 1698175906
transform 1 0 111328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1046
timestamp 1698175906
transform 1 0 118496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1052
timestamp 1698175906
transform 1 0 119168 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1116
timestamp 1698175906
transform 1 0 126336 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1122
timestamp 1698175906
transform 1 0 127008 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1186
timestamp 1698175906
transform 1 0 134176 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1192
timestamp 1698175906
transform 1 0 134848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1256
timestamp 1698175906
transform 1 0 142016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1262
timestamp 1698175906
transform 1 0 142688 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1326
timestamp 1698175906
transform 1 0 149856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1332
timestamp 1698175906
transform 1 0 150528 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1396
timestamp 1698175906
transform 1 0 157696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1402
timestamp 1698175906
transform 1 0 158368 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1466
timestamp 1698175906
transform 1 0 165536 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1472
timestamp 1698175906
transform 1 0 166208 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1536
timestamp 1698175906
transform 1 0 173376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1542
timestamp 1698175906
transform 1 0 174048 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1606
timestamp 1698175906
transform 1 0 181216 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1612
timestamp 1698175906
transform 1 0 181888 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1676
timestamp 1698175906
transform 1 0 189056 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1682
timestamp 1698175906
transform 1 0 189728 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1746
timestamp 1698175906
transform 1 0 196896 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1752
timestamp 1698175906
transform 1 0 197568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1816
timestamp 1698175906
transform 1 0 204736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1822
timestamp 1698175906
transform 1 0 205408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1886
timestamp 1698175906
transform 1 0 212576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1892
timestamp 1698175906
transform 1 0 213248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1956
timestamp 1698175906
transform 1 0 220416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1962
timestamp 1698175906
transform 1 0 221088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2026
timestamp 1698175906
transform 1 0 228256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2032
timestamp 1698175906
transform 1 0 228928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2096
timestamp 1698175906
transform 1 0 236096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2102
timestamp 1698175906
transform 1 0 236768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2166
timestamp 1698175906
transform 1 0 243936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2172
timestamp 1698175906
transform 1 0 244608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2236
timestamp 1698175906
transform 1 0 251776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2242
timestamp 1698175906
transform 1 0 252448 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2306
timestamp 1698175906
transform 1 0 259616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2312
timestamp 1698175906
transform 1 0 260288 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2376
timestamp 1698175906
transform 1 0 267456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2382
timestamp 1698175906
transform 1 0 268128 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2446
timestamp 1698175906
transform 1 0 275296 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2452
timestamp 1698175906
transform 1 0 275968 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2516
timestamp 1698175906
transform 1 0 283136 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2522
timestamp 1698175906
transform 1 0 283808 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2586
timestamp 1698175906
transform 1 0 290976 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2592
timestamp 1698175906
transform 1 0 291648 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_2624
timestamp 1698175906
transform 1 0 295232 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_2640
timestamp 1698175906
transform 1 0 297024 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2648
timestamp 1698175906
transform 1 0 297920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698175906
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698175906
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698175906
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_457
timestamp 1698175906
transform 1 0 52528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_521
timestamp 1698175906
transform 1 0 59696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_527
timestamp 1698175906
transform 1 0 60368 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_591
timestamp 1698175906
transform 1 0 67536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_597
timestamp 1698175906
transform 1 0 68208 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_661
timestamp 1698175906
transform 1 0 75376 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_667
timestamp 1698175906
transform 1 0 76048 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_731
timestamp 1698175906
transform 1 0 83216 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_737
timestamp 1698175906
transform 1 0 83888 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_801
timestamp 1698175906
transform 1 0 91056 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_807
timestamp 1698175906
transform 1 0 91728 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_871
timestamp 1698175906
transform 1 0 98896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_877
timestamp 1698175906
transform 1 0 99568 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_941
timestamp 1698175906
transform 1 0 106736 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_947
timestamp 1698175906
transform 1 0 107408 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1011
timestamp 1698175906
transform 1 0 114576 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1017
timestamp 1698175906
transform 1 0 115248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1081
timestamp 1698175906
transform 1 0 122416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1087
timestamp 1698175906
transform 1 0 123088 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1151
timestamp 1698175906
transform 1 0 130256 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1157
timestamp 1698175906
transform 1 0 130928 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1221
timestamp 1698175906
transform 1 0 138096 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1227
timestamp 1698175906
transform 1 0 138768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1291
timestamp 1698175906
transform 1 0 145936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1297
timestamp 1698175906
transform 1 0 146608 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1361
timestamp 1698175906
transform 1 0 153776 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1367
timestamp 1698175906
transform 1 0 154448 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1431
timestamp 1698175906
transform 1 0 161616 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1437
timestamp 1698175906
transform 1 0 162288 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1501
timestamp 1698175906
transform 1 0 169456 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1507
timestamp 1698175906
transform 1 0 170128 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1571
timestamp 1698175906
transform 1 0 177296 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1577
timestamp 1698175906
transform 1 0 177968 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1641
timestamp 1698175906
transform 1 0 185136 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1647
timestamp 1698175906
transform 1 0 185808 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1711
timestamp 1698175906
transform 1 0 192976 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1717
timestamp 1698175906
transform 1 0 193648 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1781
timestamp 1698175906
transform 1 0 200816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1787
timestamp 1698175906
transform 1 0 201488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1851
timestamp 1698175906
transform 1 0 208656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1857
timestamp 1698175906
transform 1 0 209328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1921
timestamp 1698175906
transform 1 0 216496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1927
timestamp 1698175906
transform 1 0 217168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1991
timestamp 1698175906
transform 1 0 224336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1997
timestamp 1698175906
transform 1 0 225008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2061
timestamp 1698175906
transform 1 0 232176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_2067
timestamp 1698175906
transform 1 0 232848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2131
timestamp 1698175906
transform 1 0 240016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_2137
timestamp 1698175906
transform 1 0 240688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2201
timestamp 1698175906
transform 1 0 247856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_2207
timestamp 1698175906
transform 1 0 248528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2271
timestamp 1698175906
transform 1 0 255696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_2277
timestamp 1698175906
transform 1 0 256368 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2341
timestamp 1698175906
transform 1 0 263536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_2347
timestamp 1698175906
transform 1 0 264208 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2411
timestamp 1698175906
transform 1 0 271376 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_2417
timestamp 1698175906
transform 1 0 272048 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2481
timestamp 1698175906
transform 1 0 279216 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_2487
timestamp 1698175906
transform 1 0 279888 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2551
timestamp 1698175906
transform 1 0 287056 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_2557
timestamp 1698175906
transform 1 0 287728 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2621
timestamp 1698175906
transform 1 0 294896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2627
timestamp 1698175906
transform 1 0 295568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_2643
timestamp 1698175906
transform 1 0 297360 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_2651
timestamp 1698175906
transform 1 0 298256 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698175906
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698175906
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698175906
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698175906
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_492
timestamp 1698175906
transform 1 0 56448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_556
timestamp 1698175906
transform 1 0 63616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_562
timestamp 1698175906
transform 1 0 64288 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_626
timestamp 1698175906
transform 1 0 71456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_632
timestamp 1698175906
transform 1 0 72128 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_696
timestamp 1698175906
transform 1 0 79296 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_702
timestamp 1698175906
transform 1 0 79968 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_766
timestamp 1698175906
transform 1 0 87136 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_772
timestamp 1698175906
transform 1 0 87808 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_836
timestamp 1698175906
transform 1 0 94976 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_842
timestamp 1698175906
transform 1 0 95648 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_906
timestamp 1698175906
transform 1 0 102816 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_912
timestamp 1698175906
transform 1 0 103488 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_976
timestamp 1698175906
transform 1 0 110656 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_982
timestamp 1698175906
transform 1 0 111328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1046
timestamp 1698175906
transform 1 0 118496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1052
timestamp 1698175906
transform 1 0 119168 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1116
timestamp 1698175906
transform 1 0 126336 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1122
timestamp 1698175906
transform 1 0 127008 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1186
timestamp 1698175906
transform 1 0 134176 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1192
timestamp 1698175906
transform 1 0 134848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1256
timestamp 1698175906
transform 1 0 142016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1262
timestamp 1698175906
transform 1 0 142688 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1326
timestamp 1698175906
transform 1 0 149856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1332
timestamp 1698175906
transform 1 0 150528 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1396
timestamp 1698175906
transform 1 0 157696 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1402
timestamp 1698175906
transform 1 0 158368 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1466
timestamp 1698175906
transform 1 0 165536 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1472
timestamp 1698175906
transform 1 0 166208 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1536
timestamp 1698175906
transform 1 0 173376 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1542
timestamp 1698175906
transform 1 0 174048 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1606
timestamp 1698175906
transform 1 0 181216 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1612
timestamp 1698175906
transform 1 0 181888 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1676
timestamp 1698175906
transform 1 0 189056 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1682
timestamp 1698175906
transform 1 0 189728 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1746
timestamp 1698175906
transform 1 0 196896 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1752
timestamp 1698175906
transform 1 0 197568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1816
timestamp 1698175906
transform 1 0 204736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1822
timestamp 1698175906
transform 1 0 205408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1886
timestamp 1698175906
transform 1 0 212576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1892
timestamp 1698175906
transform 1 0 213248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1956
timestamp 1698175906
transform 1 0 220416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1962
timestamp 1698175906
transform 1 0 221088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2026
timestamp 1698175906
transform 1 0 228256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2032
timestamp 1698175906
transform 1 0 228928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2096
timestamp 1698175906
transform 1 0 236096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2102
timestamp 1698175906
transform 1 0 236768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2166
timestamp 1698175906
transform 1 0 243936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2172
timestamp 1698175906
transform 1 0 244608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2236
timestamp 1698175906
transform 1 0 251776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2242
timestamp 1698175906
transform 1 0 252448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2306
timestamp 1698175906
transform 1 0 259616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2312
timestamp 1698175906
transform 1 0 260288 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2376
timestamp 1698175906
transform 1 0 267456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2382
timestamp 1698175906
transform 1 0 268128 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2446
timestamp 1698175906
transform 1 0 275296 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2452
timestamp 1698175906
transform 1 0 275968 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2516
timestamp 1698175906
transform 1 0 283136 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2522
timestamp 1698175906
transform 1 0 283808 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2586
timestamp 1698175906
transform 1 0 290976 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_2592
timestamp 1698175906
transform 1 0 291648 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_2624
timestamp 1698175906
transform 1 0 295232 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_2640
timestamp 1698175906
transform 1 0 297024 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2648
timestamp 1698175906
transform 1 0 297920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698175906
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698175906
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698175906
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_457
timestamp 1698175906
transform 1 0 52528 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_521
timestamp 1698175906
transform 1 0 59696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_527
timestamp 1698175906
transform 1 0 60368 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_591
timestamp 1698175906
transform 1 0 67536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_597
timestamp 1698175906
transform 1 0 68208 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_661
timestamp 1698175906
transform 1 0 75376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_667
timestamp 1698175906
transform 1 0 76048 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_731
timestamp 1698175906
transform 1 0 83216 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_737
timestamp 1698175906
transform 1 0 83888 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_801
timestamp 1698175906
transform 1 0 91056 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_807
timestamp 1698175906
transform 1 0 91728 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_871
timestamp 1698175906
transform 1 0 98896 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_877
timestamp 1698175906
transform 1 0 99568 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_941
timestamp 1698175906
transform 1 0 106736 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_947
timestamp 1698175906
transform 1 0 107408 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1011
timestamp 1698175906
transform 1 0 114576 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1017
timestamp 1698175906
transform 1 0 115248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1081
timestamp 1698175906
transform 1 0 122416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1087
timestamp 1698175906
transform 1 0 123088 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1151
timestamp 1698175906
transform 1 0 130256 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1157
timestamp 1698175906
transform 1 0 130928 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1221
timestamp 1698175906
transform 1 0 138096 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1227
timestamp 1698175906
transform 1 0 138768 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1291
timestamp 1698175906
transform 1 0 145936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1297
timestamp 1698175906
transform 1 0 146608 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1361
timestamp 1698175906
transform 1 0 153776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1367
timestamp 1698175906
transform 1 0 154448 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1431
timestamp 1698175906
transform 1 0 161616 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1437
timestamp 1698175906
transform 1 0 162288 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1501
timestamp 1698175906
transform 1 0 169456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1507
timestamp 1698175906
transform 1 0 170128 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1571
timestamp 1698175906
transform 1 0 177296 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1577
timestamp 1698175906
transform 1 0 177968 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1641
timestamp 1698175906
transform 1 0 185136 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1647
timestamp 1698175906
transform 1 0 185808 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1711
timestamp 1698175906
transform 1 0 192976 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1717
timestamp 1698175906
transform 1 0 193648 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1781
timestamp 1698175906
transform 1 0 200816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1787
timestamp 1698175906
transform 1 0 201488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1851
timestamp 1698175906
transform 1 0 208656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1857
timestamp 1698175906
transform 1 0 209328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1921
timestamp 1698175906
transform 1 0 216496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1927
timestamp 1698175906
transform 1 0 217168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1991
timestamp 1698175906
transform 1 0 224336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1997
timestamp 1698175906
transform 1 0 225008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2061
timestamp 1698175906
transform 1 0 232176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_2067
timestamp 1698175906
transform 1 0 232848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2131
timestamp 1698175906
transform 1 0 240016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_2137
timestamp 1698175906
transform 1 0 240688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2201
timestamp 1698175906
transform 1 0 247856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_2207
timestamp 1698175906
transform 1 0 248528 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2271
timestamp 1698175906
transform 1 0 255696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_2277
timestamp 1698175906
transform 1 0 256368 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2341
timestamp 1698175906
transform 1 0 263536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_2347
timestamp 1698175906
transform 1 0 264208 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2411
timestamp 1698175906
transform 1 0 271376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_2417
timestamp 1698175906
transform 1 0 272048 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2481
timestamp 1698175906
transform 1 0 279216 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_2487
timestamp 1698175906
transform 1 0 279888 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2551
timestamp 1698175906
transform 1 0 287056 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_2557
timestamp 1698175906
transform 1 0 287728 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2621
timestamp 1698175906
transform 1 0 294896 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2627
timestamp 1698175906
transform 1 0 295568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_2643
timestamp 1698175906
transform 1 0 297360 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_2651
timestamp 1698175906
transform 1 0 298256 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698175906
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698175906
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698175906
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698175906
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_492
timestamp 1698175906
transform 1 0 56448 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_556
timestamp 1698175906
transform 1 0 63616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_562
timestamp 1698175906
transform 1 0 64288 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_626
timestamp 1698175906
transform 1 0 71456 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_632
timestamp 1698175906
transform 1 0 72128 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_696
timestamp 1698175906
transform 1 0 79296 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_702
timestamp 1698175906
transform 1 0 79968 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_766
timestamp 1698175906
transform 1 0 87136 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_772
timestamp 1698175906
transform 1 0 87808 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_836
timestamp 1698175906
transform 1 0 94976 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_842
timestamp 1698175906
transform 1 0 95648 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_906
timestamp 1698175906
transform 1 0 102816 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_912
timestamp 1698175906
transform 1 0 103488 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_976
timestamp 1698175906
transform 1 0 110656 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_982
timestamp 1698175906
transform 1 0 111328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1046
timestamp 1698175906
transform 1 0 118496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1052
timestamp 1698175906
transform 1 0 119168 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1116
timestamp 1698175906
transform 1 0 126336 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1122
timestamp 1698175906
transform 1 0 127008 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1186
timestamp 1698175906
transform 1 0 134176 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1192
timestamp 1698175906
transform 1 0 134848 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1256
timestamp 1698175906
transform 1 0 142016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1262
timestamp 1698175906
transform 1 0 142688 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1326
timestamp 1698175906
transform 1 0 149856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1332
timestamp 1698175906
transform 1 0 150528 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1396
timestamp 1698175906
transform 1 0 157696 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1402
timestamp 1698175906
transform 1 0 158368 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1466
timestamp 1698175906
transform 1 0 165536 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1472
timestamp 1698175906
transform 1 0 166208 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1536
timestamp 1698175906
transform 1 0 173376 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1542
timestamp 1698175906
transform 1 0 174048 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1606
timestamp 1698175906
transform 1 0 181216 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1612
timestamp 1698175906
transform 1 0 181888 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1676
timestamp 1698175906
transform 1 0 189056 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1682
timestamp 1698175906
transform 1 0 189728 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1746
timestamp 1698175906
transform 1 0 196896 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1752
timestamp 1698175906
transform 1 0 197568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1816
timestamp 1698175906
transform 1 0 204736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1822
timestamp 1698175906
transform 1 0 205408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1886
timestamp 1698175906
transform 1 0 212576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1892
timestamp 1698175906
transform 1 0 213248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1956
timestamp 1698175906
transform 1 0 220416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1962
timestamp 1698175906
transform 1 0 221088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2026
timestamp 1698175906
transform 1 0 228256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2032
timestamp 1698175906
transform 1 0 228928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2096
timestamp 1698175906
transform 1 0 236096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2102
timestamp 1698175906
transform 1 0 236768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2166
timestamp 1698175906
transform 1 0 243936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2172
timestamp 1698175906
transform 1 0 244608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2236
timestamp 1698175906
transform 1 0 251776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2242
timestamp 1698175906
transform 1 0 252448 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2306
timestamp 1698175906
transform 1 0 259616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2312
timestamp 1698175906
transform 1 0 260288 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2376
timestamp 1698175906
transform 1 0 267456 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2382
timestamp 1698175906
transform 1 0 268128 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2446
timestamp 1698175906
transform 1 0 275296 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2452
timestamp 1698175906
transform 1 0 275968 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2516
timestamp 1698175906
transform 1 0 283136 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2522
timestamp 1698175906
transform 1 0 283808 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2586
timestamp 1698175906
transform 1 0 290976 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_2592
timestamp 1698175906
transform 1 0 291648 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_2624
timestamp 1698175906
transform 1 0 295232 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2640
timestamp 1698175906
transform 1 0 297024 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2648
timestamp 1698175906
transform 1 0 297920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698175906
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698175906
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698175906
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_457
timestamp 1698175906
transform 1 0 52528 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_521
timestamp 1698175906
transform 1 0 59696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_527
timestamp 1698175906
transform 1 0 60368 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_591
timestamp 1698175906
transform 1 0 67536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_597
timestamp 1698175906
transform 1 0 68208 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_661
timestamp 1698175906
transform 1 0 75376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_667
timestamp 1698175906
transform 1 0 76048 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_731
timestamp 1698175906
transform 1 0 83216 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_737
timestamp 1698175906
transform 1 0 83888 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_801
timestamp 1698175906
transform 1 0 91056 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_807
timestamp 1698175906
transform 1 0 91728 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_871
timestamp 1698175906
transform 1 0 98896 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_877
timestamp 1698175906
transform 1 0 99568 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_941
timestamp 1698175906
transform 1 0 106736 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_947
timestamp 1698175906
transform 1 0 107408 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1011
timestamp 1698175906
transform 1 0 114576 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1017
timestamp 1698175906
transform 1 0 115248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1081
timestamp 1698175906
transform 1 0 122416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1087
timestamp 1698175906
transform 1 0 123088 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1151
timestamp 1698175906
transform 1 0 130256 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1157
timestamp 1698175906
transform 1 0 130928 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1221
timestamp 1698175906
transform 1 0 138096 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1227
timestamp 1698175906
transform 1 0 138768 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1291
timestamp 1698175906
transform 1 0 145936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1297
timestamp 1698175906
transform 1 0 146608 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1361
timestamp 1698175906
transform 1 0 153776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1367
timestamp 1698175906
transform 1 0 154448 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1431
timestamp 1698175906
transform 1 0 161616 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1437
timestamp 1698175906
transform 1 0 162288 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1501
timestamp 1698175906
transform 1 0 169456 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1507
timestamp 1698175906
transform 1 0 170128 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1571
timestamp 1698175906
transform 1 0 177296 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1577
timestamp 1698175906
transform 1 0 177968 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1641
timestamp 1698175906
transform 1 0 185136 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1647
timestamp 1698175906
transform 1 0 185808 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1711
timestamp 1698175906
transform 1 0 192976 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1717
timestamp 1698175906
transform 1 0 193648 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1781
timestamp 1698175906
transform 1 0 200816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1787
timestamp 1698175906
transform 1 0 201488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1851
timestamp 1698175906
transform 1 0 208656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1857
timestamp 1698175906
transform 1 0 209328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1921
timestamp 1698175906
transform 1 0 216496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1927
timestamp 1698175906
transform 1 0 217168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1991
timestamp 1698175906
transform 1 0 224336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1997
timestamp 1698175906
transform 1 0 225008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2061
timestamp 1698175906
transform 1 0 232176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_2067
timestamp 1698175906
transform 1 0 232848 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2131
timestamp 1698175906
transform 1 0 240016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_2137
timestamp 1698175906
transform 1 0 240688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2201
timestamp 1698175906
transform 1 0 247856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_2207
timestamp 1698175906
transform 1 0 248528 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2271
timestamp 1698175906
transform 1 0 255696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_2277
timestamp 1698175906
transform 1 0 256368 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2341
timestamp 1698175906
transform 1 0 263536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_2347
timestamp 1698175906
transform 1 0 264208 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2411
timestamp 1698175906
transform 1 0 271376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_2417
timestamp 1698175906
transform 1 0 272048 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2481
timestamp 1698175906
transform 1 0 279216 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_2487
timestamp 1698175906
transform 1 0 279888 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2551
timestamp 1698175906
transform 1 0 287056 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_2557
timestamp 1698175906
transform 1 0 287728 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2621
timestamp 1698175906
transform 1 0 294896 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_2627
timestamp 1698175906
transform 1 0 295568 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_2643
timestamp 1698175906
transform 1 0 297360 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_2651
timestamp 1698175906
transform 1 0 298256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698175906
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698175906
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698175906
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698175906
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_492
timestamp 1698175906
transform 1 0 56448 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_556
timestamp 1698175906
transform 1 0 63616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_562
timestamp 1698175906
transform 1 0 64288 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_626
timestamp 1698175906
transform 1 0 71456 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_632
timestamp 1698175906
transform 1 0 72128 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_696
timestamp 1698175906
transform 1 0 79296 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_702
timestamp 1698175906
transform 1 0 79968 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_766
timestamp 1698175906
transform 1 0 87136 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_772
timestamp 1698175906
transform 1 0 87808 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_836
timestamp 1698175906
transform 1 0 94976 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_842
timestamp 1698175906
transform 1 0 95648 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_906
timestamp 1698175906
transform 1 0 102816 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_912
timestamp 1698175906
transform 1 0 103488 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_976
timestamp 1698175906
transform 1 0 110656 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_982
timestamp 1698175906
transform 1 0 111328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1046
timestamp 1698175906
transform 1 0 118496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1052
timestamp 1698175906
transform 1 0 119168 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1116
timestamp 1698175906
transform 1 0 126336 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1122
timestamp 1698175906
transform 1 0 127008 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1186
timestamp 1698175906
transform 1 0 134176 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1192
timestamp 1698175906
transform 1 0 134848 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1256
timestamp 1698175906
transform 1 0 142016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1262
timestamp 1698175906
transform 1 0 142688 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1326
timestamp 1698175906
transform 1 0 149856 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1332
timestamp 1698175906
transform 1 0 150528 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1396
timestamp 1698175906
transform 1 0 157696 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1402
timestamp 1698175906
transform 1 0 158368 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1466
timestamp 1698175906
transform 1 0 165536 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1472
timestamp 1698175906
transform 1 0 166208 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1536
timestamp 1698175906
transform 1 0 173376 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1542
timestamp 1698175906
transform 1 0 174048 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1606
timestamp 1698175906
transform 1 0 181216 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1612
timestamp 1698175906
transform 1 0 181888 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1676
timestamp 1698175906
transform 1 0 189056 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1682
timestamp 1698175906
transform 1 0 189728 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1746
timestamp 1698175906
transform 1 0 196896 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1752
timestamp 1698175906
transform 1 0 197568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1816
timestamp 1698175906
transform 1 0 204736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1822
timestamp 1698175906
transform 1 0 205408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1886
timestamp 1698175906
transform 1 0 212576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1892
timestamp 1698175906
transform 1 0 213248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1956
timestamp 1698175906
transform 1 0 220416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1962
timestamp 1698175906
transform 1 0 221088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2026
timestamp 1698175906
transform 1 0 228256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2032
timestamp 1698175906
transform 1 0 228928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2096
timestamp 1698175906
transform 1 0 236096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2102
timestamp 1698175906
transform 1 0 236768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2166
timestamp 1698175906
transform 1 0 243936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2172
timestamp 1698175906
transform 1 0 244608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2236
timestamp 1698175906
transform 1 0 251776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2242
timestamp 1698175906
transform 1 0 252448 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2306
timestamp 1698175906
transform 1 0 259616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2312
timestamp 1698175906
transform 1 0 260288 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2376
timestamp 1698175906
transform 1 0 267456 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2382
timestamp 1698175906
transform 1 0 268128 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2446
timestamp 1698175906
transform 1 0 275296 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2452
timestamp 1698175906
transform 1 0 275968 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2516
timestamp 1698175906
transform 1 0 283136 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2522
timestamp 1698175906
transform 1 0 283808 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2586
timestamp 1698175906
transform 1 0 290976 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_2592
timestamp 1698175906
transform 1 0 291648 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_2624
timestamp 1698175906
transform 1 0 295232 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_2640
timestamp 1698175906
transform 1 0 297024 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2648
timestamp 1698175906
transform 1 0 297920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698175906
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_381
timestamp 1698175906
transform 1 0 44016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698175906
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698175906
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_457
timestamp 1698175906
transform 1 0 52528 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_521
timestamp 1698175906
transform 1 0 59696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_527
timestamp 1698175906
transform 1 0 60368 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_591
timestamp 1698175906
transform 1 0 67536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_597
timestamp 1698175906
transform 1 0 68208 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_661
timestamp 1698175906
transform 1 0 75376 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_667
timestamp 1698175906
transform 1 0 76048 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_731
timestamp 1698175906
transform 1 0 83216 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_737
timestamp 1698175906
transform 1 0 83888 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_801
timestamp 1698175906
transform 1 0 91056 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_807
timestamp 1698175906
transform 1 0 91728 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_871
timestamp 1698175906
transform 1 0 98896 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_877
timestamp 1698175906
transform 1 0 99568 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_941
timestamp 1698175906
transform 1 0 106736 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_947
timestamp 1698175906
transform 1 0 107408 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1011
timestamp 1698175906
transform 1 0 114576 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1017
timestamp 1698175906
transform 1 0 115248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1081
timestamp 1698175906
transform 1 0 122416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1087
timestamp 1698175906
transform 1 0 123088 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1151
timestamp 1698175906
transform 1 0 130256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1157
timestamp 1698175906
transform 1 0 130928 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1221
timestamp 1698175906
transform 1 0 138096 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1227
timestamp 1698175906
transform 1 0 138768 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1291
timestamp 1698175906
transform 1 0 145936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1297
timestamp 1698175906
transform 1 0 146608 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1361
timestamp 1698175906
transform 1 0 153776 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1367
timestamp 1698175906
transform 1 0 154448 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1431
timestamp 1698175906
transform 1 0 161616 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1437
timestamp 1698175906
transform 1 0 162288 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1501
timestamp 1698175906
transform 1 0 169456 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1507
timestamp 1698175906
transform 1 0 170128 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1571
timestamp 1698175906
transform 1 0 177296 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1577
timestamp 1698175906
transform 1 0 177968 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1641
timestamp 1698175906
transform 1 0 185136 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1647
timestamp 1698175906
transform 1 0 185808 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1711
timestamp 1698175906
transform 1 0 192976 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1717
timestamp 1698175906
transform 1 0 193648 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1781
timestamp 1698175906
transform 1 0 200816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1787
timestamp 1698175906
transform 1 0 201488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1851
timestamp 1698175906
transform 1 0 208656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1857
timestamp 1698175906
transform 1 0 209328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1921
timestamp 1698175906
transform 1 0 216496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1927
timestamp 1698175906
transform 1 0 217168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1991
timestamp 1698175906
transform 1 0 224336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1997
timestamp 1698175906
transform 1 0 225008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2061
timestamp 1698175906
transform 1 0 232176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_2067
timestamp 1698175906
transform 1 0 232848 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2131
timestamp 1698175906
transform 1 0 240016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_2137
timestamp 1698175906
transform 1 0 240688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2201
timestamp 1698175906
transform 1 0 247856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_2207
timestamp 1698175906
transform 1 0 248528 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2271
timestamp 1698175906
transform 1 0 255696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_2277
timestamp 1698175906
transform 1 0 256368 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2341
timestamp 1698175906
transform 1 0 263536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_2347
timestamp 1698175906
transform 1 0 264208 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2411
timestamp 1698175906
transform 1 0 271376 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_2417
timestamp 1698175906
transform 1 0 272048 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2481
timestamp 1698175906
transform 1 0 279216 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_2487
timestamp 1698175906
transform 1 0 279888 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2551
timestamp 1698175906
transform 1 0 287056 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_2557
timestamp 1698175906
transform 1 0 287728 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2621
timestamp 1698175906
transform 1 0 294896 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_2627
timestamp 1698175906
transform 1 0 295568 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_2643
timestamp 1698175906
transform 1 0 297360 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_2651
timestamp 1698175906
transform 1 0 298256 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698175906
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_352
timestamp 1698175906
transform 1 0 40768 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698175906
transform 1 0 47936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698175906
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698175906
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_492
timestamp 1698175906
transform 1 0 56448 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_556
timestamp 1698175906
transform 1 0 63616 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_562
timestamp 1698175906
transform 1 0 64288 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_626
timestamp 1698175906
transform 1 0 71456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_632
timestamp 1698175906
transform 1 0 72128 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_696
timestamp 1698175906
transform 1 0 79296 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_702
timestamp 1698175906
transform 1 0 79968 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_766
timestamp 1698175906
transform 1 0 87136 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_772
timestamp 1698175906
transform 1 0 87808 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_836
timestamp 1698175906
transform 1 0 94976 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_842
timestamp 1698175906
transform 1 0 95648 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_906
timestamp 1698175906
transform 1 0 102816 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_912
timestamp 1698175906
transform 1 0 103488 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_976
timestamp 1698175906
transform 1 0 110656 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_982
timestamp 1698175906
transform 1 0 111328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1046
timestamp 1698175906
transform 1 0 118496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1052
timestamp 1698175906
transform 1 0 119168 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1116
timestamp 1698175906
transform 1 0 126336 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1122
timestamp 1698175906
transform 1 0 127008 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1186
timestamp 1698175906
transform 1 0 134176 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1192
timestamp 1698175906
transform 1 0 134848 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1256
timestamp 1698175906
transform 1 0 142016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1262
timestamp 1698175906
transform 1 0 142688 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1326
timestamp 1698175906
transform 1 0 149856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1332
timestamp 1698175906
transform 1 0 150528 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1396
timestamp 1698175906
transform 1 0 157696 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1402
timestamp 1698175906
transform 1 0 158368 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1466
timestamp 1698175906
transform 1 0 165536 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1472
timestamp 1698175906
transform 1 0 166208 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1536
timestamp 1698175906
transform 1 0 173376 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1542
timestamp 1698175906
transform 1 0 174048 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1606
timestamp 1698175906
transform 1 0 181216 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1612
timestamp 1698175906
transform 1 0 181888 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1676
timestamp 1698175906
transform 1 0 189056 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1682
timestamp 1698175906
transform 1 0 189728 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1746
timestamp 1698175906
transform 1 0 196896 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1752
timestamp 1698175906
transform 1 0 197568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1816
timestamp 1698175906
transform 1 0 204736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1822
timestamp 1698175906
transform 1 0 205408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1886
timestamp 1698175906
transform 1 0 212576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1892
timestamp 1698175906
transform 1 0 213248 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1956
timestamp 1698175906
transform 1 0 220416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1962
timestamp 1698175906
transform 1 0 221088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2026
timestamp 1698175906
transform 1 0 228256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2032
timestamp 1698175906
transform 1 0 228928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2096
timestamp 1698175906
transform 1 0 236096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2102
timestamp 1698175906
transform 1 0 236768 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2166
timestamp 1698175906
transform 1 0 243936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2172
timestamp 1698175906
transform 1 0 244608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2236
timestamp 1698175906
transform 1 0 251776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2242
timestamp 1698175906
transform 1 0 252448 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2306
timestamp 1698175906
transform 1 0 259616 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2312
timestamp 1698175906
transform 1 0 260288 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2376
timestamp 1698175906
transform 1 0 267456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2382
timestamp 1698175906
transform 1 0 268128 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2446
timestamp 1698175906
transform 1 0 275296 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2452
timestamp 1698175906
transform 1 0 275968 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2516
timestamp 1698175906
transform 1 0 283136 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2522
timestamp 1698175906
transform 1 0 283808 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2586
timestamp 1698175906
transform 1 0 290976 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_2592
timestamp 1698175906
transform 1 0 291648 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_2624
timestamp 1698175906
transform 1 0 295232 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_2640
timestamp 1698175906
transform 1 0 297024 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2648
timestamp 1698175906
transform 1 0 297920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698175906
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_381
timestamp 1698175906
transform 1 0 44016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_387
timestamp 1698175906
transform 1 0 44688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698175906
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_457
timestamp 1698175906
transform 1 0 52528 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_521
timestamp 1698175906
transform 1 0 59696 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_527
timestamp 1698175906
transform 1 0 60368 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_591
timestamp 1698175906
transform 1 0 67536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_597
timestamp 1698175906
transform 1 0 68208 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_661
timestamp 1698175906
transform 1 0 75376 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_667
timestamp 1698175906
transform 1 0 76048 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_731
timestamp 1698175906
transform 1 0 83216 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_737
timestamp 1698175906
transform 1 0 83888 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_801
timestamp 1698175906
transform 1 0 91056 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_807
timestamp 1698175906
transform 1 0 91728 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_871
timestamp 1698175906
transform 1 0 98896 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_877
timestamp 1698175906
transform 1 0 99568 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_941
timestamp 1698175906
transform 1 0 106736 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_947
timestamp 1698175906
transform 1 0 107408 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1011
timestamp 1698175906
transform 1 0 114576 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1017
timestamp 1698175906
transform 1 0 115248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1081
timestamp 1698175906
transform 1 0 122416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1087
timestamp 1698175906
transform 1 0 123088 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1151
timestamp 1698175906
transform 1 0 130256 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1157
timestamp 1698175906
transform 1 0 130928 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1221
timestamp 1698175906
transform 1 0 138096 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1227
timestamp 1698175906
transform 1 0 138768 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1291
timestamp 1698175906
transform 1 0 145936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1297
timestamp 1698175906
transform 1 0 146608 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1361
timestamp 1698175906
transform 1 0 153776 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1367
timestamp 1698175906
transform 1 0 154448 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1431
timestamp 1698175906
transform 1 0 161616 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1437
timestamp 1698175906
transform 1 0 162288 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1501
timestamp 1698175906
transform 1 0 169456 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1507
timestamp 1698175906
transform 1 0 170128 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1571
timestamp 1698175906
transform 1 0 177296 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1577
timestamp 1698175906
transform 1 0 177968 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1641
timestamp 1698175906
transform 1 0 185136 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1647
timestamp 1698175906
transform 1 0 185808 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1711
timestamp 1698175906
transform 1 0 192976 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1717
timestamp 1698175906
transform 1 0 193648 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1781
timestamp 1698175906
transform 1 0 200816 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1787
timestamp 1698175906
transform 1 0 201488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1851
timestamp 1698175906
transform 1 0 208656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1857
timestamp 1698175906
transform 1 0 209328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1921
timestamp 1698175906
transform 1 0 216496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1927
timestamp 1698175906
transform 1 0 217168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1991
timestamp 1698175906
transform 1 0 224336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1997
timestamp 1698175906
transform 1 0 225008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2061
timestamp 1698175906
transform 1 0 232176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_2067
timestamp 1698175906
transform 1 0 232848 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2131
timestamp 1698175906
transform 1 0 240016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_2137
timestamp 1698175906
transform 1 0 240688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2201
timestamp 1698175906
transform 1 0 247856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_2207
timestamp 1698175906
transform 1 0 248528 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2271
timestamp 1698175906
transform 1 0 255696 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_2277
timestamp 1698175906
transform 1 0 256368 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2341
timestamp 1698175906
transform 1 0 263536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_2347
timestamp 1698175906
transform 1 0 264208 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2411
timestamp 1698175906
transform 1 0 271376 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_2417
timestamp 1698175906
transform 1 0 272048 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2481
timestamp 1698175906
transform 1 0 279216 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_2487
timestamp 1698175906
transform 1 0 279888 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2551
timestamp 1698175906
transform 1 0 287056 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_2557
timestamp 1698175906
transform 1 0 287728 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2621
timestamp 1698175906
transform 1 0 294896 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_2627
timestamp 1698175906
transform 1 0 295568 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_2643
timestamp 1698175906
transform 1 0 297360 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_2651
timestamp 1698175906
transform 1 0 298256 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_346
timestamp 1698175906
transform 1 0 40096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_352
timestamp 1698175906
transform 1 0 40768 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698175906
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_422
timestamp 1698175906
transform 1 0 48608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698175906
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_492
timestamp 1698175906
transform 1 0 56448 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_556
timestamp 1698175906
transform 1 0 63616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_562
timestamp 1698175906
transform 1 0 64288 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_626
timestamp 1698175906
transform 1 0 71456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_632
timestamp 1698175906
transform 1 0 72128 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_696
timestamp 1698175906
transform 1 0 79296 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_702
timestamp 1698175906
transform 1 0 79968 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_766
timestamp 1698175906
transform 1 0 87136 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_772
timestamp 1698175906
transform 1 0 87808 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_836
timestamp 1698175906
transform 1 0 94976 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_842
timestamp 1698175906
transform 1 0 95648 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_906
timestamp 1698175906
transform 1 0 102816 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_912
timestamp 1698175906
transform 1 0 103488 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_976
timestamp 1698175906
transform 1 0 110656 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_982
timestamp 1698175906
transform 1 0 111328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1046
timestamp 1698175906
transform 1 0 118496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1052
timestamp 1698175906
transform 1 0 119168 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1116
timestamp 1698175906
transform 1 0 126336 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1122
timestamp 1698175906
transform 1 0 127008 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1186
timestamp 1698175906
transform 1 0 134176 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1192
timestamp 1698175906
transform 1 0 134848 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1256
timestamp 1698175906
transform 1 0 142016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1262
timestamp 1698175906
transform 1 0 142688 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1326
timestamp 1698175906
transform 1 0 149856 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1332
timestamp 1698175906
transform 1 0 150528 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1396
timestamp 1698175906
transform 1 0 157696 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1402
timestamp 1698175906
transform 1 0 158368 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1466
timestamp 1698175906
transform 1 0 165536 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1472
timestamp 1698175906
transform 1 0 166208 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1536
timestamp 1698175906
transform 1 0 173376 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1542
timestamp 1698175906
transform 1 0 174048 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1606
timestamp 1698175906
transform 1 0 181216 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1612
timestamp 1698175906
transform 1 0 181888 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1676
timestamp 1698175906
transform 1 0 189056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1682
timestamp 1698175906
transform 1 0 189728 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1746
timestamp 1698175906
transform 1 0 196896 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1752
timestamp 1698175906
transform 1 0 197568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1816
timestamp 1698175906
transform 1 0 204736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1822
timestamp 1698175906
transform 1 0 205408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1886
timestamp 1698175906
transform 1 0 212576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1892
timestamp 1698175906
transform 1 0 213248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1956
timestamp 1698175906
transform 1 0 220416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1962
timestamp 1698175906
transform 1 0 221088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2026
timestamp 1698175906
transform 1 0 228256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2032
timestamp 1698175906
transform 1 0 228928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2096
timestamp 1698175906
transform 1 0 236096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2102
timestamp 1698175906
transform 1 0 236768 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2166
timestamp 1698175906
transform 1 0 243936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2172
timestamp 1698175906
transform 1 0 244608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2236
timestamp 1698175906
transform 1 0 251776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2242
timestamp 1698175906
transform 1 0 252448 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2306
timestamp 1698175906
transform 1 0 259616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2312
timestamp 1698175906
transform 1 0 260288 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2376
timestamp 1698175906
transform 1 0 267456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2382
timestamp 1698175906
transform 1 0 268128 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2446
timestamp 1698175906
transform 1 0 275296 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2452
timestamp 1698175906
transform 1 0 275968 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2516
timestamp 1698175906
transform 1 0 283136 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2522
timestamp 1698175906
transform 1 0 283808 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2586
timestamp 1698175906
transform 1 0 290976 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_2592
timestamp 1698175906
transform 1 0 291648 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_2624
timestamp 1698175906
transform 1 0 295232 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2640
timestamp 1698175906
transform 1 0 297024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2648
timestamp 1698175906
transform 1 0 297920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698175906
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698175906
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_381
timestamp 1698175906
transform 1 0 44016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_387
timestamp 1698175906
transform 1 0 44688 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_451
timestamp 1698175906
transform 1 0 51856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_457
timestamp 1698175906
transform 1 0 52528 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_521
timestamp 1698175906
transform 1 0 59696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_527
timestamp 1698175906
transform 1 0 60368 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_591
timestamp 1698175906
transform 1 0 67536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_597
timestamp 1698175906
transform 1 0 68208 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_661
timestamp 1698175906
transform 1 0 75376 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_667
timestamp 1698175906
transform 1 0 76048 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_731
timestamp 1698175906
transform 1 0 83216 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_737
timestamp 1698175906
transform 1 0 83888 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_801
timestamp 1698175906
transform 1 0 91056 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_807
timestamp 1698175906
transform 1 0 91728 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_871
timestamp 1698175906
transform 1 0 98896 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_877
timestamp 1698175906
transform 1 0 99568 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_941
timestamp 1698175906
transform 1 0 106736 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_947
timestamp 1698175906
transform 1 0 107408 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1011
timestamp 1698175906
transform 1 0 114576 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1017
timestamp 1698175906
transform 1 0 115248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1081
timestamp 1698175906
transform 1 0 122416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1087
timestamp 1698175906
transform 1 0 123088 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1151
timestamp 1698175906
transform 1 0 130256 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1157
timestamp 1698175906
transform 1 0 130928 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1221
timestamp 1698175906
transform 1 0 138096 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1227
timestamp 1698175906
transform 1 0 138768 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1291
timestamp 1698175906
transform 1 0 145936 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1297
timestamp 1698175906
transform 1 0 146608 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1361
timestamp 1698175906
transform 1 0 153776 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1367
timestamp 1698175906
transform 1 0 154448 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1431
timestamp 1698175906
transform 1 0 161616 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1437
timestamp 1698175906
transform 1 0 162288 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1501
timestamp 1698175906
transform 1 0 169456 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1507
timestamp 1698175906
transform 1 0 170128 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1571
timestamp 1698175906
transform 1 0 177296 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1577
timestamp 1698175906
transform 1 0 177968 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1641
timestamp 1698175906
transform 1 0 185136 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1647
timestamp 1698175906
transform 1 0 185808 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1711
timestamp 1698175906
transform 1 0 192976 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1717
timestamp 1698175906
transform 1 0 193648 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1781
timestamp 1698175906
transform 1 0 200816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1787
timestamp 1698175906
transform 1 0 201488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1851
timestamp 1698175906
transform 1 0 208656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1857
timestamp 1698175906
transform 1 0 209328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1921
timestamp 1698175906
transform 1 0 216496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1927
timestamp 1698175906
transform 1 0 217168 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1991
timestamp 1698175906
transform 1 0 224336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1997
timestamp 1698175906
transform 1 0 225008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2061
timestamp 1698175906
transform 1 0 232176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_2067
timestamp 1698175906
transform 1 0 232848 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2131
timestamp 1698175906
transform 1 0 240016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_2137
timestamp 1698175906
transform 1 0 240688 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2201
timestamp 1698175906
transform 1 0 247856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_2207
timestamp 1698175906
transform 1 0 248528 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2271
timestamp 1698175906
transform 1 0 255696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_2277
timestamp 1698175906
transform 1 0 256368 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2341
timestamp 1698175906
transform 1 0 263536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_2347
timestamp 1698175906
transform 1 0 264208 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2411
timestamp 1698175906
transform 1 0 271376 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_2417
timestamp 1698175906
transform 1 0 272048 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2481
timestamp 1698175906
transform 1 0 279216 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_2487
timestamp 1698175906
transform 1 0 279888 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2551
timestamp 1698175906
transform 1 0 287056 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_2557
timestamp 1698175906
transform 1 0 287728 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2621
timestamp 1698175906
transform 1 0 294896 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_2627
timestamp 1698175906
transform 1 0 295568 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_2643
timestamp 1698175906
transform 1 0 297360 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_2651
timestamp 1698175906
transform 1 0 298256 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698175906
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_352
timestamp 1698175906
transform 1 0 40768 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698175906
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_422
timestamp 1698175906
transform 1 0 48608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698175906
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_492
timestamp 1698175906
transform 1 0 56448 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_556
timestamp 1698175906
transform 1 0 63616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_562
timestamp 1698175906
transform 1 0 64288 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_626
timestamp 1698175906
transform 1 0 71456 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_632
timestamp 1698175906
transform 1 0 72128 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_696
timestamp 1698175906
transform 1 0 79296 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_702
timestamp 1698175906
transform 1 0 79968 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_766
timestamp 1698175906
transform 1 0 87136 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_772
timestamp 1698175906
transform 1 0 87808 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_836
timestamp 1698175906
transform 1 0 94976 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_842
timestamp 1698175906
transform 1 0 95648 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_906
timestamp 1698175906
transform 1 0 102816 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_912
timestamp 1698175906
transform 1 0 103488 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_976
timestamp 1698175906
transform 1 0 110656 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_982
timestamp 1698175906
transform 1 0 111328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1046
timestamp 1698175906
transform 1 0 118496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1052
timestamp 1698175906
transform 1 0 119168 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1116
timestamp 1698175906
transform 1 0 126336 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1122
timestamp 1698175906
transform 1 0 127008 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1186
timestamp 1698175906
transform 1 0 134176 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1192
timestamp 1698175906
transform 1 0 134848 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1256
timestamp 1698175906
transform 1 0 142016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1262
timestamp 1698175906
transform 1 0 142688 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1326
timestamp 1698175906
transform 1 0 149856 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1332
timestamp 1698175906
transform 1 0 150528 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1396
timestamp 1698175906
transform 1 0 157696 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1402
timestamp 1698175906
transform 1 0 158368 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1466
timestamp 1698175906
transform 1 0 165536 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1472
timestamp 1698175906
transform 1 0 166208 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1536
timestamp 1698175906
transform 1 0 173376 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1542
timestamp 1698175906
transform 1 0 174048 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1606
timestamp 1698175906
transform 1 0 181216 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1612
timestamp 1698175906
transform 1 0 181888 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1676
timestamp 1698175906
transform 1 0 189056 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1682
timestamp 1698175906
transform 1 0 189728 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1746
timestamp 1698175906
transform 1 0 196896 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1752
timestamp 1698175906
transform 1 0 197568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1816
timestamp 1698175906
transform 1 0 204736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1822
timestamp 1698175906
transform 1 0 205408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1886
timestamp 1698175906
transform 1 0 212576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1892
timestamp 1698175906
transform 1 0 213248 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1956
timestamp 1698175906
transform 1 0 220416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1962
timestamp 1698175906
transform 1 0 221088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2026
timestamp 1698175906
transform 1 0 228256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2032
timestamp 1698175906
transform 1 0 228928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2096
timestamp 1698175906
transform 1 0 236096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2102
timestamp 1698175906
transform 1 0 236768 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2166
timestamp 1698175906
transform 1 0 243936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2172
timestamp 1698175906
transform 1 0 244608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2236
timestamp 1698175906
transform 1 0 251776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2242
timestamp 1698175906
transform 1 0 252448 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2306
timestamp 1698175906
transform 1 0 259616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2312
timestamp 1698175906
transform 1 0 260288 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2376
timestamp 1698175906
transform 1 0 267456 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2382
timestamp 1698175906
transform 1 0 268128 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2446
timestamp 1698175906
transform 1 0 275296 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2452
timestamp 1698175906
transform 1 0 275968 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2516
timestamp 1698175906
transform 1 0 283136 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2522
timestamp 1698175906
transform 1 0 283808 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2586
timestamp 1698175906
transform 1 0 290976 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_2592
timestamp 1698175906
transform 1 0 291648 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2624
timestamp 1698175906
transform 1 0 295232 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_2640
timestamp 1698175906
transform 1 0 297024 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2648
timestamp 1698175906
transform 1 0 297920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_381
timestamp 1698175906
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_387
timestamp 1698175906
transform 1 0 44688 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_451
timestamp 1698175906
transform 1 0 51856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_457
timestamp 1698175906
transform 1 0 52528 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_521
timestamp 1698175906
transform 1 0 59696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_527
timestamp 1698175906
transform 1 0 60368 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_591
timestamp 1698175906
transform 1 0 67536 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_597
timestamp 1698175906
transform 1 0 68208 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_661
timestamp 1698175906
transform 1 0 75376 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_667
timestamp 1698175906
transform 1 0 76048 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_731
timestamp 1698175906
transform 1 0 83216 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_737
timestamp 1698175906
transform 1 0 83888 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_801
timestamp 1698175906
transform 1 0 91056 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_807
timestamp 1698175906
transform 1 0 91728 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_871
timestamp 1698175906
transform 1 0 98896 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_877
timestamp 1698175906
transform 1 0 99568 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_941
timestamp 1698175906
transform 1 0 106736 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_947
timestamp 1698175906
transform 1 0 107408 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1011
timestamp 1698175906
transform 1 0 114576 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1017
timestamp 1698175906
transform 1 0 115248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1081
timestamp 1698175906
transform 1 0 122416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1087
timestamp 1698175906
transform 1 0 123088 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1151
timestamp 1698175906
transform 1 0 130256 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1157
timestamp 1698175906
transform 1 0 130928 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1221
timestamp 1698175906
transform 1 0 138096 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1227
timestamp 1698175906
transform 1 0 138768 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1291
timestamp 1698175906
transform 1 0 145936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1297
timestamp 1698175906
transform 1 0 146608 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1361
timestamp 1698175906
transform 1 0 153776 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1367
timestamp 1698175906
transform 1 0 154448 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1431
timestamp 1698175906
transform 1 0 161616 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1437
timestamp 1698175906
transform 1 0 162288 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1501
timestamp 1698175906
transform 1 0 169456 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1507
timestamp 1698175906
transform 1 0 170128 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1571
timestamp 1698175906
transform 1 0 177296 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1577
timestamp 1698175906
transform 1 0 177968 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1641
timestamp 1698175906
transform 1 0 185136 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1647
timestamp 1698175906
transform 1 0 185808 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1711
timestamp 1698175906
transform 1 0 192976 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1717
timestamp 1698175906
transform 1 0 193648 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1781
timestamp 1698175906
transform 1 0 200816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1787
timestamp 1698175906
transform 1 0 201488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1851
timestamp 1698175906
transform 1 0 208656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1857
timestamp 1698175906
transform 1 0 209328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1921
timestamp 1698175906
transform 1 0 216496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1927
timestamp 1698175906
transform 1 0 217168 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1991
timestamp 1698175906
transform 1 0 224336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1997
timestamp 1698175906
transform 1 0 225008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2061
timestamp 1698175906
transform 1 0 232176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_2067
timestamp 1698175906
transform 1 0 232848 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2131
timestamp 1698175906
transform 1 0 240016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_2137
timestamp 1698175906
transform 1 0 240688 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2201
timestamp 1698175906
transform 1 0 247856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_2207
timestamp 1698175906
transform 1 0 248528 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2271
timestamp 1698175906
transform 1 0 255696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_2277
timestamp 1698175906
transform 1 0 256368 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2341
timestamp 1698175906
transform 1 0 263536 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_2347
timestamp 1698175906
transform 1 0 264208 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2411
timestamp 1698175906
transform 1 0 271376 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_2417
timestamp 1698175906
transform 1 0 272048 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2481
timestamp 1698175906
transform 1 0 279216 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_2487
timestamp 1698175906
transform 1 0 279888 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2551
timestamp 1698175906
transform 1 0 287056 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_2557
timestamp 1698175906
transform 1 0 287728 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2621
timestamp 1698175906
transform 1 0 294896 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_2627
timestamp 1698175906
transform 1 0 295568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_2643
timestamp 1698175906
transform 1 0 297360 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_2651
timestamp 1698175906
transform 1 0 298256 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_352
timestamp 1698175906
transform 1 0 40768 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698175906
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698175906
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698175906
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_492
timestamp 1698175906
transform 1 0 56448 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_556
timestamp 1698175906
transform 1 0 63616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_562
timestamp 1698175906
transform 1 0 64288 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_626
timestamp 1698175906
transform 1 0 71456 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_632
timestamp 1698175906
transform 1 0 72128 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_696
timestamp 1698175906
transform 1 0 79296 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_702
timestamp 1698175906
transform 1 0 79968 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_766
timestamp 1698175906
transform 1 0 87136 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_772
timestamp 1698175906
transform 1 0 87808 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_836
timestamp 1698175906
transform 1 0 94976 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_842
timestamp 1698175906
transform 1 0 95648 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_906
timestamp 1698175906
transform 1 0 102816 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_912
timestamp 1698175906
transform 1 0 103488 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_976
timestamp 1698175906
transform 1 0 110656 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_982
timestamp 1698175906
transform 1 0 111328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1046
timestamp 1698175906
transform 1 0 118496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1052
timestamp 1698175906
transform 1 0 119168 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1116
timestamp 1698175906
transform 1 0 126336 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1122
timestamp 1698175906
transform 1 0 127008 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1186
timestamp 1698175906
transform 1 0 134176 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1192
timestamp 1698175906
transform 1 0 134848 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1256
timestamp 1698175906
transform 1 0 142016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1262
timestamp 1698175906
transform 1 0 142688 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1326
timestamp 1698175906
transform 1 0 149856 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1332
timestamp 1698175906
transform 1 0 150528 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1396
timestamp 1698175906
transform 1 0 157696 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1402
timestamp 1698175906
transform 1 0 158368 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1466
timestamp 1698175906
transform 1 0 165536 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1472
timestamp 1698175906
transform 1 0 166208 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1536
timestamp 1698175906
transform 1 0 173376 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1542
timestamp 1698175906
transform 1 0 174048 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1606
timestamp 1698175906
transform 1 0 181216 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1612
timestamp 1698175906
transform 1 0 181888 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1676
timestamp 1698175906
transform 1 0 189056 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1682
timestamp 1698175906
transform 1 0 189728 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1746
timestamp 1698175906
transform 1 0 196896 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1752
timestamp 1698175906
transform 1 0 197568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1816
timestamp 1698175906
transform 1 0 204736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1822
timestamp 1698175906
transform 1 0 205408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1886
timestamp 1698175906
transform 1 0 212576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1892
timestamp 1698175906
transform 1 0 213248 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1956
timestamp 1698175906
transform 1 0 220416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1962
timestamp 1698175906
transform 1 0 221088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2026
timestamp 1698175906
transform 1 0 228256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2032
timestamp 1698175906
transform 1 0 228928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2096
timestamp 1698175906
transform 1 0 236096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2102
timestamp 1698175906
transform 1 0 236768 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2166
timestamp 1698175906
transform 1 0 243936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2172
timestamp 1698175906
transform 1 0 244608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2236
timestamp 1698175906
transform 1 0 251776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2242
timestamp 1698175906
transform 1 0 252448 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2306
timestamp 1698175906
transform 1 0 259616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2312
timestamp 1698175906
transform 1 0 260288 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2376
timestamp 1698175906
transform 1 0 267456 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2382
timestamp 1698175906
transform 1 0 268128 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2446
timestamp 1698175906
transform 1 0 275296 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2452
timestamp 1698175906
transform 1 0 275968 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2516
timestamp 1698175906
transform 1 0 283136 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2522
timestamp 1698175906
transform 1 0 283808 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2586
timestamp 1698175906
transform 1 0 290976 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_2592
timestamp 1698175906
transform 1 0 291648 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_2624
timestamp 1698175906
transform 1 0 295232 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_2640
timestamp 1698175906
transform 1 0 297024 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2648
timestamp 1698175906
transform 1 0 297920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698175906
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_381
timestamp 1698175906
transform 1 0 44016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_387
timestamp 1698175906
transform 1 0 44688 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698175906
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_457
timestamp 1698175906
transform 1 0 52528 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_521
timestamp 1698175906
transform 1 0 59696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_527
timestamp 1698175906
transform 1 0 60368 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_591
timestamp 1698175906
transform 1 0 67536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_597
timestamp 1698175906
transform 1 0 68208 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_661
timestamp 1698175906
transform 1 0 75376 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_667
timestamp 1698175906
transform 1 0 76048 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_731
timestamp 1698175906
transform 1 0 83216 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_737
timestamp 1698175906
transform 1 0 83888 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_801
timestamp 1698175906
transform 1 0 91056 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_807
timestamp 1698175906
transform 1 0 91728 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_871
timestamp 1698175906
transform 1 0 98896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_877
timestamp 1698175906
transform 1 0 99568 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_941
timestamp 1698175906
transform 1 0 106736 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_947
timestamp 1698175906
transform 1 0 107408 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1011
timestamp 1698175906
transform 1 0 114576 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1017
timestamp 1698175906
transform 1 0 115248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1081
timestamp 1698175906
transform 1 0 122416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1087
timestamp 1698175906
transform 1 0 123088 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1151
timestamp 1698175906
transform 1 0 130256 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1157
timestamp 1698175906
transform 1 0 130928 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1221
timestamp 1698175906
transform 1 0 138096 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1227
timestamp 1698175906
transform 1 0 138768 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1291
timestamp 1698175906
transform 1 0 145936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1297
timestamp 1698175906
transform 1 0 146608 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1361
timestamp 1698175906
transform 1 0 153776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1367
timestamp 1698175906
transform 1 0 154448 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1431
timestamp 1698175906
transform 1 0 161616 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1437
timestamp 1698175906
transform 1 0 162288 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1501
timestamp 1698175906
transform 1 0 169456 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1507
timestamp 1698175906
transform 1 0 170128 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1571
timestamp 1698175906
transform 1 0 177296 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1577
timestamp 1698175906
transform 1 0 177968 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1641
timestamp 1698175906
transform 1 0 185136 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1647
timestamp 1698175906
transform 1 0 185808 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1711
timestamp 1698175906
transform 1 0 192976 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1717
timestamp 1698175906
transform 1 0 193648 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1781
timestamp 1698175906
transform 1 0 200816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1787
timestamp 1698175906
transform 1 0 201488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1851
timestamp 1698175906
transform 1 0 208656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1857
timestamp 1698175906
transform 1 0 209328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1921
timestamp 1698175906
transform 1 0 216496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1927
timestamp 1698175906
transform 1 0 217168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1991
timestamp 1698175906
transform 1 0 224336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1997
timestamp 1698175906
transform 1 0 225008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2061
timestamp 1698175906
transform 1 0 232176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_2067
timestamp 1698175906
transform 1 0 232848 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2131
timestamp 1698175906
transform 1 0 240016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_2137
timestamp 1698175906
transform 1 0 240688 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2201
timestamp 1698175906
transform 1 0 247856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_2207
timestamp 1698175906
transform 1 0 248528 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2271
timestamp 1698175906
transform 1 0 255696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_2277
timestamp 1698175906
transform 1 0 256368 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2341
timestamp 1698175906
transform 1 0 263536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_2347
timestamp 1698175906
transform 1 0 264208 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2411
timestamp 1698175906
transform 1 0 271376 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_2417
timestamp 1698175906
transform 1 0 272048 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2481
timestamp 1698175906
transform 1 0 279216 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_2487
timestamp 1698175906
transform 1 0 279888 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2551
timestamp 1698175906
transform 1 0 287056 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_2557
timestamp 1698175906
transform 1 0 287728 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2621
timestamp 1698175906
transform 1 0 294896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_2627
timestamp 1698175906
transform 1 0 295568 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_2643
timestamp 1698175906
transform 1 0 297360 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_2651
timestamp 1698175906
transform 1 0 298256 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698175906
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_352
timestamp 1698175906
transform 1 0 40768 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_416
timestamp 1698175906
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_422
timestamp 1698175906
transform 1 0 48608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698175906
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_492
timestamp 1698175906
transform 1 0 56448 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_556
timestamp 1698175906
transform 1 0 63616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_562
timestamp 1698175906
transform 1 0 64288 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_626
timestamp 1698175906
transform 1 0 71456 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_632
timestamp 1698175906
transform 1 0 72128 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_696
timestamp 1698175906
transform 1 0 79296 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_702
timestamp 1698175906
transform 1 0 79968 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_766
timestamp 1698175906
transform 1 0 87136 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_772
timestamp 1698175906
transform 1 0 87808 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_836
timestamp 1698175906
transform 1 0 94976 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_842
timestamp 1698175906
transform 1 0 95648 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_906
timestamp 1698175906
transform 1 0 102816 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_912
timestamp 1698175906
transform 1 0 103488 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_976
timestamp 1698175906
transform 1 0 110656 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_982
timestamp 1698175906
transform 1 0 111328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1046
timestamp 1698175906
transform 1 0 118496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1052
timestamp 1698175906
transform 1 0 119168 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1116
timestamp 1698175906
transform 1 0 126336 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1122
timestamp 1698175906
transform 1 0 127008 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1186
timestamp 1698175906
transform 1 0 134176 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1192
timestamp 1698175906
transform 1 0 134848 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1256
timestamp 1698175906
transform 1 0 142016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1262
timestamp 1698175906
transform 1 0 142688 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1326
timestamp 1698175906
transform 1 0 149856 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1332
timestamp 1698175906
transform 1 0 150528 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1396
timestamp 1698175906
transform 1 0 157696 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1402
timestamp 1698175906
transform 1 0 158368 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1466
timestamp 1698175906
transform 1 0 165536 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1472
timestamp 1698175906
transform 1 0 166208 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1536
timestamp 1698175906
transform 1 0 173376 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1542
timestamp 1698175906
transform 1 0 174048 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1606
timestamp 1698175906
transform 1 0 181216 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1612
timestamp 1698175906
transform 1 0 181888 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1676
timestamp 1698175906
transform 1 0 189056 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1682
timestamp 1698175906
transform 1 0 189728 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1746
timestamp 1698175906
transform 1 0 196896 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1752
timestamp 1698175906
transform 1 0 197568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1816
timestamp 1698175906
transform 1 0 204736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1822
timestamp 1698175906
transform 1 0 205408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1886
timestamp 1698175906
transform 1 0 212576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1892
timestamp 1698175906
transform 1 0 213248 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1956
timestamp 1698175906
transform 1 0 220416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1962
timestamp 1698175906
transform 1 0 221088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2026
timestamp 1698175906
transform 1 0 228256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2032
timestamp 1698175906
transform 1 0 228928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2096
timestamp 1698175906
transform 1 0 236096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2102
timestamp 1698175906
transform 1 0 236768 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2166
timestamp 1698175906
transform 1 0 243936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2172
timestamp 1698175906
transform 1 0 244608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2236
timestamp 1698175906
transform 1 0 251776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2242
timestamp 1698175906
transform 1 0 252448 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2306
timestamp 1698175906
transform 1 0 259616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2312
timestamp 1698175906
transform 1 0 260288 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2376
timestamp 1698175906
transform 1 0 267456 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2382
timestamp 1698175906
transform 1 0 268128 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2446
timestamp 1698175906
transform 1 0 275296 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2452
timestamp 1698175906
transform 1 0 275968 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2516
timestamp 1698175906
transform 1 0 283136 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2522
timestamp 1698175906
transform 1 0 283808 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2586
timestamp 1698175906
transform 1 0 290976 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2592
timestamp 1698175906
transform 1 0 291648 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2624
timestamp 1698175906
transform 1 0 295232 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_2640
timestamp 1698175906
transform 1 0 297024 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2648
timestamp 1698175906
transform 1 0 297920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_381
timestamp 1698175906
transform 1 0 44016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698175906
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698175906
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_457
timestamp 1698175906
transform 1 0 52528 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_521
timestamp 1698175906
transform 1 0 59696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_527
timestamp 1698175906
transform 1 0 60368 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_591
timestamp 1698175906
transform 1 0 67536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_597
timestamp 1698175906
transform 1 0 68208 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_661
timestamp 1698175906
transform 1 0 75376 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_667
timestamp 1698175906
transform 1 0 76048 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_731
timestamp 1698175906
transform 1 0 83216 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_737
timestamp 1698175906
transform 1 0 83888 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_801
timestamp 1698175906
transform 1 0 91056 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_807
timestamp 1698175906
transform 1 0 91728 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_871
timestamp 1698175906
transform 1 0 98896 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_877
timestamp 1698175906
transform 1 0 99568 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_941
timestamp 1698175906
transform 1 0 106736 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_947
timestamp 1698175906
transform 1 0 107408 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1011
timestamp 1698175906
transform 1 0 114576 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1017
timestamp 1698175906
transform 1 0 115248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1081
timestamp 1698175906
transform 1 0 122416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1087
timestamp 1698175906
transform 1 0 123088 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1151
timestamp 1698175906
transform 1 0 130256 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1157
timestamp 1698175906
transform 1 0 130928 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1221
timestamp 1698175906
transform 1 0 138096 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1227
timestamp 1698175906
transform 1 0 138768 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1291
timestamp 1698175906
transform 1 0 145936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1297
timestamp 1698175906
transform 1 0 146608 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1361
timestamp 1698175906
transform 1 0 153776 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1367
timestamp 1698175906
transform 1 0 154448 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1431
timestamp 1698175906
transform 1 0 161616 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1437
timestamp 1698175906
transform 1 0 162288 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1501
timestamp 1698175906
transform 1 0 169456 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1507
timestamp 1698175906
transform 1 0 170128 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1571
timestamp 1698175906
transform 1 0 177296 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1577
timestamp 1698175906
transform 1 0 177968 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1641
timestamp 1698175906
transform 1 0 185136 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1647
timestamp 1698175906
transform 1 0 185808 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1711
timestamp 1698175906
transform 1 0 192976 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1717
timestamp 1698175906
transform 1 0 193648 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1781
timestamp 1698175906
transform 1 0 200816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1787
timestamp 1698175906
transform 1 0 201488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1851
timestamp 1698175906
transform 1 0 208656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1857
timestamp 1698175906
transform 1 0 209328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1921
timestamp 1698175906
transform 1 0 216496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1927
timestamp 1698175906
transform 1 0 217168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1991
timestamp 1698175906
transform 1 0 224336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1997
timestamp 1698175906
transform 1 0 225008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2061
timestamp 1698175906
transform 1 0 232176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_2067
timestamp 1698175906
transform 1 0 232848 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2131
timestamp 1698175906
transform 1 0 240016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_2137
timestamp 1698175906
transform 1 0 240688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2201
timestamp 1698175906
transform 1 0 247856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_2207
timestamp 1698175906
transform 1 0 248528 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2271
timestamp 1698175906
transform 1 0 255696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_2277
timestamp 1698175906
transform 1 0 256368 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2341
timestamp 1698175906
transform 1 0 263536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_2347
timestamp 1698175906
transform 1 0 264208 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2411
timestamp 1698175906
transform 1 0 271376 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_2417
timestamp 1698175906
transform 1 0 272048 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2481
timestamp 1698175906
transform 1 0 279216 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_2487
timestamp 1698175906
transform 1 0 279888 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2551
timestamp 1698175906
transform 1 0 287056 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_2557
timestamp 1698175906
transform 1 0 287728 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2621
timestamp 1698175906
transform 1 0 294896 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_2627
timestamp 1698175906
transform 1 0 295568 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_2643
timestamp 1698175906
transform 1 0 297360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_2651
timestamp 1698175906
transform 1 0 298256 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_352
timestamp 1698175906
transform 1 0 40768 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698175906
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698175906
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698175906
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_492
timestamp 1698175906
transform 1 0 56448 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_556
timestamp 1698175906
transform 1 0 63616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_562
timestamp 1698175906
transform 1 0 64288 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_626
timestamp 1698175906
transform 1 0 71456 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_632
timestamp 1698175906
transform 1 0 72128 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_696
timestamp 1698175906
transform 1 0 79296 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_702
timestamp 1698175906
transform 1 0 79968 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_766
timestamp 1698175906
transform 1 0 87136 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_772
timestamp 1698175906
transform 1 0 87808 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_836
timestamp 1698175906
transform 1 0 94976 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_842
timestamp 1698175906
transform 1 0 95648 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_906
timestamp 1698175906
transform 1 0 102816 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_912
timestamp 1698175906
transform 1 0 103488 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_976
timestamp 1698175906
transform 1 0 110656 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_982
timestamp 1698175906
transform 1 0 111328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1046
timestamp 1698175906
transform 1 0 118496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1052
timestamp 1698175906
transform 1 0 119168 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1116
timestamp 1698175906
transform 1 0 126336 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1122
timestamp 1698175906
transform 1 0 127008 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1186
timestamp 1698175906
transform 1 0 134176 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1192
timestamp 1698175906
transform 1 0 134848 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1256
timestamp 1698175906
transform 1 0 142016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1262
timestamp 1698175906
transform 1 0 142688 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1326
timestamp 1698175906
transform 1 0 149856 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1332
timestamp 1698175906
transform 1 0 150528 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1396
timestamp 1698175906
transform 1 0 157696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1402
timestamp 1698175906
transform 1 0 158368 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1466
timestamp 1698175906
transform 1 0 165536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1472
timestamp 1698175906
transform 1 0 166208 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1536
timestamp 1698175906
transform 1 0 173376 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1542
timestamp 1698175906
transform 1 0 174048 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1606
timestamp 1698175906
transform 1 0 181216 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1612
timestamp 1698175906
transform 1 0 181888 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1676
timestamp 1698175906
transform 1 0 189056 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1682
timestamp 1698175906
transform 1 0 189728 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1746
timestamp 1698175906
transform 1 0 196896 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1752
timestamp 1698175906
transform 1 0 197568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1816
timestamp 1698175906
transform 1 0 204736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1822
timestamp 1698175906
transform 1 0 205408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1886
timestamp 1698175906
transform 1 0 212576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1892
timestamp 1698175906
transform 1 0 213248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1956
timestamp 1698175906
transform 1 0 220416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1962
timestamp 1698175906
transform 1 0 221088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2026
timestamp 1698175906
transform 1 0 228256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2032
timestamp 1698175906
transform 1 0 228928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2096
timestamp 1698175906
transform 1 0 236096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2102
timestamp 1698175906
transform 1 0 236768 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2166
timestamp 1698175906
transform 1 0 243936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2172
timestamp 1698175906
transform 1 0 244608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2236
timestamp 1698175906
transform 1 0 251776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2242
timestamp 1698175906
transform 1 0 252448 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2306
timestamp 1698175906
transform 1 0 259616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2312
timestamp 1698175906
transform 1 0 260288 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2376
timestamp 1698175906
transform 1 0 267456 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2382
timestamp 1698175906
transform 1 0 268128 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2446
timestamp 1698175906
transform 1 0 275296 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2452
timestamp 1698175906
transform 1 0 275968 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2516
timestamp 1698175906
transform 1 0 283136 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2522
timestamp 1698175906
transform 1 0 283808 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2586
timestamp 1698175906
transform 1 0 290976 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_2592
timestamp 1698175906
transform 1 0 291648 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2624
timestamp 1698175906
transform 1 0 295232 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_2640
timestamp 1698175906
transform 1 0 297024 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2648
timestamp 1698175906
transform 1 0 297920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_381
timestamp 1698175906
transform 1 0 44016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698175906
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698175906
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_457
timestamp 1698175906
transform 1 0 52528 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_521
timestamp 1698175906
transform 1 0 59696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_527
timestamp 1698175906
transform 1 0 60368 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_591
timestamp 1698175906
transform 1 0 67536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_597
timestamp 1698175906
transform 1 0 68208 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_661
timestamp 1698175906
transform 1 0 75376 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_667
timestamp 1698175906
transform 1 0 76048 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_731
timestamp 1698175906
transform 1 0 83216 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_737
timestamp 1698175906
transform 1 0 83888 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_801
timestamp 1698175906
transform 1 0 91056 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_807
timestamp 1698175906
transform 1 0 91728 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_871
timestamp 1698175906
transform 1 0 98896 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_877
timestamp 1698175906
transform 1 0 99568 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_941
timestamp 1698175906
transform 1 0 106736 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_947
timestamp 1698175906
transform 1 0 107408 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1011
timestamp 1698175906
transform 1 0 114576 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1017
timestamp 1698175906
transform 1 0 115248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1081
timestamp 1698175906
transform 1 0 122416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1087
timestamp 1698175906
transform 1 0 123088 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1151
timestamp 1698175906
transform 1 0 130256 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1157
timestamp 1698175906
transform 1 0 130928 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1221
timestamp 1698175906
transform 1 0 138096 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1227
timestamp 1698175906
transform 1 0 138768 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1291
timestamp 1698175906
transform 1 0 145936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1297
timestamp 1698175906
transform 1 0 146608 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1361
timestamp 1698175906
transform 1 0 153776 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1367
timestamp 1698175906
transform 1 0 154448 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1431
timestamp 1698175906
transform 1 0 161616 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1437
timestamp 1698175906
transform 1 0 162288 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1501
timestamp 1698175906
transform 1 0 169456 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1507
timestamp 1698175906
transform 1 0 170128 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1571
timestamp 1698175906
transform 1 0 177296 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1577
timestamp 1698175906
transform 1 0 177968 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1641
timestamp 1698175906
transform 1 0 185136 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1647
timestamp 1698175906
transform 1 0 185808 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1711
timestamp 1698175906
transform 1 0 192976 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1717
timestamp 1698175906
transform 1 0 193648 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1781
timestamp 1698175906
transform 1 0 200816 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1787
timestamp 1698175906
transform 1 0 201488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1851
timestamp 1698175906
transform 1 0 208656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1857
timestamp 1698175906
transform 1 0 209328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1921
timestamp 1698175906
transform 1 0 216496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1927
timestamp 1698175906
transform 1 0 217168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1991
timestamp 1698175906
transform 1 0 224336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1997
timestamp 1698175906
transform 1 0 225008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2061
timestamp 1698175906
transform 1 0 232176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_2067
timestamp 1698175906
transform 1 0 232848 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2131
timestamp 1698175906
transform 1 0 240016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_2137
timestamp 1698175906
transform 1 0 240688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2201
timestamp 1698175906
transform 1 0 247856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_2207
timestamp 1698175906
transform 1 0 248528 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2271
timestamp 1698175906
transform 1 0 255696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_2277
timestamp 1698175906
transform 1 0 256368 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2341
timestamp 1698175906
transform 1 0 263536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_2347
timestamp 1698175906
transform 1 0 264208 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2411
timestamp 1698175906
transform 1 0 271376 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_2417
timestamp 1698175906
transform 1 0 272048 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2481
timestamp 1698175906
transform 1 0 279216 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_2487
timestamp 1698175906
transform 1 0 279888 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2551
timestamp 1698175906
transform 1 0 287056 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_2557
timestamp 1698175906
transform 1 0 287728 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2621
timestamp 1698175906
transform 1 0 294896 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_2627
timestamp 1698175906
transform 1 0 295568 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_2643
timestamp 1698175906
transform 1 0 297360 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_2651
timestamp 1698175906
transform 1 0 298256 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_352
timestamp 1698175906
transform 1 0 40768 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698175906
transform 1 0 47936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698175906
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698175906
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_492
timestamp 1698175906
transform 1 0 56448 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_556
timestamp 1698175906
transform 1 0 63616 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_562
timestamp 1698175906
transform 1 0 64288 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_626
timestamp 1698175906
transform 1 0 71456 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_632
timestamp 1698175906
transform 1 0 72128 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_696
timestamp 1698175906
transform 1 0 79296 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_702
timestamp 1698175906
transform 1 0 79968 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_766
timestamp 1698175906
transform 1 0 87136 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_772
timestamp 1698175906
transform 1 0 87808 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_836
timestamp 1698175906
transform 1 0 94976 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_842
timestamp 1698175906
transform 1 0 95648 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_906
timestamp 1698175906
transform 1 0 102816 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_912
timestamp 1698175906
transform 1 0 103488 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_976
timestamp 1698175906
transform 1 0 110656 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_982
timestamp 1698175906
transform 1 0 111328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1046
timestamp 1698175906
transform 1 0 118496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1052
timestamp 1698175906
transform 1 0 119168 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1116
timestamp 1698175906
transform 1 0 126336 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1122
timestamp 1698175906
transform 1 0 127008 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1186
timestamp 1698175906
transform 1 0 134176 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1192
timestamp 1698175906
transform 1 0 134848 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1256
timestamp 1698175906
transform 1 0 142016 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1262
timestamp 1698175906
transform 1 0 142688 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1326
timestamp 1698175906
transform 1 0 149856 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1332
timestamp 1698175906
transform 1 0 150528 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1396
timestamp 1698175906
transform 1 0 157696 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1402
timestamp 1698175906
transform 1 0 158368 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1466
timestamp 1698175906
transform 1 0 165536 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1472
timestamp 1698175906
transform 1 0 166208 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1536
timestamp 1698175906
transform 1 0 173376 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1542
timestamp 1698175906
transform 1 0 174048 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1606
timestamp 1698175906
transform 1 0 181216 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1612
timestamp 1698175906
transform 1 0 181888 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1676
timestamp 1698175906
transform 1 0 189056 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1682
timestamp 1698175906
transform 1 0 189728 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1746
timestamp 1698175906
transform 1 0 196896 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1752
timestamp 1698175906
transform 1 0 197568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1816
timestamp 1698175906
transform 1 0 204736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1822
timestamp 1698175906
transform 1 0 205408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1886
timestamp 1698175906
transform 1 0 212576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1892
timestamp 1698175906
transform 1 0 213248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1956
timestamp 1698175906
transform 1 0 220416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1962
timestamp 1698175906
transform 1 0 221088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2026
timestamp 1698175906
transform 1 0 228256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2032
timestamp 1698175906
transform 1 0 228928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2096
timestamp 1698175906
transform 1 0 236096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2102
timestamp 1698175906
transform 1 0 236768 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2166
timestamp 1698175906
transform 1 0 243936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2172
timestamp 1698175906
transform 1 0 244608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2236
timestamp 1698175906
transform 1 0 251776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2242
timestamp 1698175906
transform 1 0 252448 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2306
timestamp 1698175906
transform 1 0 259616 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2312
timestamp 1698175906
transform 1 0 260288 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2376
timestamp 1698175906
transform 1 0 267456 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2382
timestamp 1698175906
transform 1 0 268128 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2446
timestamp 1698175906
transform 1 0 275296 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2452
timestamp 1698175906
transform 1 0 275968 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2516
timestamp 1698175906
transform 1 0 283136 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2522
timestamp 1698175906
transform 1 0 283808 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2586
timestamp 1698175906
transform 1 0 290976 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_2592
timestamp 1698175906
transform 1 0 291648 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_2624
timestamp 1698175906
transform 1 0 295232 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_2640
timestamp 1698175906
transform 1 0 297024 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2648
timestamp 1698175906
transform 1 0 297920 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698175906
transform 1 0 44016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_387
timestamp 1698175906
transform 1 0 44688 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698175906
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_457
timestamp 1698175906
transform 1 0 52528 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_521
timestamp 1698175906
transform 1 0 59696 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_527
timestamp 1698175906
transform 1 0 60368 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_591
timestamp 1698175906
transform 1 0 67536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_597
timestamp 1698175906
transform 1 0 68208 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_661
timestamp 1698175906
transform 1 0 75376 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_667
timestamp 1698175906
transform 1 0 76048 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_731
timestamp 1698175906
transform 1 0 83216 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_737
timestamp 1698175906
transform 1 0 83888 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_801
timestamp 1698175906
transform 1 0 91056 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_807
timestamp 1698175906
transform 1 0 91728 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_871
timestamp 1698175906
transform 1 0 98896 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_877
timestamp 1698175906
transform 1 0 99568 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_941
timestamp 1698175906
transform 1 0 106736 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_947
timestamp 1698175906
transform 1 0 107408 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1011
timestamp 1698175906
transform 1 0 114576 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1017
timestamp 1698175906
transform 1 0 115248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1081
timestamp 1698175906
transform 1 0 122416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1087
timestamp 1698175906
transform 1 0 123088 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1151
timestamp 1698175906
transform 1 0 130256 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1157
timestamp 1698175906
transform 1 0 130928 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1221
timestamp 1698175906
transform 1 0 138096 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1227
timestamp 1698175906
transform 1 0 138768 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1291
timestamp 1698175906
transform 1 0 145936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1297
timestamp 1698175906
transform 1 0 146608 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1361
timestamp 1698175906
transform 1 0 153776 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1367
timestamp 1698175906
transform 1 0 154448 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1431
timestamp 1698175906
transform 1 0 161616 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1437
timestamp 1698175906
transform 1 0 162288 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1501
timestamp 1698175906
transform 1 0 169456 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1507
timestamp 1698175906
transform 1 0 170128 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1571
timestamp 1698175906
transform 1 0 177296 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1577
timestamp 1698175906
transform 1 0 177968 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1641
timestamp 1698175906
transform 1 0 185136 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1647
timestamp 1698175906
transform 1 0 185808 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1711
timestamp 1698175906
transform 1 0 192976 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1717
timestamp 1698175906
transform 1 0 193648 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1781
timestamp 1698175906
transform 1 0 200816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1787
timestamp 1698175906
transform 1 0 201488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1851
timestamp 1698175906
transform 1 0 208656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1857
timestamp 1698175906
transform 1 0 209328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1921
timestamp 1698175906
transform 1 0 216496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1927
timestamp 1698175906
transform 1 0 217168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1991
timestamp 1698175906
transform 1 0 224336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1997
timestamp 1698175906
transform 1 0 225008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2061
timestamp 1698175906
transform 1 0 232176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_2067
timestamp 1698175906
transform 1 0 232848 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2131
timestamp 1698175906
transform 1 0 240016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_2137
timestamp 1698175906
transform 1 0 240688 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2201
timestamp 1698175906
transform 1 0 247856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_2207
timestamp 1698175906
transform 1 0 248528 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2271
timestamp 1698175906
transform 1 0 255696 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_2277
timestamp 1698175906
transform 1 0 256368 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2341
timestamp 1698175906
transform 1 0 263536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_2347
timestamp 1698175906
transform 1 0 264208 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2411
timestamp 1698175906
transform 1 0 271376 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_2417
timestamp 1698175906
transform 1 0 272048 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2481
timestamp 1698175906
transform 1 0 279216 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_2487
timestamp 1698175906
transform 1 0 279888 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2551
timestamp 1698175906
transform 1 0 287056 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_2557
timestamp 1698175906
transform 1 0 287728 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2621
timestamp 1698175906
transform 1 0 294896 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_2627
timestamp 1698175906
transform 1 0 295568 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_2643
timestamp 1698175906
transform 1 0 297360 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_2651
timestamp 1698175906
transform 1 0 298256 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_352
timestamp 1698175906
transform 1 0 40768 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_416
timestamp 1698175906
transform 1 0 47936 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698175906
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698175906
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_492
timestamp 1698175906
transform 1 0 56448 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_556
timestamp 1698175906
transform 1 0 63616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_562
timestamp 1698175906
transform 1 0 64288 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_626
timestamp 1698175906
transform 1 0 71456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_632
timestamp 1698175906
transform 1 0 72128 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_696
timestamp 1698175906
transform 1 0 79296 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_702
timestamp 1698175906
transform 1 0 79968 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_766
timestamp 1698175906
transform 1 0 87136 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_772
timestamp 1698175906
transform 1 0 87808 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_836
timestamp 1698175906
transform 1 0 94976 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_842
timestamp 1698175906
transform 1 0 95648 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_906
timestamp 1698175906
transform 1 0 102816 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_912
timestamp 1698175906
transform 1 0 103488 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_976
timestamp 1698175906
transform 1 0 110656 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_982
timestamp 1698175906
transform 1 0 111328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1046
timestamp 1698175906
transform 1 0 118496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1052
timestamp 1698175906
transform 1 0 119168 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1116
timestamp 1698175906
transform 1 0 126336 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1122
timestamp 1698175906
transform 1 0 127008 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1186
timestamp 1698175906
transform 1 0 134176 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1192
timestamp 1698175906
transform 1 0 134848 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1256
timestamp 1698175906
transform 1 0 142016 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1262
timestamp 1698175906
transform 1 0 142688 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1326
timestamp 1698175906
transform 1 0 149856 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1332
timestamp 1698175906
transform 1 0 150528 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1396
timestamp 1698175906
transform 1 0 157696 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1402
timestamp 1698175906
transform 1 0 158368 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1466
timestamp 1698175906
transform 1 0 165536 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1472
timestamp 1698175906
transform 1 0 166208 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1536
timestamp 1698175906
transform 1 0 173376 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1542
timestamp 1698175906
transform 1 0 174048 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1606
timestamp 1698175906
transform 1 0 181216 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1612
timestamp 1698175906
transform 1 0 181888 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1676
timestamp 1698175906
transform 1 0 189056 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1682
timestamp 1698175906
transform 1 0 189728 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1746
timestamp 1698175906
transform 1 0 196896 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1752
timestamp 1698175906
transform 1 0 197568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1816
timestamp 1698175906
transform 1 0 204736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1822
timestamp 1698175906
transform 1 0 205408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1886
timestamp 1698175906
transform 1 0 212576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1892
timestamp 1698175906
transform 1 0 213248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1956
timestamp 1698175906
transform 1 0 220416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1962
timestamp 1698175906
transform 1 0 221088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2026
timestamp 1698175906
transform 1 0 228256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2032
timestamp 1698175906
transform 1 0 228928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2096
timestamp 1698175906
transform 1 0 236096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2102
timestamp 1698175906
transform 1 0 236768 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2166
timestamp 1698175906
transform 1 0 243936 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2172
timestamp 1698175906
transform 1 0 244608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2236
timestamp 1698175906
transform 1 0 251776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2242
timestamp 1698175906
transform 1 0 252448 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2306
timestamp 1698175906
transform 1 0 259616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2312
timestamp 1698175906
transform 1 0 260288 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2376
timestamp 1698175906
transform 1 0 267456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2382
timestamp 1698175906
transform 1 0 268128 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2446
timestamp 1698175906
transform 1 0 275296 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2452
timestamp 1698175906
transform 1 0 275968 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2516
timestamp 1698175906
transform 1 0 283136 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2522
timestamp 1698175906
transform 1 0 283808 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2586
timestamp 1698175906
transform 1 0 290976 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_2592
timestamp 1698175906
transform 1 0 291648 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_2624
timestamp 1698175906
transform 1 0 295232 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_2640
timestamp 1698175906
transform 1 0 297024 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2648
timestamp 1698175906
transform 1 0 297920 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_381
timestamp 1698175906
transform 1 0 44016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_387
timestamp 1698175906
transform 1 0 44688 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1698175906
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_457
timestamp 1698175906
transform 1 0 52528 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_521
timestamp 1698175906
transform 1 0 59696 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_527
timestamp 1698175906
transform 1 0 60368 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_591
timestamp 1698175906
transform 1 0 67536 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_597
timestamp 1698175906
transform 1 0 68208 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_661
timestamp 1698175906
transform 1 0 75376 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_667
timestamp 1698175906
transform 1 0 76048 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_731
timestamp 1698175906
transform 1 0 83216 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_737
timestamp 1698175906
transform 1 0 83888 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_801
timestamp 1698175906
transform 1 0 91056 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_807
timestamp 1698175906
transform 1 0 91728 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_871
timestamp 1698175906
transform 1 0 98896 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_877
timestamp 1698175906
transform 1 0 99568 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_941
timestamp 1698175906
transform 1 0 106736 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_947
timestamp 1698175906
transform 1 0 107408 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1011
timestamp 1698175906
transform 1 0 114576 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1017
timestamp 1698175906
transform 1 0 115248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1081
timestamp 1698175906
transform 1 0 122416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1087
timestamp 1698175906
transform 1 0 123088 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1151
timestamp 1698175906
transform 1 0 130256 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1157
timestamp 1698175906
transform 1 0 130928 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1221
timestamp 1698175906
transform 1 0 138096 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1227
timestamp 1698175906
transform 1 0 138768 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1291
timestamp 1698175906
transform 1 0 145936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1297
timestamp 1698175906
transform 1 0 146608 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1361
timestamp 1698175906
transform 1 0 153776 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1367
timestamp 1698175906
transform 1 0 154448 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1431
timestamp 1698175906
transform 1 0 161616 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1437
timestamp 1698175906
transform 1 0 162288 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1501
timestamp 1698175906
transform 1 0 169456 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1507
timestamp 1698175906
transform 1 0 170128 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1571
timestamp 1698175906
transform 1 0 177296 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1577
timestamp 1698175906
transform 1 0 177968 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1641
timestamp 1698175906
transform 1 0 185136 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1647
timestamp 1698175906
transform 1 0 185808 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1711
timestamp 1698175906
transform 1 0 192976 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1717
timestamp 1698175906
transform 1 0 193648 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1781
timestamp 1698175906
transform 1 0 200816 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1787
timestamp 1698175906
transform 1 0 201488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1851
timestamp 1698175906
transform 1 0 208656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1857
timestamp 1698175906
transform 1 0 209328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1921
timestamp 1698175906
transform 1 0 216496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1927
timestamp 1698175906
transform 1 0 217168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1991
timestamp 1698175906
transform 1 0 224336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1997
timestamp 1698175906
transform 1 0 225008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2061
timestamp 1698175906
transform 1 0 232176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_2067
timestamp 1698175906
transform 1 0 232848 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2131
timestamp 1698175906
transform 1 0 240016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_2137
timestamp 1698175906
transform 1 0 240688 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2201
timestamp 1698175906
transform 1 0 247856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_2207
timestamp 1698175906
transform 1 0 248528 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2271
timestamp 1698175906
transform 1 0 255696 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_2277
timestamp 1698175906
transform 1 0 256368 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2341
timestamp 1698175906
transform 1 0 263536 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_2347
timestamp 1698175906
transform 1 0 264208 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2411
timestamp 1698175906
transform 1 0 271376 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_2417
timestamp 1698175906
transform 1 0 272048 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2481
timestamp 1698175906
transform 1 0 279216 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_2487
timestamp 1698175906
transform 1 0 279888 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2551
timestamp 1698175906
transform 1 0 287056 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_2557
timestamp 1698175906
transform 1 0 287728 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2621
timestamp 1698175906
transform 1 0 294896 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_2627
timestamp 1698175906
transform 1 0 295568 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_2643
timestamp 1698175906
transform 1 0 297360 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_2651
timestamp 1698175906
transform 1 0 298256 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_352
timestamp 1698175906
transform 1 0 40768 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_416
timestamp 1698175906
transform 1 0 47936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698175906
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698175906
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_492
timestamp 1698175906
transform 1 0 56448 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_556
timestamp 1698175906
transform 1 0 63616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_562
timestamp 1698175906
transform 1 0 64288 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_626
timestamp 1698175906
transform 1 0 71456 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_632
timestamp 1698175906
transform 1 0 72128 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_696
timestamp 1698175906
transform 1 0 79296 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_702
timestamp 1698175906
transform 1 0 79968 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_766
timestamp 1698175906
transform 1 0 87136 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_772
timestamp 1698175906
transform 1 0 87808 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_836
timestamp 1698175906
transform 1 0 94976 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_842
timestamp 1698175906
transform 1 0 95648 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_906
timestamp 1698175906
transform 1 0 102816 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_912
timestamp 1698175906
transform 1 0 103488 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_976
timestamp 1698175906
transform 1 0 110656 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_982
timestamp 1698175906
transform 1 0 111328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1046
timestamp 1698175906
transform 1 0 118496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1052
timestamp 1698175906
transform 1 0 119168 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1116
timestamp 1698175906
transform 1 0 126336 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1122
timestamp 1698175906
transform 1 0 127008 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1186
timestamp 1698175906
transform 1 0 134176 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1192
timestamp 1698175906
transform 1 0 134848 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1256
timestamp 1698175906
transform 1 0 142016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1262
timestamp 1698175906
transform 1 0 142688 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1326
timestamp 1698175906
transform 1 0 149856 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1332
timestamp 1698175906
transform 1 0 150528 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1396
timestamp 1698175906
transform 1 0 157696 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1402
timestamp 1698175906
transform 1 0 158368 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1466
timestamp 1698175906
transform 1 0 165536 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1472
timestamp 1698175906
transform 1 0 166208 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1536
timestamp 1698175906
transform 1 0 173376 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1542
timestamp 1698175906
transform 1 0 174048 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1606
timestamp 1698175906
transform 1 0 181216 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1612
timestamp 1698175906
transform 1 0 181888 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1676
timestamp 1698175906
transform 1 0 189056 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1682
timestamp 1698175906
transform 1 0 189728 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1746
timestamp 1698175906
transform 1 0 196896 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1752
timestamp 1698175906
transform 1 0 197568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1816
timestamp 1698175906
transform 1 0 204736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1822
timestamp 1698175906
transform 1 0 205408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1886
timestamp 1698175906
transform 1 0 212576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1892
timestamp 1698175906
transform 1 0 213248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1956
timestamp 1698175906
transform 1 0 220416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1962
timestamp 1698175906
transform 1 0 221088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2026
timestamp 1698175906
transform 1 0 228256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2032
timestamp 1698175906
transform 1 0 228928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2096
timestamp 1698175906
transform 1 0 236096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2102
timestamp 1698175906
transform 1 0 236768 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2166
timestamp 1698175906
transform 1 0 243936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2172
timestamp 1698175906
transform 1 0 244608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2236
timestamp 1698175906
transform 1 0 251776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2242
timestamp 1698175906
transform 1 0 252448 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2306
timestamp 1698175906
transform 1 0 259616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2312
timestamp 1698175906
transform 1 0 260288 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2376
timestamp 1698175906
transform 1 0 267456 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2382
timestamp 1698175906
transform 1 0 268128 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2446
timestamp 1698175906
transform 1 0 275296 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2452
timestamp 1698175906
transform 1 0 275968 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2516
timestamp 1698175906
transform 1 0 283136 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2522
timestamp 1698175906
transform 1 0 283808 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2586
timestamp 1698175906
transform 1 0 290976 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_2592
timestamp 1698175906
transform 1 0 291648 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_2624
timestamp 1698175906
transform 1 0 295232 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_2640
timestamp 1698175906
transform 1 0 297024 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2648
timestamp 1698175906
transform 1 0 297920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698175906
transform 1 0 44016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_387
timestamp 1698175906
transform 1 0 44688 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_451
timestamp 1698175906
transform 1 0 51856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_457
timestamp 1698175906
transform 1 0 52528 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_521
timestamp 1698175906
transform 1 0 59696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_527
timestamp 1698175906
transform 1 0 60368 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_591
timestamp 1698175906
transform 1 0 67536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_597
timestamp 1698175906
transform 1 0 68208 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_661
timestamp 1698175906
transform 1 0 75376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_667
timestamp 1698175906
transform 1 0 76048 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_731
timestamp 1698175906
transform 1 0 83216 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_737
timestamp 1698175906
transform 1 0 83888 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_801
timestamp 1698175906
transform 1 0 91056 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_807
timestamp 1698175906
transform 1 0 91728 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_871
timestamp 1698175906
transform 1 0 98896 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_877
timestamp 1698175906
transform 1 0 99568 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_941
timestamp 1698175906
transform 1 0 106736 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_947
timestamp 1698175906
transform 1 0 107408 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1011
timestamp 1698175906
transform 1 0 114576 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1017
timestamp 1698175906
transform 1 0 115248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1081
timestamp 1698175906
transform 1 0 122416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1087
timestamp 1698175906
transform 1 0 123088 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1151
timestamp 1698175906
transform 1 0 130256 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1157
timestamp 1698175906
transform 1 0 130928 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1221
timestamp 1698175906
transform 1 0 138096 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1227
timestamp 1698175906
transform 1 0 138768 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1291
timestamp 1698175906
transform 1 0 145936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1297
timestamp 1698175906
transform 1 0 146608 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1361
timestamp 1698175906
transform 1 0 153776 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1367
timestamp 1698175906
transform 1 0 154448 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1431
timestamp 1698175906
transform 1 0 161616 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1437
timestamp 1698175906
transform 1 0 162288 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1501
timestamp 1698175906
transform 1 0 169456 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1507
timestamp 1698175906
transform 1 0 170128 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1571
timestamp 1698175906
transform 1 0 177296 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1577
timestamp 1698175906
transform 1 0 177968 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1641
timestamp 1698175906
transform 1 0 185136 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1647
timestamp 1698175906
transform 1 0 185808 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1711
timestamp 1698175906
transform 1 0 192976 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1717
timestamp 1698175906
transform 1 0 193648 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1781
timestamp 1698175906
transform 1 0 200816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1787
timestamp 1698175906
transform 1 0 201488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1851
timestamp 1698175906
transform 1 0 208656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1857
timestamp 1698175906
transform 1 0 209328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1921
timestamp 1698175906
transform 1 0 216496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1927
timestamp 1698175906
transform 1 0 217168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1991
timestamp 1698175906
transform 1 0 224336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1997
timestamp 1698175906
transform 1 0 225008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2061
timestamp 1698175906
transform 1 0 232176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_2067
timestamp 1698175906
transform 1 0 232848 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2131
timestamp 1698175906
transform 1 0 240016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_2137
timestamp 1698175906
transform 1 0 240688 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2201
timestamp 1698175906
transform 1 0 247856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_2207
timestamp 1698175906
transform 1 0 248528 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2271
timestamp 1698175906
transform 1 0 255696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_2277
timestamp 1698175906
transform 1 0 256368 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2341
timestamp 1698175906
transform 1 0 263536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_2347
timestamp 1698175906
transform 1 0 264208 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2411
timestamp 1698175906
transform 1 0 271376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_2417
timestamp 1698175906
transform 1 0 272048 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2481
timestamp 1698175906
transform 1 0 279216 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_2487
timestamp 1698175906
transform 1 0 279888 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2551
timestamp 1698175906
transform 1 0 287056 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_2557
timestamp 1698175906
transform 1 0 287728 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2621
timestamp 1698175906
transform 1 0 294896 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_2627
timestamp 1698175906
transform 1 0 295568 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_2643
timestamp 1698175906
transform 1 0 297360 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_2651
timestamp 1698175906
transform 1 0 298256 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_352
timestamp 1698175906
transform 1 0 40768 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1698175906
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_422
timestamp 1698175906
transform 1 0 48608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698175906
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_492
timestamp 1698175906
transform 1 0 56448 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_556
timestamp 1698175906
transform 1 0 63616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_562
timestamp 1698175906
transform 1 0 64288 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_626
timestamp 1698175906
transform 1 0 71456 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_632
timestamp 1698175906
transform 1 0 72128 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_696
timestamp 1698175906
transform 1 0 79296 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_702
timestamp 1698175906
transform 1 0 79968 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_766
timestamp 1698175906
transform 1 0 87136 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_772
timestamp 1698175906
transform 1 0 87808 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_836
timestamp 1698175906
transform 1 0 94976 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_842
timestamp 1698175906
transform 1 0 95648 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_906
timestamp 1698175906
transform 1 0 102816 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_912
timestamp 1698175906
transform 1 0 103488 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_976
timestamp 1698175906
transform 1 0 110656 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_982
timestamp 1698175906
transform 1 0 111328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1046
timestamp 1698175906
transform 1 0 118496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1052
timestamp 1698175906
transform 1 0 119168 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1116
timestamp 1698175906
transform 1 0 126336 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1122
timestamp 1698175906
transform 1 0 127008 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1186
timestamp 1698175906
transform 1 0 134176 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1192
timestamp 1698175906
transform 1 0 134848 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1256
timestamp 1698175906
transform 1 0 142016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1262
timestamp 1698175906
transform 1 0 142688 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1326
timestamp 1698175906
transform 1 0 149856 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1332
timestamp 1698175906
transform 1 0 150528 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1396
timestamp 1698175906
transform 1 0 157696 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1402
timestamp 1698175906
transform 1 0 158368 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1466
timestamp 1698175906
transform 1 0 165536 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1472
timestamp 1698175906
transform 1 0 166208 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1536
timestamp 1698175906
transform 1 0 173376 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1542
timestamp 1698175906
transform 1 0 174048 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1606
timestamp 1698175906
transform 1 0 181216 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1612
timestamp 1698175906
transform 1 0 181888 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1676
timestamp 1698175906
transform 1 0 189056 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1682
timestamp 1698175906
transform 1 0 189728 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1746
timestamp 1698175906
transform 1 0 196896 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1752
timestamp 1698175906
transform 1 0 197568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1816
timestamp 1698175906
transform 1 0 204736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1822
timestamp 1698175906
transform 1 0 205408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1886
timestamp 1698175906
transform 1 0 212576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1892
timestamp 1698175906
transform 1 0 213248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1956
timestamp 1698175906
transform 1 0 220416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1962
timestamp 1698175906
transform 1 0 221088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2026
timestamp 1698175906
transform 1 0 228256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2032
timestamp 1698175906
transform 1 0 228928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2096
timestamp 1698175906
transform 1 0 236096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2102
timestamp 1698175906
transform 1 0 236768 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2166
timestamp 1698175906
transform 1 0 243936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2172
timestamp 1698175906
transform 1 0 244608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2236
timestamp 1698175906
transform 1 0 251776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2242
timestamp 1698175906
transform 1 0 252448 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2306
timestamp 1698175906
transform 1 0 259616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2312
timestamp 1698175906
transform 1 0 260288 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2376
timestamp 1698175906
transform 1 0 267456 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2382
timestamp 1698175906
transform 1 0 268128 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2446
timestamp 1698175906
transform 1 0 275296 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2452
timestamp 1698175906
transform 1 0 275968 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2516
timestamp 1698175906
transform 1 0 283136 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2522
timestamp 1698175906
transform 1 0 283808 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2586
timestamp 1698175906
transform 1 0 290976 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_2592
timestamp 1698175906
transform 1 0 291648 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_2624
timestamp 1698175906
transform 1 0 295232 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_2640
timestamp 1698175906
transform 1 0 297024 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2648
timestamp 1698175906
transform 1 0 297920 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_381
timestamp 1698175906
transform 1 0 44016 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_387
timestamp 1698175906
transform 1 0 44688 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_451
timestamp 1698175906
transform 1 0 51856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_457
timestamp 1698175906
transform 1 0 52528 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_521
timestamp 1698175906
transform 1 0 59696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_527
timestamp 1698175906
transform 1 0 60368 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_591
timestamp 1698175906
transform 1 0 67536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_597
timestamp 1698175906
transform 1 0 68208 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_661
timestamp 1698175906
transform 1 0 75376 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_667
timestamp 1698175906
transform 1 0 76048 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_731
timestamp 1698175906
transform 1 0 83216 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_737
timestamp 1698175906
transform 1 0 83888 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_801
timestamp 1698175906
transform 1 0 91056 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_807
timestamp 1698175906
transform 1 0 91728 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_871
timestamp 1698175906
transform 1 0 98896 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_877
timestamp 1698175906
transform 1 0 99568 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_941
timestamp 1698175906
transform 1 0 106736 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_947
timestamp 1698175906
transform 1 0 107408 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1011
timestamp 1698175906
transform 1 0 114576 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1017
timestamp 1698175906
transform 1 0 115248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1081
timestamp 1698175906
transform 1 0 122416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1087
timestamp 1698175906
transform 1 0 123088 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1151
timestamp 1698175906
transform 1 0 130256 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1157
timestamp 1698175906
transform 1 0 130928 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1221
timestamp 1698175906
transform 1 0 138096 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1227
timestamp 1698175906
transform 1 0 138768 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1291
timestamp 1698175906
transform 1 0 145936 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1297
timestamp 1698175906
transform 1 0 146608 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1361
timestamp 1698175906
transform 1 0 153776 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1367
timestamp 1698175906
transform 1 0 154448 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1431
timestamp 1698175906
transform 1 0 161616 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1437
timestamp 1698175906
transform 1 0 162288 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1501
timestamp 1698175906
transform 1 0 169456 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1507
timestamp 1698175906
transform 1 0 170128 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1571
timestamp 1698175906
transform 1 0 177296 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1577
timestamp 1698175906
transform 1 0 177968 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1641
timestamp 1698175906
transform 1 0 185136 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1647
timestamp 1698175906
transform 1 0 185808 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1711
timestamp 1698175906
transform 1 0 192976 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1717
timestamp 1698175906
transform 1 0 193648 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1781
timestamp 1698175906
transform 1 0 200816 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1787
timestamp 1698175906
transform 1 0 201488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1851
timestamp 1698175906
transform 1 0 208656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1857
timestamp 1698175906
transform 1 0 209328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1921
timestamp 1698175906
transform 1 0 216496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1927
timestamp 1698175906
transform 1 0 217168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1991
timestamp 1698175906
transform 1 0 224336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1997
timestamp 1698175906
transform 1 0 225008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2061
timestamp 1698175906
transform 1 0 232176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_2067
timestamp 1698175906
transform 1 0 232848 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2131
timestamp 1698175906
transform 1 0 240016 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_2137
timestamp 1698175906
transform 1 0 240688 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2201
timestamp 1698175906
transform 1 0 247856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_2207
timestamp 1698175906
transform 1 0 248528 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2271
timestamp 1698175906
transform 1 0 255696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_2277
timestamp 1698175906
transform 1 0 256368 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2341
timestamp 1698175906
transform 1 0 263536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_2347
timestamp 1698175906
transform 1 0 264208 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2411
timestamp 1698175906
transform 1 0 271376 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_2417
timestamp 1698175906
transform 1 0 272048 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2481
timestamp 1698175906
transform 1 0 279216 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_2487
timestamp 1698175906
transform 1 0 279888 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2551
timestamp 1698175906
transform 1 0 287056 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_2557
timestamp 1698175906
transform 1 0 287728 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2621
timestamp 1698175906
transform 1 0 294896 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_2627
timestamp 1698175906
transform 1 0 295568 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_2643
timestamp 1698175906
transform 1 0 297360 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_2651
timestamp 1698175906
transform 1 0 298256 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_352
timestamp 1698175906
transform 1 0 40768 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698175906
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_422
timestamp 1698175906
transform 1 0 48608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698175906
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_492
timestamp 1698175906
transform 1 0 56448 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_556
timestamp 1698175906
transform 1 0 63616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_562
timestamp 1698175906
transform 1 0 64288 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_626
timestamp 1698175906
transform 1 0 71456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_632
timestamp 1698175906
transform 1 0 72128 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_696
timestamp 1698175906
transform 1 0 79296 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_702
timestamp 1698175906
transform 1 0 79968 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_766
timestamp 1698175906
transform 1 0 87136 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_772
timestamp 1698175906
transform 1 0 87808 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_836
timestamp 1698175906
transform 1 0 94976 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_842
timestamp 1698175906
transform 1 0 95648 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_906
timestamp 1698175906
transform 1 0 102816 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_912
timestamp 1698175906
transform 1 0 103488 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_976
timestamp 1698175906
transform 1 0 110656 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_982
timestamp 1698175906
transform 1 0 111328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1046
timestamp 1698175906
transform 1 0 118496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1052
timestamp 1698175906
transform 1 0 119168 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1116
timestamp 1698175906
transform 1 0 126336 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1122
timestamp 1698175906
transform 1 0 127008 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1186
timestamp 1698175906
transform 1 0 134176 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1192
timestamp 1698175906
transform 1 0 134848 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1256
timestamp 1698175906
transform 1 0 142016 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1262
timestamp 1698175906
transform 1 0 142688 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1326
timestamp 1698175906
transform 1 0 149856 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1332
timestamp 1698175906
transform 1 0 150528 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1396
timestamp 1698175906
transform 1 0 157696 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1402
timestamp 1698175906
transform 1 0 158368 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1466
timestamp 1698175906
transform 1 0 165536 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1472
timestamp 1698175906
transform 1 0 166208 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1536
timestamp 1698175906
transform 1 0 173376 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1542
timestamp 1698175906
transform 1 0 174048 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1606
timestamp 1698175906
transform 1 0 181216 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1612
timestamp 1698175906
transform 1 0 181888 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1676
timestamp 1698175906
transform 1 0 189056 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1682
timestamp 1698175906
transform 1 0 189728 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1746
timestamp 1698175906
transform 1 0 196896 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1752
timestamp 1698175906
transform 1 0 197568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1816
timestamp 1698175906
transform 1 0 204736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1822
timestamp 1698175906
transform 1 0 205408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1886
timestamp 1698175906
transform 1 0 212576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1892
timestamp 1698175906
transform 1 0 213248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1956
timestamp 1698175906
transform 1 0 220416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1962
timestamp 1698175906
transform 1 0 221088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2026
timestamp 1698175906
transform 1 0 228256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2032
timestamp 1698175906
transform 1 0 228928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2096
timestamp 1698175906
transform 1 0 236096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2102
timestamp 1698175906
transform 1 0 236768 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2166
timestamp 1698175906
transform 1 0 243936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2172
timestamp 1698175906
transform 1 0 244608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2236
timestamp 1698175906
transform 1 0 251776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2242
timestamp 1698175906
transform 1 0 252448 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2306
timestamp 1698175906
transform 1 0 259616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2312
timestamp 1698175906
transform 1 0 260288 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2376
timestamp 1698175906
transform 1 0 267456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2382
timestamp 1698175906
transform 1 0 268128 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2446
timestamp 1698175906
transform 1 0 275296 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2452
timestamp 1698175906
transform 1 0 275968 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2516
timestamp 1698175906
transform 1 0 283136 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2522
timestamp 1698175906
transform 1 0 283808 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2586
timestamp 1698175906
transform 1 0 290976 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_2592
timestamp 1698175906
transform 1 0 291648 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_2624
timestamp 1698175906
transform 1 0 295232 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_2640
timestamp 1698175906
transform 1 0 297024 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2648
timestamp 1698175906
transform 1 0 297920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_381
timestamp 1698175906
transform 1 0 44016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_387
timestamp 1698175906
transform 1 0 44688 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_451
timestamp 1698175906
transform 1 0 51856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_457
timestamp 1698175906
transform 1 0 52528 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_521
timestamp 1698175906
transform 1 0 59696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_527
timestamp 1698175906
transform 1 0 60368 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_591
timestamp 1698175906
transform 1 0 67536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_597
timestamp 1698175906
transform 1 0 68208 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_661
timestamp 1698175906
transform 1 0 75376 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_667
timestamp 1698175906
transform 1 0 76048 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_731
timestamp 1698175906
transform 1 0 83216 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_737
timestamp 1698175906
transform 1 0 83888 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_801
timestamp 1698175906
transform 1 0 91056 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_807
timestamp 1698175906
transform 1 0 91728 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_871
timestamp 1698175906
transform 1 0 98896 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_877
timestamp 1698175906
transform 1 0 99568 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_941
timestamp 1698175906
transform 1 0 106736 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_947
timestamp 1698175906
transform 1 0 107408 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1011
timestamp 1698175906
transform 1 0 114576 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1017
timestamp 1698175906
transform 1 0 115248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1081
timestamp 1698175906
transform 1 0 122416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1087
timestamp 1698175906
transform 1 0 123088 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1151
timestamp 1698175906
transform 1 0 130256 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1157
timestamp 1698175906
transform 1 0 130928 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1221
timestamp 1698175906
transform 1 0 138096 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1227
timestamp 1698175906
transform 1 0 138768 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1291
timestamp 1698175906
transform 1 0 145936 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1297
timestamp 1698175906
transform 1 0 146608 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1361
timestamp 1698175906
transform 1 0 153776 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1367
timestamp 1698175906
transform 1 0 154448 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1431
timestamp 1698175906
transform 1 0 161616 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1437
timestamp 1698175906
transform 1 0 162288 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1501
timestamp 1698175906
transform 1 0 169456 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1507
timestamp 1698175906
transform 1 0 170128 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1571
timestamp 1698175906
transform 1 0 177296 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1577
timestamp 1698175906
transform 1 0 177968 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1641
timestamp 1698175906
transform 1 0 185136 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1647
timestamp 1698175906
transform 1 0 185808 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1711
timestamp 1698175906
transform 1 0 192976 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1717
timestamp 1698175906
transform 1 0 193648 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1781
timestamp 1698175906
transform 1 0 200816 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1787
timestamp 1698175906
transform 1 0 201488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1851
timestamp 1698175906
transform 1 0 208656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1857
timestamp 1698175906
transform 1 0 209328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1921
timestamp 1698175906
transform 1 0 216496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1927
timestamp 1698175906
transform 1 0 217168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1991
timestamp 1698175906
transform 1 0 224336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1997
timestamp 1698175906
transform 1 0 225008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2061
timestamp 1698175906
transform 1 0 232176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_2067
timestamp 1698175906
transform 1 0 232848 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2131
timestamp 1698175906
transform 1 0 240016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_2137
timestamp 1698175906
transform 1 0 240688 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2201
timestamp 1698175906
transform 1 0 247856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_2207
timestamp 1698175906
transform 1 0 248528 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2271
timestamp 1698175906
transform 1 0 255696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_2277
timestamp 1698175906
transform 1 0 256368 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2341
timestamp 1698175906
transform 1 0 263536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_2347
timestamp 1698175906
transform 1 0 264208 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2411
timestamp 1698175906
transform 1 0 271376 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_2417
timestamp 1698175906
transform 1 0 272048 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2481
timestamp 1698175906
transform 1 0 279216 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_2487
timestamp 1698175906
transform 1 0 279888 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2551
timestamp 1698175906
transform 1 0 287056 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_2557
timestamp 1698175906
transform 1 0 287728 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2621
timestamp 1698175906
transform 1 0 294896 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_2627
timestamp 1698175906
transform 1 0 295568 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_2643
timestamp 1698175906
transform 1 0 297360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_2651
timestamp 1698175906
transform 1 0 298256 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698175906
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698175906
transform 1 0 40768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698175906
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698175906
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698175906
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_492
timestamp 1698175906
transform 1 0 56448 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_556
timestamp 1698175906
transform 1 0 63616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_562
timestamp 1698175906
transform 1 0 64288 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_626
timestamp 1698175906
transform 1 0 71456 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_632
timestamp 1698175906
transform 1 0 72128 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_696
timestamp 1698175906
transform 1 0 79296 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_702
timestamp 1698175906
transform 1 0 79968 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_766
timestamp 1698175906
transform 1 0 87136 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_772
timestamp 1698175906
transform 1 0 87808 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_836
timestamp 1698175906
transform 1 0 94976 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_842
timestamp 1698175906
transform 1 0 95648 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_906
timestamp 1698175906
transform 1 0 102816 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_912
timestamp 1698175906
transform 1 0 103488 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_976
timestamp 1698175906
transform 1 0 110656 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_982
timestamp 1698175906
transform 1 0 111328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1046
timestamp 1698175906
transform 1 0 118496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1052
timestamp 1698175906
transform 1 0 119168 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1116
timestamp 1698175906
transform 1 0 126336 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1122
timestamp 1698175906
transform 1 0 127008 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1186
timestamp 1698175906
transform 1 0 134176 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1192
timestamp 1698175906
transform 1 0 134848 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1256
timestamp 1698175906
transform 1 0 142016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1262
timestamp 1698175906
transform 1 0 142688 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1326
timestamp 1698175906
transform 1 0 149856 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1332
timestamp 1698175906
transform 1 0 150528 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1396
timestamp 1698175906
transform 1 0 157696 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1402
timestamp 1698175906
transform 1 0 158368 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1466
timestamp 1698175906
transform 1 0 165536 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1472
timestamp 1698175906
transform 1 0 166208 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1536
timestamp 1698175906
transform 1 0 173376 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1542
timestamp 1698175906
transform 1 0 174048 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1606
timestamp 1698175906
transform 1 0 181216 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1612
timestamp 1698175906
transform 1 0 181888 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1676
timestamp 1698175906
transform 1 0 189056 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1682
timestamp 1698175906
transform 1 0 189728 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1746
timestamp 1698175906
transform 1 0 196896 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1752
timestamp 1698175906
transform 1 0 197568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1816
timestamp 1698175906
transform 1 0 204736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1822
timestamp 1698175906
transform 1 0 205408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1886
timestamp 1698175906
transform 1 0 212576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1892
timestamp 1698175906
transform 1 0 213248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1956
timestamp 1698175906
transform 1 0 220416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1962
timestamp 1698175906
transform 1 0 221088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2026
timestamp 1698175906
transform 1 0 228256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2032
timestamp 1698175906
transform 1 0 228928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2096
timestamp 1698175906
transform 1 0 236096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2102
timestamp 1698175906
transform 1 0 236768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2166
timestamp 1698175906
transform 1 0 243936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2172
timestamp 1698175906
transform 1 0 244608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2236
timestamp 1698175906
transform 1 0 251776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2242
timestamp 1698175906
transform 1 0 252448 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2306
timestamp 1698175906
transform 1 0 259616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2312
timestamp 1698175906
transform 1 0 260288 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2376
timestamp 1698175906
transform 1 0 267456 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2382
timestamp 1698175906
transform 1 0 268128 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2446
timestamp 1698175906
transform 1 0 275296 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2452
timestamp 1698175906
transform 1 0 275968 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2516
timestamp 1698175906
transform 1 0 283136 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2522
timestamp 1698175906
transform 1 0 283808 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2586
timestamp 1698175906
transform 1 0 290976 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_2592
timestamp 1698175906
transform 1 0 291648 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_2624
timestamp 1698175906
transform 1 0 295232 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_2640
timestamp 1698175906
transform 1 0 297024 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2648
timestamp 1698175906
transform 1 0 297920 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698175906
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698175906
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698175906
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698175906
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698175906
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698175906
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698175906
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698175906
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_317
timestamp 1698175906
transform 1 0 36848 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_381
timestamp 1698175906
transform 1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698175906
transform 1 0 44688 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698175906
transform 1 0 51856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_457
timestamp 1698175906
transform 1 0 52528 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_521
timestamp 1698175906
transform 1 0 59696 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_527
timestamp 1698175906
transform 1 0 60368 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_591
timestamp 1698175906
transform 1 0 67536 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_597
timestamp 1698175906
transform 1 0 68208 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_661
timestamp 1698175906
transform 1 0 75376 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_667
timestamp 1698175906
transform 1 0 76048 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_731
timestamp 1698175906
transform 1 0 83216 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_737
timestamp 1698175906
transform 1 0 83888 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_801
timestamp 1698175906
transform 1 0 91056 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_807
timestamp 1698175906
transform 1 0 91728 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_871
timestamp 1698175906
transform 1 0 98896 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_877
timestamp 1698175906
transform 1 0 99568 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_941
timestamp 1698175906
transform 1 0 106736 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_947
timestamp 1698175906
transform 1 0 107408 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1011
timestamp 1698175906
transform 1 0 114576 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1017
timestamp 1698175906
transform 1 0 115248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1081
timestamp 1698175906
transform 1 0 122416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1087
timestamp 1698175906
transform 1 0 123088 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1151
timestamp 1698175906
transform 1 0 130256 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1157
timestamp 1698175906
transform 1 0 130928 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1221
timestamp 1698175906
transform 1 0 138096 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1227
timestamp 1698175906
transform 1 0 138768 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1291
timestamp 1698175906
transform 1 0 145936 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1297
timestamp 1698175906
transform 1 0 146608 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1361
timestamp 1698175906
transform 1 0 153776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1367
timestamp 1698175906
transform 1 0 154448 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1431
timestamp 1698175906
transform 1 0 161616 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1437
timestamp 1698175906
transform 1 0 162288 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1501
timestamp 1698175906
transform 1 0 169456 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1507
timestamp 1698175906
transform 1 0 170128 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1571
timestamp 1698175906
transform 1 0 177296 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1577
timestamp 1698175906
transform 1 0 177968 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1641
timestamp 1698175906
transform 1 0 185136 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1647
timestamp 1698175906
transform 1 0 185808 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1711
timestamp 1698175906
transform 1 0 192976 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1717
timestamp 1698175906
transform 1 0 193648 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1781
timestamp 1698175906
transform 1 0 200816 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1787
timestamp 1698175906
transform 1 0 201488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1851
timestamp 1698175906
transform 1 0 208656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1857
timestamp 1698175906
transform 1 0 209328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1921
timestamp 1698175906
transform 1 0 216496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1927
timestamp 1698175906
transform 1 0 217168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1991
timestamp 1698175906
transform 1 0 224336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1997
timestamp 1698175906
transform 1 0 225008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2061
timestamp 1698175906
transform 1 0 232176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_2067
timestamp 1698175906
transform 1 0 232848 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2131
timestamp 1698175906
transform 1 0 240016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_2137
timestamp 1698175906
transform 1 0 240688 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2201
timestamp 1698175906
transform 1 0 247856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_2207
timestamp 1698175906
transform 1 0 248528 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2271
timestamp 1698175906
transform 1 0 255696 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_2277
timestamp 1698175906
transform 1 0 256368 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2341
timestamp 1698175906
transform 1 0 263536 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_2347
timestamp 1698175906
transform 1 0 264208 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2411
timestamp 1698175906
transform 1 0 271376 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_2417
timestamp 1698175906
transform 1 0 272048 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2481
timestamp 1698175906
transform 1 0 279216 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_2487
timestamp 1698175906
transform 1 0 279888 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2551
timestamp 1698175906
transform 1 0 287056 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_2557
timestamp 1698175906
transform 1 0 287728 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2621
timestamp 1698175906
transform 1 0 294896 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_2627
timestamp 1698175906
transform 1 0 295568 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_2643
timestamp 1698175906
transform 1 0 297360 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_2651
timestamp 1698175906
transform 1 0 298256 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698175906
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698175906
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698175906
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698175906
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698175906
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698175906
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698175906
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698175906
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698175906
transform 1 0 32928 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698175906
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_352
timestamp 1698175906
transform 1 0 40768 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_416
timestamp 1698175906
transform 1 0 47936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698175906
transform 1 0 48608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698175906
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_492
timestamp 1698175906
transform 1 0 56448 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_556
timestamp 1698175906
transform 1 0 63616 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_562
timestamp 1698175906
transform 1 0 64288 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_626
timestamp 1698175906
transform 1 0 71456 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_632
timestamp 1698175906
transform 1 0 72128 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_696
timestamp 1698175906
transform 1 0 79296 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_702
timestamp 1698175906
transform 1 0 79968 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_766
timestamp 1698175906
transform 1 0 87136 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_772
timestamp 1698175906
transform 1 0 87808 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_836
timestamp 1698175906
transform 1 0 94976 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_842
timestamp 1698175906
transform 1 0 95648 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_906
timestamp 1698175906
transform 1 0 102816 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_912
timestamp 1698175906
transform 1 0 103488 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_976
timestamp 1698175906
transform 1 0 110656 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_982
timestamp 1698175906
transform 1 0 111328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1046
timestamp 1698175906
transform 1 0 118496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1052
timestamp 1698175906
transform 1 0 119168 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1116
timestamp 1698175906
transform 1 0 126336 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1122
timestamp 1698175906
transform 1 0 127008 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1186
timestamp 1698175906
transform 1 0 134176 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1192
timestamp 1698175906
transform 1 0 134848 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1256
timestamp 1698175906
transform 1 0 142016 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1262
timestamp 1698175906
transform 1 0 142688 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1326
timestamp 1698175906
transform 1 0 149856 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1332
timestamp 1698175906
transform 1 0 150528 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1396
timestamp 1698175906
transform 1 0 157696 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1402
timestamp 1698175906
transform 1 0 158368 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1466
timestamp 1698175906
transform 1 0 165536 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1472
timestamp 1698175906
transform 1 0 166208 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1536
timestamp 1698175906
transform 1 0 173376 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1542
timestamp 1698175906
transform 1 0 174048 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1606
timestamp 1698175906
transform 1 0 181216 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1612
timestamp 1698175906
transform 1 0 181888 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1676
timestamp 1698175906
transform 1 0 189056 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1682
timestamp 1698175906
transform 1 0 189728 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1746
timestamp 1698175906
transform 1 0 196896 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1752
timestamp 1698175906
transform 1 0 197568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1816
timestamp 1698175906
transform 1 0 204736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1822
timestamp 1698175906
transform 1 0 205408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1886
timestamp 1698175906
transform 1 0 212576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1892
timestamp 1698175906
transform 1 0 213248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1956
timestamp 1698175906
transform 1 0 220416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1962
timestamp 1698175906
transform 1 0 221088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2026
timestamp 1698175906
transform 1 0 228256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2032
timestamp 1698175906
transform 1 0 228928 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2096
timestamp 1698175906
transform 1 0 236096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2102
timestamp 1698175906
transform 1 0 236768 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2166
timestamp 1698175906
transform 1 0 243936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2172
timestamp 1698175906
transform 1 0 244608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2236
timestamp 1698175906
transform 1 0 251776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2242
timestamp 1698175906
transform 1 0 252448 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2306
timestamp 1698175906
transform 1 0 259616 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2312
timestamp 1698175906
transform 1 0 260288 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2376
timestamp 1698175906
transform 1 0 267456 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2382
timestamp 1698175906
transform 1 0 268128 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2446
timestamp 1698175906
transform 1 0 275296 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2452
timestamp 1698175906
transform 1 0 275968 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2516
timestamp 1698175906
transform 1 0 283136 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2522
timestamp 1698175906
transform 1 0 283808 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2586
timestamp 1698175906
transform 1 0 290976 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_2592
timestamp 1698175906
transform 1 0 291648 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_2624
timestamp 1698175906
transform 1 0 295232 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_2640
timestamp 1698175906
transform 1 0 297024 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2648
timestamp 1698175906
transform 1 0 297920 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698175906
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698175906
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698175906
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698175906
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698175906
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698175906
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698175906
transform 1 0 21168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698175906
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698175906
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698175906
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698175906
transform 1 0 36848 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698175906
transform 1 0 44016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_387
timestamp 1698175906
transform 1 0 44688 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_451
timestamp 1698175906
transform 1 0 51856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_457
timestamp 1698175906
transform 1 0 52528 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_521
timestamp 1698175906
transform 1 0 59696 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_527
timestamp 1698175906
transform 1 0 60368 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_591
timestamp 1698175906
transform 1 0 67536 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_597
timestamp 1698175906
transform 1 0 68208 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_661
timestamp 1698175906
transform 1 0 75376 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_667
timestamp 1698175906
transform 1 0 76048 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_731
timestamp 1698175906
transform 1 0 83216 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_737
timestamp 1698175906
transform 1 0 83888 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_801
timestamp 1698175906
transform 1 0 91056 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_807
timestamp 1698175906
transform 1 0 91728 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_871
timestamp 1698175906
transform 1 0 98896 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_877
timestamp 1698175906
transform 1 0 99568 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_941
timestamp 1698175906
transform 1 0 106736 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_947
timestamp 1698175906
transform 1 0 107408 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1011
timestamp 1698175906
transform 1 0 114576 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1017
timestamp 1698175906
transform 1 0 115248 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1081
timestamp 1698175906
transform 1 0 122416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1087
timestamp 1698175906
transform 1 0 123088 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1151
timestamp 1698175906
transform 1 0 130256 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1157
timestamp 1698175906
transform 1 0 130928 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1221
timestamp 1698175906
transform 1 0 138096 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1227
timestamp 1698175906
transform 1 0 138768 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1291
timestamp 1698175906
transform 1 0 145936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1297
timestamp 1698175906
transform 1 0 146608 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1361
timestamp 1698175906
transform 1 0 153776 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1367
timestamp 1698175906
transform 1 0 154448 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1431
timestamp 1698175906
transform 1 0 161616 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1437
timestamp 1698175906
transform 1 0 162288 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1501
timestamp 1698175906
transform 1 0 169456 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1507
timestamp 1698175906
transform 1 0 170128 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1571
timestamp 1698175906
transform 1 0 177296 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1577
timestamp 1698175906
transform 1 0 177968 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1641
timestamp 1698175906
transform 1 0 185136 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1647
timestamp 1698175906
transform 1 0 185808 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1711
timestamp 1698175906
transform 1 0 192976 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1717
timestamp 1698175906
transform 1 0 193648 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1781
timestamp 1698175906
transform 1 0 200816 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1787
timestamp 1698175906
transform 1 0 201488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1851
timestamp 1698175906
transform 1 0 208656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1857
timestamp 1698175906
transform 1 0 209328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1921
timestamp 1698175906
transform 1 0 216496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1927
timestamp 1698175906
transform 1 0 217168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1991
timestamp 1698175906
transform 1 0 224336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1997
timestamp 1698175906
transform 1 0 225008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2061
timestamp 1698175906
transform 1 0 232176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_2067
timestamp 1698175906
transform 1 0 232848 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2131
timestamp 1698175906
transform 1 0 240016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_2137
timestamp 1698175906
transform 1 0 240688 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2201
timestamp 1698175906
transform 1 0 247856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_2207
timestamp 1698175906
transform 1 0 248528 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2271
timestamp 1698175906
transform 1 0 255696 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_2277
timestamp 1698175906
transform 1 0 256368 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2341
timestamp 1698175906
transform 1 0 263536 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_2347
timestamp 1698175906
transform 1 0 264208 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2411
timestamp 1698175906
transform 1 0 271376 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_2417
timestamp 1698175906
transform 1 0 272048 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2481
timestamp 1698175906
transform 1 0 279216 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_2487
timestamp 1698175906
transform 1 0 279888 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2551
timestamp 1698175906
transform 1 0 287056 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_2557
timestamp 1698175906
transform 1 0 287728 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2621
timestamp 1698175906
transform 1 0 294896 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_2627
timestamp 1698175906
transform 1 0 295568 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_2643
timestamp 1698175906
transform 1 0 297360 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_2651
timestamp 1698175906
transform 1 0 298256 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698175906
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698175906
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698175906
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698175906
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698175906
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698175906
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698175906
transform 1 0 25088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698175906
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_282
timestamp 1698175906
transform 1 0 32928 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698175906
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698175906
transform 1 0 40768 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698175906
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_422
timestamp 1698175906
transform 1 0 48608 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698175906
transform 1 0 55776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_492
timestamp 1698175906
transform 1 0 56448 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_556
timestamp 1698175906
transform 1 0 63616 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_562
timestamp 1698175906
transform 1 0 64288 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_626
timestamp 1698175906
transform 1 0 71456 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_632
timestamp 1698175906
transform 1 0 72128 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_696
timestamp 1698175906
transform 1 0 79296 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_702
timestamp 1698175906
transform 1 0 79968 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_766
timestamp 1698175906
transform 1 0 87136 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_772
timestamp 1698175906
transform 1 0 87808 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_836
timestamp 1698175906
transform 1 0 94976 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_842
timestamp 1698175906
transform 1 0 95648 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_906
timestamp 1698175906
transform 1 0 102816 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_912
timestamp 1698175906
transform 1 0 103488 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_976
timestamp 1698175906
transform 1 0 110656 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_982
timestamp 1698175906
transform 1 0 111328 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1046
timestamp 1698175906
transform 1 0 118496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1052
timestamp 1698175906
transform 1 0 119168 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1116
timestamp 1698175906
transform 1 0 126336 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1122
timestamp 1698175906
transform 1 0 127008 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1186
timestamp 1698175906
transform 1 0 134176 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1192
timestamp 1698175906
transform 1 0 134848 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1256
timestamp 1698175906
transform 1 0 142016 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1262
timestamp 1698175906
transform 1 0 142688 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1326
timestamp 1698175906
transform 1 0 149856 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1332
timestamp 1698175906
transform 1 0 150528 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1396
timestamp 1698175906
transform 1 0 157696 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1402
timestamp 1698175906
transform 1 0 158368 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1466
timestamp 1698175906
transform 1 0 165536 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1472
timestamp 1698175906
transform 1 0 166208 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1536
timestamp 1698175906
transform 1 0 173376 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1542
timestamp 1698175906
transform 1 0 174048 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1606
timestamp 1698175906
transform 1 0 181216 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1612
timestamp 1698175906
transform 1 0 181888 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1676
timestamp 1698175906
transform 1 0 189056 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1682
timestamp 1698175906
transform 1 0 189728 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1746
timestamp 1698175906
transform 1 0 196896 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1752
timestamp 1698175906
transform 1 0 197568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1816
timestamp 1698175906
transform 1 0 204736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1822
timestamp 1698175906
transform 1 0 205408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1886
timestamp 1698175906
transform 1 0 212576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1892
timestamp 1698175906
transform 1 0 213248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1956
timestamp 1698175906
transform 1 0 220416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1962
timestamp 1698175906
transform 1 0 221088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2026
timestamp 1698175906
transform 1 0 228256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2032
timestamp 1698175906
transform 1 0 228928 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2096
timestamp 1698175906
transform 1 0 236096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2102
timestamp 1698175906
transform 1 0 236768 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2166
timestamp 1698175906
transform 1 0 243936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2172
timestamp 1698175906
transform 1 0 244608 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2236
timestamp 1698175906
transform 1 0 251776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2242
timestamp 1698175906
transform 1 0 252448 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2306
timestamp 1698175906
transform 1 0 259616 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2312
timestamp 1698175906
transform 1 0 260288 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2376
timestamp 1698175906
transform 1 0 267456 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2382
timestamp 1698175906
transform 1 0 268128 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2446
timestamp 1698175906
transform 1 0 275296 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2452
timestamp 1698175906
transform 1 0 275968 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2516
timestamp 1698175906
transform 1 0 283136 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2522
timestamp 1698175906
transform 1 0 283808 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2586
timestamp 1698175906
transform 1 0 290976 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_2592
timestamp 1698175906
transform 1 0 291648 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_2624
timestamp 1698175906
transform 1 0 295232 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_2640
timestamp 1698175906
transform 1 0 297024 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2648
timestamp 1698175906
transform 1 0 297920 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698175906
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698175906
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698175906
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698175906
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698175906
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698175906
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698175906
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698175906
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698175906
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698175906
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698175906
transform 1 0 36848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698175906
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_387
timestamp 1698175906
transform 1 0 44688 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698175906
transform 1 0 51856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_457
timestamp 1698175906
transform 1 0 52528 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_521
timestamp 1698175906
transform 1 0 59696 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_527
timestamp 1698175906
transform 1 0 60368 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_591
timestamp 1698175906
transform 1 0 67536 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_597
timestamp 1698175906
transform 1 0 68208 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_661
timestamp 1698175906
transform 1 0 75376 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_667
timestamp 1698175906
transform 1 0 76048 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_731
timestamp 1698175906
transform 1 0 83216 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_737
timestamp 1698175906
transform 1 0 83888 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_801
timestamp 1698175906
transform 1 0 91056 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_807
timestamp 1698175906
transform 1 0 91728 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_871
timestamp 1698175906
transform 1 0 98896 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_877
timestamp 1698175906
transform 1 0 99568 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_941
timestamp 1698175906
transform 1 0 106736 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_947
timestamp 1698175906
transform 1 0 107408 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1011
timestamp 1698175906
transform 1 0 114576 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1017
timestamp 1698175906
transform 1 0 115248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1081
timestamp 1698175906
transform 1 0 122416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1087
timestamp 1698175906
transform 1 0 123088 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1151
timestamp 1698175906
transform 1 0 130256 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1157
timestamp 1698175906
transform 1 0 130928 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1221
timestamp 1698175906
transform 1 0 138096 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1227
timestamp 1698175906
transform 1 0 138768 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1291
timestamp 1698175906
transform 1 0 145936 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1297
timestamp 1698175906
transform 1 0 146608 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1361
timestamp 1698175906
transform 1 0 153776 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1367
timestamp 1698175906
transform 1 0 154448 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1431
timestamp 1698175906
transform 1 0 161616 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1437
timestamp 1698175906
transform 1 0 162288 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1501
timestamp 1698175906
transform 1 0 169456 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1507
timestamp 1698175906
transform 1 0 170128 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1571
timestamp 1698175906
transform 1 0 177296 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1577
timestamp 1698175906
transform 1 0 177968 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1641
timestamp 1698175906
transform 1 0 185136 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1647
timestamp 1698175906
transform 1 0 185808 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1711
timestamp 1698175906
transform 1 0 192976 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1717
timestamp 1698175906
transform 1 0 193648 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1781
timestamp 1698175906
transform 1 0 200816 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1787
timestamp 1698175906
transform 1 0 201488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1851
timestamp 1698175906
transform 1 0 208656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1857
timestamp 1698175906
transform 1 0 209328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1921
timestamp 1698175906
transform 1 0 216496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1927
timestamp 1698175906
transform 1 0 217168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1991
timestamp 1698175906
transform 1 0 224336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1997
timestamp 1698175906
transform 1 0 225008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_2061
timestamp 1698175906
transform 1 0 232176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_2067
timestamp 1698175906
transform 1 0 232848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_2131
timestamp 1698175906
transform 1 0 240016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_2137
timestamp 1698175906
transform 1 0 240688 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_2201
timestamp 1698175906
transform 1 0 247856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_2207
timestamp 1698175906
transform 1 0 248528 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_2271
timestamp 1698175906
transform 1 0 255696 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_2277
timestamp 1698175906
transform 1 0 256368 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_2341
timestamp 1698175906
transform 1 0 263536 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_2347
timestamp 1698175906
transform 1 0 264208 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_2411
timestamp 1698175906
transform 1 0 271376 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_2417
timestamp 1698175906
transform 1 0 272048 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_2481
timestamp 1698175906
transform 1 0 279216 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_2487
timestamp 1698175906
transform 1 0 279888 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_2551
timestamp 1698175906
transform 1 0 287056 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_2557
timestamp 1698175906
transform 1 0 287728 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_2621
timestamp 1698175906
transform 1 0 294896 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_2627
timestamp 1698175906
transform 1 0 295568 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_2643
timestamp 1698175906
transform 1 0 297360 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_2651
timestamp 1698175906
transform 1 0 298256 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698175906
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698175906
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698175906
transform 1 0 9408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698175906
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698175906
transform 1 0 17248 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698175906
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698175906
transform 1 0 25088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698175906
transform 1 0 32256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_282
timestamp 1698175906
transform 1 0 32928 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_346
timestamp 1698175906
transform 1 0 40096 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_352
timestamp 1698175906
transform 1 0 40768 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_416
timestamp 1698175906
transform 1 0 47936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_422
timestamp 1698175906
transform 1 0 48608 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_486
timestamp 1698175906
transform 1 0 55776 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_492
timestamp 1698175906
transform 1 0 56448 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_556
timestamp 1698175906
transform 1 0 63616 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_562
timestamp 1698175906
transform 1 0 64288 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_626
timestamp 1698175906
transform 1 0 71456 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_632
timestamp 1698175906
transform 1 0 72128 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_696
timestamp 1698175906
transform 1 0 79296 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_702
timestamp 1698175906
transform 1 0 79968 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_766
timestamp 1698175906
transform 1 0 87136 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_772
timestamp 1698175906
transform 1 0 87808 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_836
timestamp 1698175906
transform 1 0 94976 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_842
timestamp 1698175906
transform 1 0 95648 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_906
timestamp 1698175906
transform 1 0 102816 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_912
timestamp 1698175906
transform 1 0 103488 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_976
timestamp 1698175906
transform 1 0 110656 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_982
timestamp 1698175906
transform 1 0 111328 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1046
timestamp 1698175906
transform 1 0 118496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1052
timestamp 1698175906
transform 1 0 119168 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1116
timestamp 1698175906
transform 1 0 126336 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1122
timestamp 1698175906
transform 1 0 127008 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1186
timestamp 1698175906
transform 1 0 134176 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1192
timestamp 1698175906
transform 1 0 134848 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1256
timestamp 1698175906
transform 1 0 142016 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1262
timestamp 1698175906
transform 1 0 142688 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1326
timestamp 1698175906
transform 1 0 149856 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1332
timestamp 1698175906
transform 1 0 150528 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1396
timestamp 1698175906
transform 1 0 157696 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1402
timestamp 1698175906
transform 1 0 158368 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1466
timestamp 1698175906
transform 1 0 165536 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1472
timestamp 1698175906
transform 1 0 166208 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1536
timestamp 1698175906
transform 1 0 173376 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1542
timestamp 1698175906
transform 1 0 174048 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1606
timestamp 1698175906
transform 1 0 181216 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1612
timestamp 1698175906
transform 1 0 181888 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1676
timestamp 1698175906
transform 1 0 189056 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1682
timestamp 1698175906
transform 1 0 189728 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1746
timestamp 1698175906
transform 1 0 196896 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1752
timestamp 1698175906
transform 1 0 197568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1816
timestamp 1698175906
transform 1 0 204736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1822
timestamp 1698175906
transform 1 0 205408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1886
timestamp 1698175906
transform 1 0 212576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1892
timestamp 1698175906
transform 1 0 213248 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1956
timestamp 1698175906
transform 1 0 220416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1962
timestamp 1698175906
transform 1 0 221088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2026
timestamp 1698175906
transform 1 0 228256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2032
timestamp 1698175906
transform 1 0 228928 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2096
timestamp 1698175906
transform 1 0 236096 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2102
timestamp 1698175906
transform 1 0 236768 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2166
timestamp 1698175906
transform 1 0 243936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2172
timestamp 1698175906
transform 1 0 244608 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2236
timestamp 1698175906
transform 1 0 251776 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2242
timestamp 1698175906
transform 1 0 252448 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2306
timestamp 1698175906
transform 1 0 259616 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2312
timestamp 1698175906
transform 1 0 260288 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2376
timestamp 1698175906
transform 1 0 267456 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2382
timestamp 1698175906
transform 1 0 268128 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2446
timestamp 1698175906
transform 1 0 275296 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2452
timestamp 1698175906
transform 1 0 275968 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2516
timestamp 1698175906
transform 1 0 283136 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2522
timestamp 1698175906
transform 1 0 283808 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2586
timestamp 1698175906
transform 1 0 290976 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2592
timestamp 1698175906
transform 1 0 291648 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_2624
timestamp 1698175906
transform 1 0 295232 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_2640
timestamp 1698175906
transform 1 0 297024 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2648
timestamp 1698175906
transform 1 0 297920 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698175906
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698175906
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698175906
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698175906
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698175906
transform 1 0 13328 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698175906
transform 1 0 20496 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698175906
transform 1 0 21168 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698175906
transform 1 0 28336 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698175906
transform 1 0 29008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698175906
transform 1 0 36176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698175906
transform 1 0 36848 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698175906
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_387
timestamp 1698175906
transform 1 0 44688 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698175906
transform 1 0 51856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_457
timestamp 1698175906
transform 1 0 52528 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_521
timestamp 1698175906
transform 1 0 59696 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_527
timestamp 1698175906
transform 1 0 60368 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_591
timestamp 1698175906
transform 1 0 67536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_597
timestamp 1698175906
transform 1 0 68208 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_661
timestamp 1698175906
transform 1 0 75376 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_667
timestamp 1698175906
transform 1 0 76048 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_731
timestamp 1698175906
transform 1 0 83216 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_737
timestamp 1698175906
transform 1 0 83888 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_801
timestamp 1698175906
transform 1 0 91056 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_807
timestamp 1698175906
transform 1 0 91728 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_871
timestamp 1698175906
transform 1 0 98896 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_877
timestamp 1698175906
transform 1 0 99568 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_941
timestamp 1698175906
transform 1 0 106736 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_947
timestamp 1698175906
transform 1 0 107408 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1011
timestamp 1698175906
transform 1 0 114576 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1017
timestamp 1698175906
transform 1 0 115248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1081
timestamp 1698175906
transform 1 0 122416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1087
timestamp 1698175906
transform 1 0 123088 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1151
timestamp 1698175906
transform 1 0 130256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1157
timestamp 1698175906
transform 1 0 130928 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1221
timestamp 1698175906
transform 1 0 138096 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1227
timestamp 1698175906
transform 1 0 138768 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1291
timestamp 1698175906
transform 1 0 145936 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1297
timestamp 1698175906
transform 1 0 146608 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1361
timestamp 1698175906
transform 1 0 153776 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1367
timestamp 1698175906
transform 1 0 154448 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1431
timestamp 1698175906
transform 1 0 161616 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1437
timestamp 1698175906
transform 1 0 162288 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1501
timestamp 1698175906
transform 1 0 169456 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1507
timestamp 1698175906
transform 1 0 170128 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1571
timestamp 1698175906
transform 1 0 177296 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1577
timestamp 1698175906
transform 1 0 177968 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1641
timestamp 1698175906
transform 1 0 185136 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1647
timestamp 1698175906
transform 1 0 185808 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1711
timestamp 1698175906
transform 1 0 192976 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1717
timestamp 1698175906
transform 1 0 193648 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1781
timestamp 1698175906
transform 1 0 200816 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1787
timestamp 1698175906
transform 1 0 201488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1851
timestamp 1698175906
transform 1 0 208656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1857
timestamp 1698175906
transform 1 0 209328 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1921
timestamp 1698175906
transform 1 0 216496 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1927
timestamp 1698175906
transform 1 0 217168 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1991
timestamp 1698175906
transform 1 0 224336 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1997
timestamp 1698175906
transform 1 0 225008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_2061
timestamp 1698175906
transform 1 0 232176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_2067
timestamp 1698175906
transform 1 0 232848 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_2131
timestamp 1698175906
transform 1 0 240016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_2137
timestamp 1698175906
transform 1 0 240688 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_2201
timestamp 1698175906
transform 1 0 247856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_2207
timestamp 1698175906
transform 1 0 248528 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_2271
timestamp 1698175906
transform 1 0 255696 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_2277
timestamp 1698175906
transform 1 0 256368 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_2341
timestamp 1698175906
transform 1 0 263536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_2347
timestamp 1698175906
transform 1 0 264208 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_2411
timestamp 1698175906
transform 1 0 271376 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_2417
timestamp 1698175906
transform 1 0 272048 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_2481
timestamp 1698175906
transform 1 0 279216 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_2487
timestamp 1698175906
transform 1 0 279888 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_2551
timestamp 1698175906
transform 1 0 287056 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_2557
timestamp 1698175906
transform 1 0 287728 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_2621
timestamp 1698175906
transform 1 0 294896 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_2627
timestamp 1698175906
transform 1 0 295568 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_2643
timestamp 1698175906
transform 1 0 297360 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_2651
timestamp 1698175906
transform 1 0 298256 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2
timestamp 1698175906
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698175906
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1698175906
transform 1 0 9408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698175906
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_142
timestamp 1698175906
transform 1 0 17248 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698175906
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_212
timestamp 1698175906
transform 1 0 25088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_276
timestamp 1698175906
transform 1 0 32256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_282
timestamp 1698175906
transform 1 0 32928 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_346
timestamp 1698175906
transform 1 0 40096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_352
timestamp 1698175906
transform 1 0 40768 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_416
timestamp 1698175906
transform 1 0 47936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_422
timestamp 1698175906
transform 1 0 48608 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_486
timestamp 1698175906
transform 1 0 55776 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_492
timestamp 1698175906
transform 1 0 56448 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_556
timestamp 1698175906
transform 1 0 63616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_562
timestamp 1698175906
transform 1 0 64288 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_626
timestamp 1698175906
transform 1 0 71456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_632
timestamp 1698175906
transform 1 0 72128 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_696
timestamp 1698175906
transform 1 0 79296 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_702
timestamp 1698175906
transform 1 0 79968 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_766
timestamp 1698175906
transform 1 0 87136 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_772
timestamp 1698175906
transform 1 0 87808 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_836
timestamp 1698175906
transform 1 0 94976 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_842
timestamp 1698175906
transform 1 0 95648 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_906
timestamp 1698175906
transform 1 0 102816 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_912
timestamp 1698175906
transform 1 0 103488 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_976
timestamp 1698175906
transform 1 0 110656 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_982
timestamp 1698175906
transform 1 0 111328 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1046
timestamp 1698175906
transform 1 0 118496 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1052
timestamp 1698175906
transform 1 0 119168 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1116
timestamp 1698175906
transform 1 0 126336 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1122
timestamp 1698175906
transform 1 0 127008 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1186
timestamp 1698175906
transform 1 0 134176 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1192
timestamp 1698175906
transform 1 0 134848 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1256
timestamp 1698175906
transform 1 0 142016 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1262
timestamp 1698175906
transform 1 0 142688 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1326
timestamp 1698175906
transform 1 0 149856 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1332
timestamp 1698175906
transform 1 0 150528 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1396
timestamp 1698175906
transform 1 0 157696 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1402
timestamp 1698175906
transform 1 0 158368 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1466
timestamp 1698175906
transform 1 0 165536 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1472
timestamp 1698175906
transform 1 0 166208 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1536
timestamp 1698175906
transform 1 0 173376 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1542
timestamp 1698175906
transform 1 0 174048 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1606
timestamp 1698175906
transform 1 0 181216 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1612
timestamp 1698175906
transform 1 0 181888 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1676
timestamp 1698175906
transform 1 0 189056 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1682
timestamp 1698175906
transform 1 0 189728 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1746
timestamp 1698175906
transform 1 0 196896 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1752
timestamp 1698175906
transform 1 0 197568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1816
timestamp 1698175906
transform 1 0 204736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1822
timestamp 1698175906
transform 1 0 205408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1886
timestamp 1698175906
transform 1 0 212576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1892
timestamp 1698175906
transform 1 0 213248 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1956
timestamp 1698175906
transform 1 0 220416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1962
timestamp 1698175906
transform 1 0 221088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2026
timestamp 1698175906
transform 1 0 228256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2032
timestamp 1698175906
transform 1 0 228928 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2096
timestamp 1698175906
transform 1 0 236096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2102
timestamp 1698175906
transform 1 0 236768 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2166
timestamp 1698175906
transform 1 0 243936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2172
timestamp 1698175906
transform 1 0 244608 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2236
timestamp 1698175906
transform 1 0 251776 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2242
timestamp 1698175906
transform 1 0 252448 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2306
timestamp 1698175906
transform 1 0 259616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2312
timestamp 1698175906
transform 1 0 260288 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2376
timestamp 1698175906
transform 1 0 267456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2382
timestamp 1698175906
transform 1 0 268128 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2446
timestamp 1698175906
transform 1 0 275296 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2452
timestamp 1698175906
transform 1 0 275968 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2516
timestamp 1698175906
transform 1 0 283136 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2522
timestamp 1698175906
transform 1 0 283808 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2586
timestamp 1698175906
transform 1 0 290976 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_2592
timestamp 1698175906
transform 1 0 291648 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_2624
timestamp 1698175906
transform 1 0 295232 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_2640
timestamp 1698175906
transform 1 0 297024 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2648
timestamp 1698175906
transform 1 0 297920 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698175906
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698175906
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698175906
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698175906
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_107
timestamp 1698175906
transform 1 0 13328 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_171
timestamp 1698175906
transform 1 0 20496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_177
timestamp 1698175906
transform 1 0 21168 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698175906
transform 1 0 28336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_247
timestamp 1698175906
transform 1 0 29008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_311
timestamp 1698175906
transform 1 0 36176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_317
timestamp 1698175906
transform 1 0 36848 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_381
timestamp 1698175906
transform 1 0 44016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_387
timestamp 1698175906
transform 1 0 44688 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_451
timestamp 1698175906
transform 1 0 51856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_457
timestamp 1698175906
transform 1 0 52528 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_521
timestamp 1698175906
transform 1 0 59696 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_527
timestamp 1698175906
transform 1 0 60368 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_591
timestamp 1698175906
transform 1 0 67536 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_597
timestamp 1698175906
transform 1 0 68208 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_661
timestamp 1698175906
transform 1 0 75376 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_667
timestamp 1698175906
transform 1 0 76048 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_731
timestamp 1698175906
transform 1 0 83216 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_737
timestamp 1698175906
transform 1 0 83888 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_801
timestamp 1698175906
transform 1 0 91056 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_807
timestamp 1698175906
transform 1 0 91728 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_871
timestamp 1698175906
transform 1 0 98896 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_877
timestamp 1698175906
transform 1 0 99568 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_941
timestamp 1698175906
transform 1 0 106736 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_947
timestamp 1698175906
transform 1 0 107408 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1011
timestamp 1698175906
transform 1 0 114576 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1017
timestamp 1698175906
transform 1 0 115248 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1081
timestamp 1698175906
transform 1 0 122416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1087
timestamp 1698175906
transform 1 0 123088 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1151
timestamp 1698175906
transform 1 0 130256 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1157
timestamp 1698175906
transform 1 0 130928 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1221
timestamp 1698175906
transform 1 0 138096 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1227
timestamp 1698175906
transform 1 0 138768 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1291
timestamp 1698175906
transform 1 0 145936 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1297
timestamp 1698175906
transform 1 0 146608 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1361
timestamp 1698175906
transform 1 0 153776 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1367
timestamp 1698175906
transform 1 0 154448 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1431
timestamp 1698175906
transform 1 0 161616 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1437
timestamp 1698175906
transform 1 0 162288 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1501
timestamp 1698175906
transform 1 0 169456 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1507
timestamp 1698175906
transform 1 0 170128 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1571
timestamp 1698175906
transform 1 0 177296 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1577
timestamp 1698175906
transform 1 0 177968 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1641
timestamp 1698175906
transform 1 0 185136 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1647
timestamp 1698175906
transform 1 0 185808 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1711
timestamp 1698175906
transform 1 0 192976 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1717
timestamp 1698175906
transform 1 0 193648 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1781
timestamp 1698175906
transform 1 0 200816 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1787
timestamp 1698175906
transform 1 0 201488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1851
timestamp 1698175906
transform 1 0 208656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1857
timestamp 1698175906
transform 1 0 209328 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1921
timestamp 1698175906
transform 1 0 216496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1927
timestamp 1698175906
transform 1 0 217168 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1991
timestamp 1698175906
transform 1 0 224336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1997
timestamp 1698175906
transform 1 0 225008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2061
timestamp 1698175906
transform 1 0 232176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_2067
timestamp 1698175906
transform 1 0 232848 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2131
timestamp 1698175906
transform 1 0 240016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_2137
timestamp 1698175906
transform 1 0 240688 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2201
timestamp 1698175906
transform 1 0 247856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_2207
timestamp 1698175906
transform 1 0 248528 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2271
timestamp 1698175906
transform 1 0 255696 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_2277
timestamp 1698175906
transform 1 0 256368 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2341
timestamp 1698175906
transform 1 0 263536 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_2347
timestamp 1698175906
transform 1 0 264208 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2411
timestamp 1698175906
transform 1 0 271376 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_2417
timestamp 1698175906
transform 1 0 272048 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2481
timestamp 1698175906
transform 1 0 279216 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_2487
timestamp 1698175906
transform 1 0 279888 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2551
timestamp 1698175906
transform 1 0 287056 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_2557
timestamp 1698175906
transform 1 0 287728 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2621
timestamp 1698175906
transform 1 0 294896 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_2627
timestamp 1698175906
transform 1 0 295568 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_2643
timestamp 1698175906
transform 1 0 297360 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_2651
timestamp 1698175906
transform 1 0 298256 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698175906
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698175906
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1698175906
transform 1 0 9408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698175906
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_142
timestamp 1698175906
transform 1 0 17248 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698175906
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_212
timestamp 1698175906
transform 1 0 25088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_276
timestamp 1698175906
transform 1 0 32256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_282
timestamp 1698175906
transform 1 0 32928 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_346
timestamp 1698175906
transform 1 0 40096 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_352
timestamp 1698175906
transform 1 0 40768 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_416
timestamp 1698175906
transform 1 0 47936 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_422
timestamp 1698175906
transform 1 0 48608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_486
timestamp 1698175906
transform 1 0 55776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_492
timestamp 1698175906
transform 1 0 56448 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_556
timestamp 1698175906
transform 1 0 63616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_562
timestamp 1698175906
transform 1 0 64288 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_626
timestamp 1698175906
transform 1 0 71456 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_632
timestamp 1698175906
transform 1 0 72128 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_696
timestamp 1698175906
transform 1 0 79296 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_702
timestamp 1698175906
transform 1 0 79968 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_766
timestamp 1698175906
transform 1 0 87136 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_772
timestamp 1698175906
transform 1 0 87808 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_836
timestamp 1698175906
transform 1 0 94976 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_842
timestamp 1698175906
transform 1 0 95648 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_906
timestamp 1698175906
transform 1 0 102816 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_912
timestamp 1698175906
transform 1 0 103488 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_976
timestamp 1698175906
transform 1 0 110656 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_982
timestamp 1698175906
transform 1 0 111328 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1046
timestamp 1698175906
transform 1 0 118496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1052
timestamp 1698175906
transform 1 0 119168 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1116
timestamp 1698175906
transform 1 0 126336 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1122
timestamp 1698175906
transform 1 0 127008 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1186
timestamp 1698175906
transform 1 0 134176 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1192
timestamp 1698175906
transform 1 0 134848 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1256
timestamp 1698175906
transform 1 0 142016 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1262
timestamp 1698175906
transform 1 0 142688 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1326
timestamp 1698175906
transform 1 0 149856 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1332
timestamp 1698175906
transform 1 0 150528 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1396
timestamp 1698175906
transform 1 0 157696 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1402
timestamp 1698175906
transform 1 0 158368 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1466
timestamp 1698175906
transform 1 0 165536 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1472
timestamp 1698175906
transform 1 0 166208 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1536
timestamp 1698175906
transform 1 0 173376 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1542
timestamp 1698175906
transform 1 0 174048 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1606
timestamp 1698175906
transform 1 0 181216 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1612
timestamp 1698175906
transform 1 0 181888 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1676
timestamp 1698175906
transform 1 0 189056 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1682
timestamp 1698175906
transform 1 0 189728 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1746
timestamp 1698175906
transform 1 0 196896 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1752
timestamp 1698175906
transform 1 0 197568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1816
timestamp 1698175906
transform 1 0 204736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1822
timestamp 1698175906
transform 1 0 205408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1886
timestamp 1698175906
transform 1 0 212576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1892
timestamp 1698175906
transform 1 0 213248 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1956
timestamp 1698175906
transform 1 0 220416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1962
timestamp 1698175906
transform 1 0 221088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2026
timestamp 1698175906
transform 1 0 228256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2032
timestamp 1698175906
transform 1 0 228928 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2096
timestamp 1698175906
transform 1 0 236096 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2102
timestamp 1698175906
transform 1 0 236768 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2166
timestamp 1698175906
transform 1 0 243936 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2172
timestamp 1698175906
transform 1 0 244608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2236
timestamp 1698175906
transform 1 0 251776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2242
timestamp 1698175906
transform 1 0 252448 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2306
timestamp 1698175906
transform 1 0 259616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2312
timestamp 1698175906
transform 1 0 260288 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2376
timestamp 1698175906
transform 1 0 267456 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2382
timestamp 1698175906
transform 1 0 268128 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2446
timestamp 1698175906
transform 1 0 275296 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2452
timestamp 1698175906
transform 1 0 275968 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2516
timestamp 1698175906
transform 1 0 283136 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2522
timestamp 1698175906
transform 1 0 283808 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2586
timestamp 1698175906
transform 1 0 290976 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_2592
timestamp 1698175906
transform 1 0 291648 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_2624
timestamp 1698175906
transform 1 0 295232 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_2640
timestamp 1698175906
transform 1 0 297024 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2648
timestamp 1698175906
transform 1 0 297920 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698175906
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698175906
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_37
timestamp 1698175906
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_101
timestamp 1698175906
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_107
timestamp 1698175906
transform 1 0 13328 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_171
timestamp 1698175906
transform 1 0 20496 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_177
timestamp 1698175906
transform 1 0 21168 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_241
timestamp 1698175906
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_247
timestamp 1698175906
transform 1 0 29008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_311
timestamp 1698175906
transform 1 0 36176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_317
timestamp 1698175906
transform 1 0 36848 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_381
timestamp 1698175906
transform 1 0 44016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_387
timestamp 1698175906
transform 1 0 44688 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698175906
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_457
timestamp 1698175906
transform 1 0 52528 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_521
timestamp 1698175906
transform 1 0 59696 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_527
timestamp 1698175906
transform 1 0 60368 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_591
timestamp 1698175906
transform 1 0 67536 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_597
timestamp 1698175906
transform 1 0 68208 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_661
timestamp 1698175906
transform 1 0 75376 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_667
timestamp 1698175906
transform 1 0 76048 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_731
timestamp 1698175906
transform 1 0 83216 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_737
timestamp 1698175906
transform 1 0 83888 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_801
timestamp 1698175906
transform 1 0 91056 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_807
timestamp 1698175906
transform 1 0 91728 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_871
timestamp 1698175906
transform 1 0 98896 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_877
timestamp 1698175906
transform 1 0 99568 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_941
timestamp 1698175906
transform 1 0 106736 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_947
timestamp 1698175906
transform 1 0 107408 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1011
timestamp 1698175906
transform 1 0 114576 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1017
timestamp 1698175906
transform 1 0 115248 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1081
timestamp 1698175906
transform 1 0 122416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1087
timestamp 1698175906
transform 1 0 123088 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1151
timestamp 1698175906
transform 1 0 130256 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1157
timestamp 1698175906
transform 1 0 130928 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1221
timestamp 1698175906
transform 1 0 138096 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1227
timestamp 1698175906
transform 1 0 138768 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1291
timestamp 1698175906
transform 1 0 145936 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1297
timestamp 1698175906
transform 1 0 146608 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1361
timestamp 1698175906
transform 1 0 153776 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1367
timestamp 1698175906
transform 1 0 154448 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1431
timestamp 1698175906
transform 1 0 161616 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1437
timestamp 1698175906
transform 1 0 162288 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1501
timestamp 1698175906
transform 1 0 169456 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1507
timestamp 1698175906
transform 1 0 170128 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1571
timestamp 1698175906
transform 1 0 177296 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1577
timestamp 1698175906
transform 1 0 177968 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1641
timestamp 1698175906
transform 1 0 185136 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1647
timestamp 1698175906
transform 1 0 185808 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1711
timestamp 1698175906
transform 1 0 192976 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1717
timestamp 1698175906
transform 1 0 193648 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1781
timestamp 1698175906
transform 1 0 200816 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1787
timestamp 1698175906
transform 1 0 201488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1851
timestamp 1698175906
transform 1 0 208656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1857
timestamp 1698175906
transform 1 0 209328 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1921
timestamp 1698175906
transform 1 0 216496 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1927
timestamp 1698175906
transform 1 0 217168 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1991
timestamp 1698175906
transform 1 0 224336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1997
timestamp 1698175906
transform 1 0 225008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2061
timestamp 1698175906
transform 1 0 232176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_2067
timestamp 1698175906
transform 1 0 232848 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2131
timestamp 1698175906
transform 1 0 240016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_2137
timestamp 1698175906
transform 1 0 240688 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2201
timestamp 1698175906
transform 1 0 247856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_2207
timestamp 1698175906
transform 1 0 248528 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2271
timestamp 1698175906
transform 1 0 255696 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_2277
timestamp 1698175906
transform 1 0 256368 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2341
timestamp 1698175906
transform 1 0 263536 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_2347
timestamp 1698175906
transform 1 0 264208 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2411
timestamp 1698175906
transform 1 0 271376 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_2417
timestamp 1698175906
transform 1 0 272048 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2481
timestamp 1698175906
transform 1 0 279216 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_2487
timestamp 1698175906
transform 1 0 279888 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2551
timestamp 1698175906
transform 1 0 287056 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_2557
timestamp 1698175906
transform 1 0 287728 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2621
timestamp 1698175906
transform 1 0 294896 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_2627
timestamp 1698175906
transform 1 0 295568 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_2643
timestamp 1698175906
transform 1 0 297360 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_2651
timestamp 1698175906
transform 1 0 298256 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2
timestamp 1698175906
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_66
timestamp 1698175906
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_72
timestamp 1698175906
transform 1 0 9408 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_136
timestamp 1698175906
transform 1 0 16576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_142
timestamp 1698175906
transform 1 0 17248 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_206
timestamp 1698175906
transform 1 0 24416 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_212
timestamp 1698175906
transform 1 0 25088 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_276
timestamp 1698175906
transform 1 0 32256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_282
timestamp 1698175906
transform 1 0 32928 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_346
timestamp 1698175906
transform 1 0 40096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_352
timestamp 1698175906
transform 1 0 40768 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_416
timestamp 1698175906
transform 1 0 47936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_422
timestamp 1698175906
transform 1 0 48608 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_486
timestamp 1698175906
transform 1 0 55776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_492
timestamp 1698175906
transform 1 0 56448 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_556
timestamp 1698175906
transform 1 0 63616 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_562
timestamp 1698175906
transform 1 0 64288 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_626
timestamp 1698175906
transform 1 0 71456 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_632
timestamp 1698175906
transform 1 0 72128 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_696
timestamp 1698175906
transform 1 0 79296 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_702
timestamp 1698175906
transform 1 0 79968 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_766
timestamp 1698175906
transform 1 0 87136 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_772
timestamp 1698175906
transform 1 0 87808 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_836
timestamp 1698175906
transform 1 0 94976 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_842
timestamp 1698175906
transform 1 0 95648 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_906
timestamp 1698175906
transform 1 0 102816 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_912
timestamp 1698175906
transform 1 0 103488 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_976
timestamp 1698175906
transform 1 0 110656 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_982
timestamp 1698175906
transform 1 0 111328 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1046
timestamp 1698175906
transform 1 0 118496 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1052
timestamp 1698175906
transform 1 0 119168 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1116
timestamp 1698175906
transform 1 0 126336 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1122
timestamp 1698175906
transform 1 0 127008 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1186
timestamp 1698175906
transform 1 0 134176 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1192
timestamp 1698175906
transform 1 0 134848 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1256
timestamp 1698175906
transform 1 0 142016 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1262
timestamp 1698175906
transform 1 0 142688 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1326
timestamp 1698175906
transform 1 0 149856 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1332
timestamp 1698175906
transform 1 0 150528 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1396
timestamp 1698175906
transform 1 0 157696 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1402
timestamp 1698175906
transform 1 0 158368 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1466
timestamp 1698175906
transform 1 0 165536 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1472
timestamp 1698175906
transform 1 0 166208 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1536
timestamp 1698175906
transform 1 0 173376 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1542
timestamp 1698175906
transform 1 0 174048 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1606
timestamp 1698175906
transform 1 0 181216 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1612
timestamp 1698175906
transform 1 0 181888 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1676
timestamp 1698175906
transform 1 0 189056 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1682
timestamp 1698175906
transform 1 0 189728 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1746
timestamp 1698175906
transform 1 0 196896 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1752
timestamp 1698175906
transform 1 0 197568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1816
timestamp 1698175906
transform 1 0 204736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1822
timestamp 1698175906
transform 1 0 205408 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1886
timestamp 1698175906
transform 1 0 212576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1892
timestamp 1698175906
transform 1 0 213248 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1956
timestamp 1698175906
transform 1 0 220416 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1962
timestamp 1698175906
transform 1 0 221088 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2026
timestamp 1698175906
transform 1 0 228256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2032
timestamp 1698175906
transform 1 0 228928 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2096
timestamp 1698175906
transform 1 0 236096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2102
timestamp 1698175906
transform 1 0 236768 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2166
timestamp 1698175906
transform 1 0 243936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2172
timestamp 1698175906
transform 1 0 244608 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2236
timestamp 1698175906
transform 1 0 251776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2242
timestamp 1698175906
transform 1 0 252448 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2306
timestamp 1698175906
transform 1 0 259616 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2312
timestamp 1698175906
transform 1 0 260288 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2376
timestamp 1698175906
transform 1 0 267456 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2382
timestamp 1698175906
transform 1 0 268128 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2446
timestamp 1698175906
transform 1 0 275296 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2452
timestamp 1698175906
transform 1 0 275968 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2516
timestamp 1698175906
transform 1 0 283136 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2522
timestamp 1698175906
transform 1 0 283808 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2586
timestamp 1698175906
transform 1 0 290976 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_2592
timestamp 1698175906
transform 1 0 291648 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_2624
timestamp 1698175906
transform 1 0 295232 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_2640
timestamp 1698175906
transform 1 0 297024 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2648
timestamp 1698175906
transform 1 0 297920 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698175906
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698175906
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_37
timestamp 1698175906
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_101
timestamp 1698175906
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_107
timestamp 1698175906
transform 1 0 13328 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698175906
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_177
timestamp 1698175906
transform 1 0 21168 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_241
timestamp 1698175906
transform 1 0 28336 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_247
timestamp 1698175906
transform 1 0 29008 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_311
timestamp 1698175906
transform 1 0 36176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_317
timestamp 1698175906
transform 1 0 36848 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_381
timestamp 1698175906
transform 1 0 44016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_387
timestamp 1698175906
transform 1 0 44688 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_451
timestamp 1698175906
transform 1 0 51856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_457
timestamp 1698175906
transform 1 0 52528 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_521
timestamp 1698175906
transform 1 0 59696 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_527
timestamp 1698175906
transform 1 0 60368 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_591
timestamp 1698175906
transform 1 0 67536 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_597
timestamp 1698175906
transform 1 0 68208 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_661
timestamp 1698175906
transform 1 0 75376 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_667
timestamp 1698175906
transform 1 0 76048 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_731
timestamp 1698175906
transform 1 0 83216 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_737
timestamp 1698175906
transform 1 0 83888 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_801
timestamp 1698175906
transform 1 0 91056 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_807
timestamp 1698175906
transform 1 0 91728 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_871
timestamp 1698175906
transform 1 0 98896 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_877
timestamp 1698175906
transform 1 0 99568 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_941
timestamp 1698175906
transform 1 0 106736 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_947
timestamp 1698175906
transform 1 0 107408 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1011
timestamp 1698175906
transform 1 0 114576 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1017
timestamp 1698175906
transform 1 0 115248 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1081
timestamp 1698175906
transform 1 0 122416 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1087
timestamp 1698175906
transform 1 0 123088 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1151
timestamp 1698175906
transform 1 0 130256 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1157
timestamp 1698175906
transform 1 0 130928 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1221
timestamp 1698175906
transform 1 0 138096 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1227
timestamp 1698175906
transform 1 0 138768 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1291
timestamp 1698175906
transform 1 0 145936 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1297
timestamp 1698175906
transform 1 0 146608 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1361
timestamp 1698175906
transform 1 0 153776 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1367
timestamp 1698175906
transform 1 0 154448 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1431
timestamp 1698175906
transform 1 0 161616 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1437
timestamp 1698175906
transform 1 0 162288 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1501
timestamp 1698175906
transform 1 0 169456 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1507
timestamp 1698175906
transform 1 0 170128 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1571
timestamp 1698175906
transform 1 0 177296 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1577
timestamp 1698175906
transform 1 0 177968 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1641
timestamp 1698175906
transform 1 0 185136 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1647
timestamp 1698175906
transform 1 0 185808 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1711
timestamp 1698175906
transform 1 0 192976 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1717
timestamp 1698175906
transform 1 0 193648 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1781
timestamp 1698175906
transform 1 0 200816 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1787
timestamp 1698175906
transform 1 0 201488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1851
timestamp 1698175906
transform 1 0 208656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1857
timestamp 1698175906
transform 1 0 209328 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1921
timestamp 1698175906
transform 1 0 216496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1927
timestamp 1698175906
transform 1 0 217168 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1991
timestamp 1698175906
transform 1 0 224336 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1997
timestamp 1698175906
transform 1 0 225008 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2061
timestamp 1698175906
transform 1 0 232176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_2067
timestamp 1698175906
transform 1 0 232848 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2131
timestamp 1698175906
transform 1 0 240016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_2137
timestamp 1698175906
transform 1 0 240688 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2201
timestamp 1698175906
transform 1 0 247856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_2207
timestamp 1698175906
transform 1 0 248528 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2271
timestamp 1698175906
transform 1 0 255696 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_2277
timestamp 1698175906
transform 1 0 256368 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2341
timestamp 1698175906
transform 1 0 263536 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_2347
timestamp 1698175906
transform 1 0 264208 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2411
timestamp 1698175906
transform 1 0 271376 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_2417
timestamp 1698175906
transform 1 0 272048 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2481
timestamp 1698175906
transform 1 0 279216 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_2487
timestamp 1698175906
transform 1 0 279888 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2551
timestamp 1698175906
transform 1 0 287056 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_2557
timestamp 1698175906
transform 1 0 287728 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2621
timestamp 1698175906
transform 1 0 294896 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_2627
timestamp 1698175906
transform 1 0 295568 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_2643
timestamp 1698175906
transform 1 0 297360 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_2651
timestamp 1698175906
transform 1 0 298256 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2
timestamp 1698175906
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_66
timestamp 1698175906
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_72
timestamp 1698175906
transform 1 0 9408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698175906
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_142
timestamp 1698175906
transform 1 0 17248 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_206
timestamp 1698175906
transform 1 0 24416 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_212
timestamp 1698175906
transform 1 0 25088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_276
timestamp 1698175906
transform 1 0 32256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_282
timestamp 1698175906
transform 1 0 32928 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_346
timestamp 1698175906
transform 1 0 40096 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_352
timestamp 1698175906
transform 1 0 40768 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_416
timestamp 1698175906
transform 1 0 47936 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_422
timestamp 1698175906
transform 1 0 48608 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_486
timestamp 1698175906
transform 1 0 55776 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_492
timestamp 1698175906
transform 1 0 56448 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_556
timestamp 1698175906
transform 1 0 63616 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_562
timestamp 1698175906
transform 1 0 64288 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_626
timestamp 1698175906
transform 1 0 71456 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_632
timestamp 1698175906
transform 1 0 72128 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_696
timestamp 1698175906
transform 1 0 79296 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_702
timestamp 1698175906
transform 1 0 79968 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_766
timestamp 1698175906
transform 1 0 87136 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_772
timestamp 1698175906
transform 1 0 87808 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_836
timestamp 1698175906
transform 1 0 94976 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_842
timestamp 1698175906
transform 1 0 95648 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_906
timestamp 1698175906
transform 1 0 102816 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_912
timestamp 1698175906
transform 1 0 103488 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_976
timestamp 1698175906
transform 1 0 110656 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_982
timestamp 1698175906
transform 1 0 111328 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1046
timestamp 1698175906
transform 1 0 118496 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1052
timestamp 1698175906
transform 1 0 119168 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1116
timestamp 1698175906
transform 1 0 126336 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1122
timestamp 1698175906
transform 1 0 127008 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1186
timestamp 1698175906
transform 1 0 134176 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1192
timestamp 1698175906
transform 1 0 134848 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1256
timestamp 1698175906
transform 1 0 142016 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1262
timestamp 1698175906
transform 1 0 142688 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1326
timestamp 1698175906
transform 1 0 149856 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1332
timestamp 1698175906
transform 1 0 150528 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1396
timestamp 1698175906
transform 1 0 157696 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1402
timestamp 1698175906
transform 1 0 158368 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1466
timestamp 1698175906
transform 1 0 165536 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1472
timestamp 1698175906
transform 1 0 166208 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1536
timestamp 1698175906
transform 1 0 173376 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1542
timestamp 1698175906
transform 1 0 174048 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1606
timestamp 1698175906
transform 1 0 181216 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1612
timestamp 1698175906
transform 1 0 181888 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1676
timestamp 1698175906
transform 1 0 189056 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1682
timestamp 1698175906
transform 1 0 189728 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1746
timestamp 1698175906
transform 1 0 196896 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1752
timestamp 1698175906
transform 1 0 197568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1816
timestamp 1698175906
transform 1 0 204736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1822
timestamp 1698175906
transform 1 0 205408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1886
timestamp 1698175906
transform 1 0 212576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1892
timestamp 1698175906
transform 1 0 213248 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1956
timestamp 1698175906
transform 1 0 220416 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1962
timestamp 1698175906
transform 1 0 221088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2026
timestamp 1698175906
transform 1 0 228256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2032
timestamp 1698175906
transform 1 0 228928 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2096
timestamp 1698175906
transform 1 0 236096 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2102
timestamp 1698175906
transform 1 0 236768 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2166
timestamp 1698175906
transform 1 0 243936 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2172
timestamp 1698175906
transform 1 0 244608 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2236
timestamp 1698175906
transform 1 0 251776 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2242
timestamp 1698175906
transform 1 0 252448 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2306
timestamp 1698175906
transform 1 0 259616 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2312
timestamp 1698175906
transform 1 0 260288 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2376
timestamp 1698175906
transform 1 0 267456 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2382
timestamp 1698175906
transform 1 0 268128 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2446
timestamp 1698175906
transform 1 0 275296 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2452
timestamp 1698175906
transform 1 0 275968 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2516
timestamp 1698175906
transform 1 0 283136 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2522
timestamp 1698175906
transform 1 0 283808 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2586
timestamp 1698175906
transform 1 0 290976 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_2592
timestamp 1698175906
transform 1 0 291648 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_2624
timestamp 1698175906
transform 1 0 295232 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_2640
timestamp 1698175906
transform 1 0 297024 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2648
timestamp 1698175906
transform 1 0 297920 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698175906
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698175906
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698175906
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698175906
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_107
timestamp 1698175906
transform 1 0 13328 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_171
timestamp 1698175906
transform 1 0 20496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_177
timestamp 1698175906
transform 1 0 21168 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_241
timestamp 1698175906
transform 1 0 28336 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_247
timestamp 1698175906
transform 1 0 29008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_311
timestamp 1698175906
transform 1 0 36176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_317
timestamp 1698175906
transform 1 0 36848 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_381
timestamp 1698175906
transform 1 0 44016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_387
timestamp 1698175906
transform 1 0 44688 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_451
timestamp 1698175906
transform 1 0 51856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_457
timestamp 1698175906
transform 1 0 52528 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_521
timestamp 1698175906
transform 1 0 59696 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_527
timestamp 1698175906
transform 1 0 60368 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_591
timestamp 1698175906
transform 1 0 67536 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_597
timestamp 1698175906
transform 1 0 68208 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_661
timestamp 1698175906
transform 1 0 75376 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_667
timestamp 1698175906
transform 1 0 76048 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_731
timestamp 1698175906
transform 1 0 83216 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_737
timestamp 1698175906
transform 1 0 83888 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_801
timestamp 1698175906
transform 1 0 91056 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_807
timestamp 1698175906
transform 1 0 91728 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_871
timestamp 1698175906
transform 1 0 98896 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_877
timestamp 1698175906
transform 1 0 99568 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_941
timestamp 1698175906
transform 1 0 106736 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_947
timestamp 1698175906
transform 1 0 107408 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1011
timestamp 1698175906
transform 1 0 114576 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1017
timestamp 1698175906
transform 1 0 115248 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1081
timestamp 1698175906
transform 1 0 122416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1087
timestamp 1698175906
transform 1 0 123088 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1151
timestamp 1698175906
transform 1 0 130256 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1157
timestamp 1698175906
transform 1 0 130928 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1221
timestamp 1698175906
transform 1 0 138096 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1227
timestamp 1698175906
transform 1 0 138768 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1291
timestamp 1698175906
transform 1 0 145936 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1297
timestamp 1698175906
transform 1 0 146608 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1361
timestamp 1698175906
transform 1 0 153776 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1367
timestamp 1698175906
transform 1 0 154448 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1431
timestamp 1698175906
transform 1 0 161616 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1437
timestamp 1698175906
transform 1 0 162288 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1501
timestamp 1698175906
transform 1 0 169456 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1507
timestamp 1698175906
transform 1 0 170128 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1571
timestamp 1698175906
transform 1 0 177296 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1577
timestamp 1698175906
transform 1 0 177968 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1641
timestamp 1698175906
transform 1 0 185136 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1647
timestamp 1698175906
transform 1 0 185808 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1711
timestamp 1698175906
transform 1 0 192976 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1717
timestamp 1698175906
transform 1 0 193648 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1781
timestamp 1698175906
transform 1 0 200816 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1787
timestamp 1698175906
transform 1 0 201488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1851
timestamp 1698175906
transform 1 0 208656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1857
timestamp 1698175906
transform 1 0 209328 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1921
timestamp 1698175906
transform 1 0 216496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1927
timestamp 1698175906
transform 1 0 217168 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1991
timestamp 1698175906
transform 1 0 224336 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1997
timestamp 1698175906
transform 1 0 225008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2061
timestamp 1698175906
transform 1 0 232176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_2067
timestamp 1698175906
transform 1 0 232848 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2131
timestamp 1698175906
transform 1 0 240016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_2137
timestamp 1698175906
transform 1 0 240688 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2201
timestamp 1698175906
transform 1 0 247856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_2207
timestamp 1698175906
transform 1 0 248528 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2271
timestamp 1698175906
transform 1 0 255696 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_2277
timestamp 1698175906
transform 1 0 256368 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2341
timestamp 1698175906
transform 1 0 263536 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_2347
timestamp 1698175906
transform 1 0 264208 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2411
timestamp 1698175906
transform 1 0 271376 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_2417
timestamp 1698175906
transform 1 0 272048 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2481
timestamp 1698175906
transform 1 0 279216 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_2487
timestamp 1698175906
transform 1 0 279888 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2551
timestamp 1698175906
transform 1 0 287056 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_2557
timestamp 1698175906
transform 1 0 287728 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2621
timestamp 1698175906
transform 1 0 294896 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_2627
timestamp 1698175906
transform 1 0 295568 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_2643
timestamp 1698175906
transform 1 0 297360 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_2651
timestamp 1698175906
transform 1 0 298256 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2
timestamp 1698175906
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1698175906
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_72
timestamp 1698175906
transform 1 0 9408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698175906
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_142
timestamp 1698175906
transform 1 0 17248 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_206
timestamp 1698175906
transform 1 0 24416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_212
timestamp 1698175906
transform 1 0 25088 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_276
timestamp 1698175906
transform 1 0 32256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_282
timestamp 1698175906
transform 1 0 32928 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_346
timestamp 1698175906
transform 1 0 40096 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_352
timestamp 1698175906
transform 1 0 40768 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_416
timestamp 1698175906
transform 1 0 47936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_422
timestamp 1698175906
transform 1 0 48608 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_486
timestamp 1698175906
transform 1 0 55776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_492
timestamp 1698175906
transform 1 0 56448 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_556
timestamp 1698175906
transform 1 0 63616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_562
timestamp 1698175906
transform 1 0 64288 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_626
timestamp 1698175906
transform 1 0 71456 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_632
timestamp 1698175906
transform 1 0 72128 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_696
timestamp 1698175906
transform 1 0 79296 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_702
timestamp 1698175906
transform 1 0 79968 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_766
timestamp 1698175906
transform 1 0 87136 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_772
timestamp 1698175906
transform 1 0 87808 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_836
timestamp 1698175906
transform 1 0 94976 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_842
timestamp 1698175906
transform 1 0 95648 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_906
timestamp 1698175906
transform 1 0 102816 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_912
timestamp 1698175906
transform 1 0 103488 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_976
timestamp 1698175906
transform 1 0 110656 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_982
timestamp 1698175906
transform 1 0 111328 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1046
timestamp 1698175906
transform 1 0 118496 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1052
timestamp 1698175906
transform 1 0 119168 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1116
timestamp 1698175906
transform 1 0 126336 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1122
timestamp 1698175906
transform 1 0 127008 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1186
timestamp 1698175906
transform 1 0 134176 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1192
timestamp 1698175906
transform 1 0 134848 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1256
timestamp 1698175906
transform 1 0 142016 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1262
timestamp 1698175906
transform 1 0 142688 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1326
timestamp 1698175906
transform 1 0 149856 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1332
timestamp 1698175906
transform 1 0 150528 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1396
timestamp 1698175906
transform 1 0 157696 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1402
timestamp 1698175906
transform 1 0 158368 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1466
timestamp 1698175906
transform 1 0 165536 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1472
timestamp 1698175906
transform 1 0 166208 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1536
timestamp 1698175906
transform 1 0 173376 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1542
timestamp 1698175906
transform 1 0 174048 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1606
timestamp 1698175906
transform 1 0 181216 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1612
timestamp 1698175906
transform 1 0 181888 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1676
timestamp 1698175906
transform 1 0 189056 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1682
timestamp 1698175906
transform 1 0 189728 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1746
timestamp 1698175906
transform 1 0 196896 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1752
timestamp 1698175906
transform 1 0 197568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1816
timestamp 1698175906
transform 1 0 204736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1822
timestamp 1698175906
transform 1 0 205408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1886
timestamp 1698175906
transform 1 0 212576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1892
timestamp 1698175906
transform 1 0 213248 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1956
timestamp 1698175906
transform 1 0 220416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1962
timestamp 1698175906
transform 1 0 221088 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_2026
timestamp 1698175906
transform 1 0 228256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2032
timestamp 1698175906
transform 1 0 228928 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_2096
timestamp 1698175906
transform 1 0 236096 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2102
timestamp 1698175906
transform 1 0 236768 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_2166
timestamp 1698175906
transform 1 0 243936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2172
timestamp 1698175906
transform 1 0 244608 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_2236
timestamp 1698175906
transform 1 0 251776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2242
timestamp 1698175906
transform 1 0 252448 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_2306
timestamp 1698175906
transform 1 0 259616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2312
timestamp 1698175906
transform 1 0 260288 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_2376
timestamp 1698175906
transform 1 0 267456 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2382
timestamp 1698175906
transform 1 0 268128 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_2446
timestamp 1698175906
transform 1 0 275296 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2452
timestamp 1698175906
transform 1 0 275968 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_2516
timestamp 1698175906
transform 1 0 283136 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2522
timestamp 1698175906
transform 1 0 283808 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_2586
timestamp 1698175906
transform 1 0 290976 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_2592
timestamp 1698175906
transform 1 0 291648 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_2624
timestamp 1698175906
transform 1 0 295232 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_2640
timestamp 1698175906
transform 1 0 297024 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_2648
timestamp 1698175906
transform 1 0 297920 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698175906
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698175906
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698175906
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698175906
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_107
timestamp 1698175906
transform 1 0 13328 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_171
timestamp 1698175906
transform 1 0 20496 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_177
timestamp 1698175906
transform 1 0 21168 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_241
timestamp 1698175906
transform 1 0 28336 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_247
timestamp 1698175906
transform 1 0 29008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_311
timestamp 1698175906
transform 1 0 36176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_317
timestamp 1698175906
transform 1 0 36848 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_381
timestamp 1698175906
transform 1 0 44016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_387
timestamp 1698175906
transform 1 0 44688 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_451
timestamp 1698175906
transform 1 0 51856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_457
timestamp 1698175906
transform 1 0 52528 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_521
timestamp 1698175906
transform 1 0 59696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_527
timestamp 1698175906
transform 1 0 60368 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_591
timestamp 1698175906
transform 1 0 67536 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_597
timestamp 1698175906
transform 1 0 68208 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_661
timestamp 1698175906
transform 1 0 75376 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_667
timestamp 1698175906
transform 1 0 76048 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_731
timestamp 1698175906
transform 1 0 83216 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_737
timestamp 1698175906
transform 1 0 83888 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_801
timestamp 1698175906
transform 1 0 91056 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_807
timestamp 1698175906
transform 1 0 91728 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_871
timestamp 1698175906
transform 1 0 98896 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_877
timestamp 1698175906
transform 1 0 99568 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_941
timestamp 1698175906
transform 1 0 106736 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_947
timestamp 1698175906
transform 1 0 107408 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1011
timestamp 1698175906
transform 1 0 114576 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1017
timestamp 1698175906
transform 1 0 115248 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1081
timestamp 1698175906
transform 1 0 122416 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1087
timestamp 1698175906
transform 1 0 123088 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1151
timestamp 1698175906
transform 1 0 130256 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1157
timestamp 1698175906
transform 1 0 130928 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1221
timestamp 1698175906
transform 1 0 138096 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1227
timestamp 1698175906
transform 1 0 138768 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1291
timestamp 1698175906
transform 1 0 145936 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1297
timestamp 1698175906
transform 1 0 146608 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1361
timestamp 1698175906
transform 1 0 153776 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1367
timestamp 1698175906
transform 1 0 154448 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1431
timestamp 1698175906
transform 1 0 161616 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1437
timestamp 1698175906
transform 1 0 162288 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1501
timestamp 1698175906
transform 1 0 169456 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1507
timestamp 1698175906
transform 1 0 170128 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1571
timestamp 1698175906
transform 1 0 177296 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1577
timestamp 1698175906
transform 1 0 177968 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1641
timestamp 1698175906
transform 1 0 185136 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1647
timestamp 1698175906
transform 1 0 185808 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1711
timestamp 1698175906
transform 1 0 192976 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1717
timestamp 1698175906
transform 1 0 193648 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1781
timestamp 1698175906
transform 1 0 200816 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1787
timestamp 1698175906
transform 1 0 201488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1851
timestamp 1698175906
transform 1 0 208656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1857
timestamp 1698175906
transform 1 0 209328 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1921
timestamp 1698175906
transform 1 0 216496 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1927
timestamp 1698175906
transform 1 0 217168 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1991
timestamp 1698175906
transform 1 0 224336 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1997
timestamp 1698175906
transform 1 0 225008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_2061
timestamp 1698175906
transform 1 0 232176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_2067
timestamp 1698175906
transform 1 0 232848 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_2131
timestamp 1698175906
transform 1 0 240016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_2137
timestamp 1698175906
transform 1 0 240688 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_2201
timestamp 1698175906
transform 1 0 247856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_2207
timestamp 1698175906
transform 1 0 248528 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_2271
timestamp 1698175906
transform 1 0 255696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_2277
timestamp 1698175906
transform 1 0 256368 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_2341
timestamp 1698175906
transform 1 0 263536 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_2347
timestamp 1698175906
transform 1 0 264208 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_2411
timestamp 1698175906
transform 1 0 271376 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_2417
timestamp 1698175906
transform 1 0 272048 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_2481
timestamp 1698175906
transform 1 0 279216 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_2487
timestamp 1698175906
transform 1 0 279888 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_2551
timestamp 1698175906
transform 1 0 287056 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_2557
timestamp 1698175906
transform 1 0 287728 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_2621
timestamp 1698175906
transform 1 0 294896 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_2627
timestamp 1698175906
transform 1 0 295568 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_2643
timestamp 1698175906
transform 1 0 297360 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_2651
timestamp 1698175906
transform 1 0 298256 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2
timestamp 1698175906
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1698175906
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_72
timestamp 1698175906
transform 1 0 9408 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_136
timestamp 1698175906
transform 1 0 16576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_142
timestamp 1698175906
transform 1 0 17248 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698175906
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_212
timestamp 1698175906
transform 1 0 25088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_276
timestamp 1698175906
transform 1 0 32256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_282
timestamp 1698175906
transform 1 0 32928 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_346
timestamp 1698175906
transform 1 0 40096 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_352
timestamp 1698175906
transform 1 0 40768 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_416
timestamp 1698175906
transform 1 0 47936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_422
timestamp 1698175906
transform 1 0 48608 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_486
timestamp 1698175906
transform 1 0 55776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_492
timestamp 1698175906
transform 1 0 56448 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_556
timestamp 1698175906
transform 1 0 63616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_562
timestamp 1698175906
transform 1 0 64288 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_626
timestamp 1698175906
transform 1 0 71456 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_632
timestamp 1698175906
transform 1 0 72128 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_696
timestamp 1698175906
transform 1 0 79296 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_702
timestamp 1698175906
transform 1 0 79968 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_766
timestamp 1698175906
transform 1 0 87136 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_772
timestamp 1698175906
transform 1 0 87808 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_836
timestamp 1698175906
transform 1 0 94976 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_842
timestamp 1698175906
transform 1 0 95648 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_906
timestamp 1698175906
transform 1 0 102816 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_912
timestamp 1698175906
transform 1 0 103488 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_976
timestamp 1698175906
transform 1 0 110656 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_982
timestamp 1698175906
transform 1 0 111328 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1046
timestamp 1698175906
transform 1 0 118496 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1052
timestamp 1698175906
transform 1 0 119168 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1116
timestamp 1698175906
transform 1 0 126336 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1122
timestamp 1698175906
transform 1 0 127008 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1186
timestamp 1698175906
transform 1 0 134176 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1192
timestamp 1698175906
transform 1 0 134848 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1256
timestamp 1698175906
transform 1 0 142016 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1262
timestamp 1698175906
transform 1 0 142688 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1326
timestamp 1698175906
transform 1 0 149856 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1332
timestamp 1698175906
transform 1 0 150528 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1396
timestamp 1698175906
transform 1 0 157696 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1402
timestamp 1698175906
transform 1 0 158368 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1466
timestamp 1698175906
transform 1 0 165536 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1472
timestamp 1698175906
transform 1 0 166208 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1536
timestamp 1698175906
transform 1 0 173376 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1542
timestamp 1698175906
transform 1 0 174048 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1606
timestamp 1698175906
transform 1 0 181216 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1612
timestamp 1698175906
transform 1 0 181888 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1676
timestamp 1698175906
transform 1 0 189056 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1682
timestamp 1698175906
transform 1 0 189728 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1746
timestamp 1698175906
transform 1 0 196896 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1752
timestamp 1698175906
transform 1 0 197568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1816
timestamp 1698175906
transform 1 0 204736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1822
timestamp 1698175906
transform 1 0 205408 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1886
timestamp 1698175906
transform 1 0 212576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1892
timestamp 1698175906
transform 1 0 213248 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1956
timestamp 1698175906
transform 1 0 220416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1962
timestamp 1698175906
transform 1 0 221088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2026
timestamp 1698175906
transform 1 0 228256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2032
timestamp 1698175906
transform 1 0 228928 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2096
timestamp 1698175906
transform 1 0 236096 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2102
timestamp 1698175906
transform 1 0 236768 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2166
timestamp 1698175906
transform 1 0 243936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2172
timestamp 1698175906
transform 1 0 244608 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2236
timestamp 1698175906
transform 1 0 251776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2242
timestamp 1698175906
transform 1 0 252448 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2306
timestamp 1698175906
transform 1 0 259616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2312
timestamp 1698175906
transform 1 0 260288 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2376
timestamp 1698175906
transform 1 0 267456 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2382
timestamp 1698175906
transform 1 0 268128 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2446
timestamp 1698175906
transform 1 0 275296 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2452
timestamp 1698175906
transform 1 0 275968 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2516
timestamp 1698175906
transform 1 0 283136 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2522
timestamp 1698175906
transform 1 0 283808 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2586
timestamp 1698175906
transform 1 0 290976 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_2592
timestamp 1698175906
transform 1 0 291648 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_2624
timestamp 1698175906
transform 1 0 295232 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_2640
timestamp 1698175906
transform 1 0 297024 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2648
timestamp 1698175906
transform 1 0 297920 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698175906
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698175906
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698175906
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698175906
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_107
timestamp 1698175906
transform 1 0 13328 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_171
timestamp 1698175906
transform 1 0 20496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_177
timestamp 1698175906
transform 1 0 21168 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_241
timestamp 1698175906
transform 1 0 28336 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_247
timestamp 1698175906
transform 1 0 29008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_311
timestamp 1698175906
transform 1 0 36176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_317
timestamp 1698175906
transform 1 0 36848 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_381
timestamp 1698175906
transform 1 0 44016 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_387
timestamp 1698175906
transform 1 0 44688 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_451
timestamp 1698175906
transform 1 0 51856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_457
timestamp 1698175906
transform 1 0 52528 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_521
timestamp 1698175906
transform 1 0 59696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_527
timestamp 1698175906
transform 1 0 60368 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_591
timestamp 1698175906
transform 1 0 67536 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_597
timestamp 1698175906
transform 1 0 68208 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_661
timestamp 1698175906
transform 1 0 75376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_667
timestamp 1698175906
transform 1 0 76048 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_731
timestamp 1698175906
transform 1 0 83216 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_737
timestamp 1698175906
transform 1 0 83888 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_801
timestamp 1698175906
transform 1 0 91056 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_807
timestamp 1698175906
transform 1 0 91728 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_871
timestamp 1698175906
transform 1 0 98896 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_877
timestamp 1698175906
transform 1 0 99568 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_941
timestamp 1698175906
transform 1 0 106736 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_947
timestamp 1698175906
transform 1 0 107408 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1011
timestamp 1698175906
transform 1 0 114576 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1017
timestamp 1698175906
transform 1 0 115248 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1081
timestamp 1698175906
transform 1 0 122416 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1087
timestamp 1698175906
transform 1 0 123088 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1151
timestamp 1698175906
transform 1 0 130256 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1157
timestamp 1698175906
transform 1 0 130928 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1221
timestamp 1698175906
transform 1 0 138096 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1227
timestamp 1698175906
transform 1 0 138768 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1291
timestamp 1698175906
transform 1 0 145936 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1297
timestamp 1698175906
transform 1 0 146608 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1361
timestamp 1698175906
transform 1 0 153776 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1367
timestamp 1698175906
transform 1 0 154448 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1431
timestamp 1698175906
transform 1 0 161616 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1437
timestamp 1698175906
transform 1 0 162288 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1501
timestamp 1698175906
transform 1 0 169456 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1507
timestamp 1698175906
transform 1 0 170128 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1571
timestamp 1698175906
transform 1 0 177296 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1577
timestamp 1698175906
transform 1 0 177968 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1641
timestamp 1698175906
transform 1 0 185136 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_1647
timestamp 1698175906
transform 1 0 185808 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1651
timestamp 1698175906
transform 1 0 186256 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1717
timestamp 1698175906
transform 1 0 193648 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1781
timestamp 1698175906
transform 1 0 200816 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1787
timestamp 1698175906
transform 1 0 201488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1851
timestamp 1698175906
transform 1 0 208656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1857
timestamp 1698175906
transform 1 0 209328 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1921
timestamp 1698175906
transform 1 0 216496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1927
timestamp 1698175906
transform 1 0 217168 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1991
timestamp 1698175906
transform 1 0 224336 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1997
timestamp 1698175906
transform 1 0 225008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_2061
timestamp 1698175906
transform 1 0 232176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_2067
timestamp 1698175906
transform 1 0 232848 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_2131
timestamp 1698175906
transform 1 0 240016 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_2137
timestamp 1698175906
transform 1 0 240688 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_2201
timestamp 1698175906
transform 1 0 247856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_2207
timestamp 1698175906
transform 1 0 248528 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_2271
timestamp 1698175906
transform 1 0 255696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_2277
timestamp 1698175906
transform 1 0 256368 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_2341
timestamp 1698175906
transform 1 0 263536 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_2347
timestamp 1698175906
transform 1 0 264208 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_2411
timestamp 1698175906
transform 1 0 271376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_2417
timestamp 1698175906
transform 1 0 272048 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_2481
timestamp 1698175906
transform 1 0 279216 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_2487
timestamp 1698175906
transform 1 0 279888 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_2551
timestamp 1698175906
transform 1 0 287056 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_2557
timestamp 1698175906
transform 1 0 287728 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_2621
timestamp 1698175906
transform 1 0 294896 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_2627
timestamp 1698175906
transform 1 0 295568 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_2643
timestamp 1698175906
transform 1 0 297360 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_2651
timestamp 1698175906
transform 1 0 298256 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1698175906
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698175906
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_72
timestamp 1698175906
transform 1 0 9408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_136
timestamp 1698175906
transform 1 0 16576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_142
timestamp 1698175906
transform 1 0 17248 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698175906
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_212
timestamp 1698175906
transform 1 0 25088 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_276
timestamp 1698175906
transform 1 0 32256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_282
timestamp 1698175906
transform 1 0 32928 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_346
timestamp 1698175906
transform 1 0 40096 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_352
timestamp 1698175906
transform 1 0 40768 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_416
timestamp 1698175906
transform 1 0 47936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_422
timestamp 1698175906
transform 1 0 48608 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_486
timestamp 1698175906
transform 1 0 55776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_492
timestamp 1698175906
transform 1 0 56448 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_556
timestamp 1698175906
transform 1 0 63616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_562
timestamp 1698175906
transform 1 0 64288 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_626
timestamp 1698175906
transform 1 0 71456 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_632
timestamp 1698175906
transform 1 0 72128 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_696
timestamp 1698175906
transform 1 0 79296 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_702
timestamp 1698175906
transform 1 0 79968 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_766
timestamp 1698175906
transform 1 0 87136 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_772
timestamp 1698175906
transform 1 0 87808 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_836
timestamp 1698175906
transform 1 0 94976 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_842
timestamp 1698175906
transform 1 0 95648 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_906
timestamp 1698175906
transform 1 0 102816 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_912
timestamp 1698175906
transform 1 0 103488 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_976
timestamp 1698175906
transform 1 0 110656 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_982
timestamp 1698175906
transform 1 0 111328 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1046
timestamp 1698175906
transform 1 0 118496 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1052
timestamp 1698175906
transform 1 0 119168 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1116
timestamp 1698175906
transform 1 0 126336 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1122
timestamp 1698175906
transform 1 0 127008 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1186
timestamp 1698175906
transform 1 0 134176 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1192
timestamp 1698175906
transform 1 0 134848 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1256
timestamp 1698175906
transform 1 0 142016 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1262
timestamp 1698175906
transform 1 0 142688 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1326
timestamp 1698175906
transform 1 0 149856 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1332
timestamp 1698175906
transform 1 0 150528 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1396
timestamp 1698175906
transform 1 0 157696 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1402
timestamp 1698175906
transform 1 0 158368 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1466
timestamp 1698175906
transform 1 0 165536 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1472
timestamp 1698175906
transform 1 0 166208 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1536
timestamp 1698175906
transform 1 0 173376 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1542
timestamp 1698175906
transform 1 0 174048 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_1606
timestamp 1698175906
transform 1 0 181216 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_1612
timestamp 1698175906
transform 1 0 181888 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_1645
timestamp 1698175906
transform 1 0 185584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_1649
timestamp 1698175906
transform 1 0 186032 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1682
timestamp 1698175906
transform 1 0 189728 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1746
timestamp 1698175906
transform 1 0 196896 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1752
timestamp 1698175906
transform 1 0 197568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1816
timestamp 1698175906
transform 1 0 204736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1822
timestamp 1698175906
transform 1 0 205408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1886
timestamp 1698175906
transform 1 0 212576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1892
timestamp 1698175906
transform 1 0 213248 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1956
timestamp 1698175906
transform 1 0 220416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1962
timestamp 1698175906
transform 1 0 221088 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2026
timestamp 1698175906
transform 1 0 228256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2032
timestamp 1698175906
transform 1 0 228928 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2096
timestamp 1698175906
transform 1 0 236096 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2102
timestamp 1698175906
transform 1 0 236768 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2166
timestamp 1698175906
transform 1 0 243936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2172
timestamp 1698175906
transform 1 0 244608 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2236
timestamp 1698175906
transform 1 0 251776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2242
timestamp 1698175906
transform 1 0 252448 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2306
timestamp 1698175906
transform 1 0 259616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2312
timestamp 1698175906
transform 1 0 260288 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2376
timestamp 1698175906
transform 1 0 267456 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2382
timestamp 1698175906
transform 1 0 268128 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2446
timestamp 1698175906
transform 1 0 275296 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2452
timestamp 1698175906
transform 1 0 275968 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2516
timestamp 1698175906
transform 1 0 283136 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2522
timestamp 1698175906
transform 1 0 283808 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2586
timestamp 1698175906
transform 1 0 290976 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_2592
timestamp 1698175906
transform 1 0 291648 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_2624
timestamp 1698175906
transform 1 0 295232 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_2640
timestamp 1698175906
transform 1 0 297024 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2648
timestamp 1698175906
transform 1 0 297920 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698175906
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698175906
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698175906
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698175906
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_107
timestamp 1698175906
transform 1 0 13328 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_171
timestamp 1698175906
transform 1 0 20496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_177
timestamp 1698175906
transform 1 0 21168 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_241
timestamp 1698175906
transform 1 0 28336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_247
timestamp 1698175906
transform 1 0 29008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698175906
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_317
timestamp 1698175906
transform 1 0 36848 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_381
timestamp 1698175906
transform 1 0 44016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_387
timestamp 1698175906
transform 1 0 44688 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698175906
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_457
timestamp 1698175906
transform 1 0 52528 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_521
timestamp 1698175906
transform 1 0 59696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_527
timestamp 1698175906
transform 1 0 60368 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_591
timestamp 1698175906
transform 1 0 67536 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_597
timestamp 1698175906
transform 1 0 68208 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_661
timestamp 1698175906
transform 1 0 75376 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_667
timestamp 1698175906
transform 1 0 76048 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_731
timestamp 1698175906
transform 1 0 83216 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_737
timestamp 1698175906
transform 1 0 83888 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_801
timestamp 1698175906
transform 1 0 91056 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_807
timestamp 1698175906
transform 1 0 91728 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_871
timestamp 1698175906
transform 1 0 98896 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_877
timestamp 1698175906
transform 1 0 99568 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_941
timestamp 1698175906
transform 1 0 106736 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_947
timestamp 1698175906
transform 1 0 107408 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1011
timestamp 1698175906
transform 1 0 114576 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1017
timestamp 1698175906
transform 1 0 115248 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1081
timestamp 1698175906
transform 1 0 122416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_1087
timestamp 1698175906
transform 1 0 123088 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_1119
timestamp 1698175906
transform 1 0 126672 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1135
timestamp 1698175906
transform 1 0 128464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1153
timestamp 1698175906
transform 1 0 130480 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1157
timestamp 1698175906
transform 1 0 130928 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1221
timestamp 1698175906
transform 1 0 138096 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_1227
timestamp 1698175906
transform 1 0 138768 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_1259
timestamp 1698175906
transform 1 0 142352 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_1275
timestamp 1698175906
transform 1 0 144144 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1293
timestamp 1698175906
transform 1 0 146160 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_1297
timestamp 1698175906
transform 1 0 146608 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1329
timestamp 1698175906
transform 1 0 150192 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_1343
timestamp 1698175906
transform 1 0 151760 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1359
timestamp 1698175906
transform 1 0 153552 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1363
timestamp 1698175906
transform 1 0 154000 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1367
timestamp 1698175906
transform 1 0 154448 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1431
timestamp 1698175906
transform 1 0 161616 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_1487
timestamp 1698175906
transform 1 0 167888 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1503
timestamp 1698175906
transform 1 0 169680 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1507
timestamp 1698175906
transform 1 0 170128 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1571
timestamp 1698175906
transform 1 0 177296 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_1627
timestamp 1698175906
transform 1 0 183568 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1643
timestamp 1698175906
transform 1 0 185360 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_1647
timestamp 1698175906
transform 1 0 185808 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_1663
timestamp 1698175906
transform 1 0 187600 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1671
timestamp 1698175906
transform 1 0 188496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1675
timestamp 1698175906
transform 1 0 188944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_1677
timestamp 1698175906
transform 1 0 189168 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1680
timestamp 1698175906
transform 1 0 189504 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1684
timestamp 1698175906
transform 1 0 189952 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1717
timestamp 1698175906
transform 1 0 193648 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1781
timestamp 1698175906
transform 1 0 200816 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1787
timestamp 1698175906
transform 1 0 201488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1851
timestamp 1698175906
transform 1 0 208656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1857
timestamp 1698175906
transform 1 0 209328 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1921
timestamp 1698175906
transform 1 0 216496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1927
timestamp 1698175906
transform 1 0 217168 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1991
timestamp 1698175906
transform 1 0 224336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1997
timestamp 1698175906
transform 1 0 225008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2061
timestamp 1698175906
transform 1 0 232176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_2067
timestamp 1698175906
transform 1 0 232848 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2131
timestamp 1698175906
transform 1 0 240016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_2137
timestamp 1698175906
transform 1 0 240688 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2201
timestamp 1698175906
transform 1 0 247856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_2207
timestamp 1698175906
transform 1 0 248528 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2271
timestamp 1698175906
transform 1 0 255696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_2277
timestamp 1698175906
transform 1 0 256368 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2341
timestamp 1698175906
transform 1 0 263536 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_2347
timestamp 1698175906
transform 1 0 264208 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2411
timestamp 1698175906
transform 1 0 271376 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_2417
timestamp 1698175906
transform 1 0 272048 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2481
timestamp 1698175906
transform 1 0 279216 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_2487
timestamp 1698175906
transform 1 0 279888 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2551
timestamp 1698175906
transform 1 0 287056 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_2557
timestamp 1698175906
transform 1 0 287728 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2621
timestamp 1698175906
transform 1 0 294896 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_2627
timestamp 1698175906
transform 1 0 295568 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_2643
timestamp 1698175906
transform 1 0 297360 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_2651
timestamp 1698175906
transform 1 0 298256 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2
timestamp 1698175906
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698175906
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698175906
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698175906
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_142
timestamp 1698175906
transform 1 0 17248 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_206
timestamp 1698175906
transform 1 0 24416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_212
timestamp 1698175906
transform 1 0 25088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_276
timestamp 1698175906
transform 1 0 32256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_282
timestamp 1698175906
transform 1 0 32928 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_346
timestamp 1698175906
transform 1 0 40096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_352
timestamp 1698175906
transform 1 0 40768 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_416
timestamp 1698175906
transform 1 0 47936 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698175906
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698175906
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_492
timestamp 1698175906
transform 1 0 56448 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_556
timestamp 1698175906
transform 1 0 63616 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_562
timestamp 1698175906
transform 1 0 64288 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_626
timestamp 1698175906
transform 1 0 71456 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_632
timestamp 1698175906
transform 1 0 72128 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_696
timestamp 1698175906
transform 1 0 79296 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_702
timestamp 1698175906
transform 1 0 79968 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_766
timestamp 1698175906
transform 1 0 87136 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_772
timestamp 1698175906
transform 1 0 87808 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_836
timestamp 1698175906
transform 1 0 94976 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_842
timestamp 1698175906
transform 1 0 95648 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_906
timestamp 1698175906
transform 1 0 102816 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_912
timestamp 1698175906
transform 1 0 103488 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_976
timestamp 1698175906
transform 1 0 110656 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_982
timestamp 1698175906
transform 1 0 111328 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1046
timestamp 1698175906
transform 1 0 118496 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1052
timestamp 1698175906
transform 1 0 119168 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1116
timestamp 1698175906
transform 1 0 126336 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_1122
timestamp 1698175906
transform 1 0 127008 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1138
timestamp 1698175906
transform 1 0 128800 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1142
timestamp 1698175906
transform 1 0 129248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1173
timestamp 1698175906
transform 1 0 132720 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_1177
timestamp 1698175906
transform 1 0 133168 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1185
timestamp 1698175906
transform 1 0 134064 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1189
timestamp 1698175906
transform 1 0 134512 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_1202
timestamp 1698175906
transform 1 0 135968 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1234
timestamp 1698175906
transform 1 0 139552 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1238
timestamp 1698175906
transform 1 0 140000 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_1249
timestamp 1698175906
transform 1 0 141232 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1257
timestamp 1698175906
transform 1 0 142128 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1259
timestamp 1698175906
transform 1 0 142352 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_1262
timestamp 1698175906
transform 1 0 142688 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1278
timestamp 1698175906
transform 1 0 144480 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1282
timestamp 1698175906
transform 1 0 144928 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1313
timestamp 1698175906
transform 1 0 148400 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_1317
timestamp 1698175906
transform 1 0 148848 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1325
timestamp 1698175906
transform 1 0 149744 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1327
timestamp 1698175906
transform 1 0 149968 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1332
timestamp 1698175906
transform 1 0 150528 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1334
timestamp 1698175906
transform 1 0 150752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_1364
timestamp 1698175906
transform 1 0 154112 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1380
timestamp 1698175906
transform 1 0 155904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1382
timestamp 1698175906
transform 1 0 156128 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1393
timestamp 1698175906
transform 1 0 157360 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1397
timestamp 1698175906
transform 1 0 157808 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1399
timestamp 1698175906
transform 1 0 158032 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_1402
timestamp 1698175906
transform 1 0 158368 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_1418
timestamp 1698175906
transform 1 0 160160 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1426
timestamp 1698175906
transform 1 0 161056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1428
timestamp 1698175906
transform 1 0 161280 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_1439
timestamp 1698175906
transform 1 0 162512 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_1455
timestamp 1698175906
transform 1 0 164304 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1463
timestamp 1698175906
transform 1 0 165200 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1467
timestamp 1698175906
transform 1 0 165648 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1469
timestamp 1698175906
transform 1 0 165872 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1472
timestamp 1698175906
transform 1 0 166208 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1476
timestamp 1698175906
transform 1 0 166656 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1478
timestamp 1698175906
transform 1 0 166880 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_1489
timestamp 1698175906
transform 1 0 168112 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1521
timestamp 1698175906
transform 1 0 171696 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_1532
timestamp 1698175906
transform 1 0 172928 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1542
timestamp 1698175906
transform 1 0 174048 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1606
timestamp 1698175906
transform 1 0 181216 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_1612
timestamp 1698175906
transform 1 0 181888 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1620
timestamp 1698175906
transform 1 0 182784 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_1652
timestamp 1698175906
transform 1 0 186368 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_1668
timestamp 1698175906
transform 1 0 188160 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1676
timestamp 1698175906
transform 1 0 189056 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_1682
timestamp 1698175906
transform 1 0 189728 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1690
timestamp 1698175906
transform 1 0 190624 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1694
timestamp 1698175906
transform 1 0 191072 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1696
timestamp 1698175906
transform 1 0 191296 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_1728
timestamp 1698175906
transform 1 0 194880 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1744
timestamp 1698175906
transform 1 0 196672 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1748
timestamp 1698175906
transform 1 0 197120 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1752
timestamp 1698175906
transform 1 0 197568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1816
timestamp 1698175906
transform 1 0 204736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1822
timestamp 1698175906
transform 1 0 205408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1886
timestamp 1698175906
transform 1 0 212576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1892
timestamp 1698175906
transform 1 0 213248 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1956
timestamp 1698175906
transform 1 0 220416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1962
timestamp 1698175906
transform 1 0 221088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2026
timestamp 1698175906
transform 1 0 228256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2032
timestamp 1698175906
transform 1 0 228928 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2096
timestamp 1698175906
transform 1 0 236096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2102
timestamp 1698175906
transform 1 0 236768 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2166
timestamp 1698175906
transform 1 0 243936 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2172
timestamp 1698175906
transform 1 0 244608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2236
timestamp 1698175906
transform 1 0 251776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2242
timestamp 1698175906
transform 1 0 252448 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2306
timestamp 1698175906
transform 1 0 259616 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2312
timestamp 1698175906
transform 1 0 260288 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2376
timestamp 1698175906
transform 1 0 267456 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2382
timestamp 1698175906
transform 1 0 268128 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2446
timestamp 1698175906
transform 1 0 275296 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2452
timestamp 1698175906
transform 1 0 275968 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2516
timestamp 1698175906
transform 1 0 283136 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2522
timestamp 1698175906
transform 1 0 283808 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2586
timestamp 1698175906
transform 1 0 290976 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_2592
timestamp 1698175906
transform 1 0 291648 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_2624
timestamp 1698175906
transform 1 0 295232 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_2640
timestamp 1698175906
transform 1 0 297024 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2648
timestamp 1698175906
transform 1 0 297920 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698175906
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698175906
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698175906
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698175906
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_107
timestamp 1698175906
transform 1 0 13328 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_171
timestamp 1698175906
transform 1 0 20496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_177
timestamp 1698175906
transform 1 0 21168 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_241
timestamp 1698175906
transform 1 0 28336 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_247
timestamp 1698175906
transform 1 0 29008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_311
timestamp 1698175906
transform 1 0 36176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_317
timestamp 1698175906
transform 1 0 36848 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_381
timestamp 1698175906
transform 1 0 44016 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_387
timestamp 1698175906
transform 1 0 44688 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_451
timestamp 1698175906
transform 1 0 51856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_457
timestamp 1698175906
transform 1 0 52528 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_521
timestamp 1698175906
transform 1 0 59696 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_527
timestamp 1698175906
transform 1 0 60368 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_591
timestamp 1698175906
transform 1 0 67536 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_597
timestamp 1698175906
transform 1 0 68208 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_629
timestamp 1698175906
transform 1 0 71792 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_657
timestamp 1698175906
transform 1 0 74928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_661
timestamp 1698175906
transform 1 0 75376 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_667
timestamp 1698175906
transform 1 0 76048 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_731
timestamp 1698175906
transform 1 0 83216 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_737
timestamp 1698175906
transform 1 0 83888 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_801
timestamp 1698175906
transform 1 0 91056 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_807
timestamp 1698175906
transform 1 0 91728 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_871
timestamp 1698175906
transform 1 0 98896 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_903
timestamp 1698175906
transform 1 0 102480 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_907
timestamp 1698175906
transform 1 0 102928 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_939
timestamp 1698175906
transform 1 0 106512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_943
timestamp 1698175906
transform 1 0 106960 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_947
timestamp 1698175906
transform 1 0 107408 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1011
timestamp 1698175906
transform 1 0 114576 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_1017
timestamp 1698175906
transform 1 0 115248 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1081
timestamp 1698175906
transform 1 0 122416 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_1087
timestamp 1698175906
transform 1 0 123088 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1151
timestamp 1698175906
transform 1 0 130256 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_1157
timestamp 1698175906
transform 1 0 130928 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1189
timestamp 1698175906
transform 1 0 134512 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1191
timestamp 1698175906
transform 1 0 134736 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1221
timestamp 1698175906
transform 1 0 138096 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1227
timestamp 1698175906
transform 1 0 138768 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1235
timestamp 1698175906
transform 1 0 139664 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1239
timestamp 1698175906
transform 1 0 140112 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1270
timestamp 1698175906
transform 1 0 143584 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1274
timestamp 1698175906
transform 1 0 144032 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1290
timestamp 1698175906
transform 1 0 145824 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1294
timestamp 1698175906
transform 1 0 146272 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1297
timestamp 1698175906
transform 1 0 146608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1301
timestamp 1698175906
transform 1 0 147056 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1303
timestamp 1698175906
transform 1 0 147280 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1354
timestamp 1698175906
transform 1 0 152992 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1358
timestamp 1698175906
transform 1 0 153440 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1362
timestamp 1698175906
transform 1 0 153888 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1364
timestamp 1698175906
transform 1 0 154112 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1367
timestamp 1698175906
transform 1 0 154448 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1414
timestamp 1698175906
transform 1 0 159712 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1430
timestamp 1698175906
transform 1 0 161504 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1432
timestamp 1698175906
transform 1 0 161728 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1466
timestamp 1698175906
transform 1 0 165536 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1474
timestamp 1698175906
transform 1 0 166432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1507
timestamp 1698175906
transform 1 0 170128 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1511
timestamp 1698175906
transform 1 0 170576 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1519
timestamp 1698175906
transform 1 0 171472 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1523
timestamp 1698175906
transform 1 0 171920 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1553
timestamp 1698175906
transform 1 0 175280 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1557
timestamp 1698175906
transform 1 0 175728 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1573
timestamp 1698175906
transform 1 0 177520 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_1577
timestamp 1698175906
transform 1 0 177968 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1585
timestamp 1698175906
transform 1 0 178864 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1618
timestamp 1698175906
transform 1 0 182560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1622
timestamp 1698175906
transform 1 0 183008 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1638
timestamp 1698175906
transform 1 0 184800 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1642
timestamp 1698175906
transform 1 0 185248 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1644
timestamp 1698175906
transform 1 0 185472 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1660
timestamp 1698175906
transform 1 0 187264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1664
timestamp 1698175906
transform 1 0 187712 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_1697
timestamp 1698175906
transform 1 0 191408 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1713
timestamp 1698175906
transform 1 0 193200 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_1717
timestamp 1698175906
transform 1 0 193648 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1781
timestamp 1698175906
transform 1 0 200816 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_1787
timestamp 1698175906
transform 1 0 201488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1851
timestamp 1698175906
transform 1 0 208656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_1857
timestamp 1698175906
transform 1 0 209328 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1921
timestamp 1698175906
transform 1 0 216496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_1927
timestamp 1698175906
transform 1 0 217168 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1991
timestamp 1698175906
transform 1 0 224336 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_1997
timestamp 1698175906
transform 1 0 225008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2061
timestamp 1698175906
transform 1 0 232176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_2067
timestamp 1698175906
transform 1 0 232848 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2131
timestamp 1698175906
transform 1 0 240016 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_2137
timestamp 1698175906
transform 1 0 240688 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2201
timestamp 1698175906
transform 1 0 247856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_2207
timestamp 1698175906
transform 1 0 248528 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2271
timestamp 1698175906
transform 1 0 255696 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_2277
timestamp 1698175906
transform 1 0 256368 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2341
timestamp 1698175906
transform 1 0 263536 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_2347
timestamp 1698175906
transform 1 0 264208 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2411
timestamp 1698175906
transform 1 0 271376 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_2417
timestamp 1698175906
transform 1 0 272048 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2481
timestamp 1698175906
transform 1 0 279216 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_2487
timestamp 1698175906
transform 1 0 279888 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2551
timestamp 1698175906
transform 1 0 287056 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_2557
timestamp 1698175906
transform 1 0 287728 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2621
timestamp 1698175906
transform 1 0 294896 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_2627
timestamp 1698175906
transform 1 0 295568 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_2643
timestamp 1698175906
transform 1 0 297360 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_2651
timestamp 1698175906
transform 1 0 298256 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_2
timestamp 1698175906
transform 1 0 1568 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_36
timestamp 1698175906
transform 1 0 5376 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_70
timestamp 1698175906
transform 1 0 9184 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_86
timestamp 1698175906
transform 1 0 10976 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_94
timestamp 1698175906
transform 1 0 11872 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_98
timestamp 1698175906
transform 1 0 12320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_110
timestamp 1698175906
transform 1 0 13664 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_126
timestamp 1698175906
transform 1 0 15456 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_134
timestamp 1698175906
transform 1 0 16352 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_138
timestamp 1698175906
transform 1 0 16800 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_146
timestamp 1698175906
transform 1 0 17696 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_148
timestamp 1698175906
transform 1 0 17920 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_161
timestamp 1698175906
transform 1 0 19376 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_169
timestamp 1698175906
transform 1 0 20272 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_172
timestamp 1698175906
transform 1 0 20608 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_188
timestamp 1698175906
transform 1 0 22400 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_196
timestamp 1698175906
transform 1 0 23296 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_200
timestamp 1698175906
transform 1 0 23744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_214
timestamp 1698175906
transform 1 0 25312 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_230
timestamp 1698175906
transform 1 0 27104 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_240
timestamp 1698175906
transform 1 0 28224 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_244
timestamp 1698175906
transform 1 0 28672 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_255
timestamp 1698175906
transform 1 0 29904 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_271
timestamp 1698175906
transform 1 0 31696 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_274
timestamp 1698175906
transform 1 0 32032 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_290
timestamp 1698175906
transform 1 0 33824 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_292
timestamp 1698175906
transform 1 0 34048 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_303
timestamp 1698175906
transform 1 0 35280 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_305
timestamp 1698175906
transform 1 0 35504 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_308
timestamp 1698175906
transform 1 0 35840 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_324
timestamp 1698175906
transform 1 0 37632 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_332
timestamp 1698175906
transform 1 0 38528 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_336
timestamp 1698175906
transform 1 0 38976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_342
timestamp 1698175906
transform 1 0 39648 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_351
timestamp 1698175906
transform 1 0 40656 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_367
timestamp 1698175906
transform 1 0 42448 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_371
timestamp 1698175906
transform 1 0 42896 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_373
timestamp 1698175906
transform 1 0 43120 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_376
timestamp 1698175906
transform 1 0 43456 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_384
timestamp 1698175906
transform 1 0 44352 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_388
timestamp 1698175906
transform 1 0 44800 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_399
timestamp 1698175906
transform 1 0 46032 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_407
timestamp 1698175906
transform 1 0 46928 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_410
timestamp 1698175906
transform 1 0 47264 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_426
timestamp 1698175906
transform 1 0 49056 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_434
timestamp 1698175906
transform 1 0 49952 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_438
timestamp 1698175906
transform 1 0 50400 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_452
timestamp 1698175906
transform 1 0 51968 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_468
timestamp 1698175906
transform 1 0 53760 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_478
timestamp 1698175906
transform 1 0 54880 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_482
timestamp 1698175906
transform 1 0 55328 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_484
timestamp 1698175906
transform 1 0 55552 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_495
timestamp 1698175906
transform 1 0 56784 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_503
timestamp 1698175906
transform 1 0 57680 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_507
timestamp 1698175906
transform 1 0 58128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_509
timestamp 1698175906
transform 1 0 58352 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_512
timestamp 1698175906
transform 1 0 58688 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_528
timestamp 1698175906
transform 1 0 60480 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_532
timestamp 1698175906
transform 1 0 60928 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_543
timestamp 1698175906
transform 1 0 62160 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_546
timestamp 1698175906
transform 1 0 62496 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_580
timestamp 1698175906
transform 1 0 66304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_582
timestamp 1698175906
transform 1 0 66528 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_609
timestamp 1698175906
transform 1 0 69552 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_611
timestamp 1698175906
transform 1 0 69776 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_614
timestamp 1698175906
transform 1 0 70112 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_618
timestamp 1698175906
transform 1 0 70560 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_634
timestamp 1698175906
transform 1 0 72352 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_642
timestamp 1698175906
transform 1 0 73248 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_648
timestamp 1698175906
transform 1 0 73920 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_708
timestamp 1698175906
transform 1 0 80640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_712
timestamp 1698175906
transform 1 0 81088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_716
timestamp 1698175906
transform 1 0 81536 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_720
timestamp 1698175906
transform 1 0 81984 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_750
timestamp 1698175906
transform 1 0 85344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_754
timestamp 1698175906
transform 1 0 85792 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_770
timestamp 1698175906
transform 1 0 87584 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_778
timestamp 1698175906
transform 1 0 88480 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_810
timestamp 1698175906
transform 1 0 92064 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_814
timestamp 1698175906
transform 1 0 92512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_818
timestamp 1698175906
transform 1 0 92960 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_822
timestamp 1698175906
transform 1 0 93408 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_849
timestamp 1698175906
transform 1 0 96432 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_852
timestamp 1698175906
transform 1 0 96768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_856
timestamp 1698175906
transform 1 0 97216 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_872
timestamp 1698175906
transform 1 0 99008 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_880
timestamp 1698175906
transform 1 0 99904 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_886
timestamp 1698175906
transform 1 0 100576 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_946
timestamp 1698175906
transform 1 0 107296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_950
timestamp 1698175906
transform 1 0 107744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_954
timestamp 1698175906
transform 1 0 108192 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_962
timestamp 1698175906
transform 1 0 109088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_964
timestamp 1698175906
transform 1 0 109312 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_975
timestamp 1698175906
transform 1 0 110544 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_983
timestamp 1698175906
transform 1 0 111440 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_985
timestamp 1698175906
transform 1 0 111664 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_988
timestamp 1698175906
transform 1 0 112000 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1004
timestamp 1698175906
transform 1 0 113792 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1012
timestamp 1698175906
transform 1 0 114688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1016
timestamp 1698175906
transform 1 0 115136 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1030
timestamp 1698175906
transform 1 0 116704 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1046
timestamp 1698175906
transform 1 0 118496 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1056
timestamp 1698175906
transform 1 0 119616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1060
timestamp 1698175906
transform 1 0 120064 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1071
timestamp 1698175906
transform 1 0 121296 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1087
timestamp 1698175906
transform 1 0 123088 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1090
timestamp 1698175906
transform 1 0 123424 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1106
timestamp 1698175906
transform 1 0 125216 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1108
timestamp 1698175906
transform 1 0 125440 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1117
timestamp 1698175906
transform 1 0 126448 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1121
timestamp 1698175906
transform 1 0 126896 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1124
timestamp 1698175906
transform 1 0 127232 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1140
timestamp 1698175906
transform 1 0 129024 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1148
timestamp 1698175906
transform 1 0 129920 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1152
timestamp 1698175906
transform 1 0 130368 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1158
timestamp 1698175906
transform 1 0 131040 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1165
timestamp 1698175906
transform 1 0 131824 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1181
timestamp 1698175906
transform 1 0 133616 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1189
timestamp 1698175906
transform 1 0 134512 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1192
timestamp 1698175906
transform 1 0 134848 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1200
timestamp 1698175906
transform 1 0 135744 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1204
timestamp 1698175906
transform 1 0 136192 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1213
timestamp 1698175906
transform 1 0 137200 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1221
timestamp 1698175906
transform 1 0 138096 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1223
timestamp 1698175906
transform 1 0 138320 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1226
timestamp 1698175906
transform 1 0 138656 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1242
timestamp 1698175906
transform 1 0 140448 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1250
timestamp 1698175906
transform 1 0 141344 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1254
timestamp 1698175906
transform 1 0 141792 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1266
timestamp 1698175906
transform 1 0 143136 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1282
timestamp 1698175906
transform 1 0 144928 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1290
timestamp 1698175906
transform 1 0 145824 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1294
timestamp 1698175906
transform 1 0 146272 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1298
timestamp 1698175906
transform 1 0 146720 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1300
timestamp 1698175906
transform 1 0 146944 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1309
timestamp 1698175906
transform 1 0 147952 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1325
timestamp 1698175906
transform 1 0 149744 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1328
timestamp 1698175906
transform 1 0 150080 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1344
timestamp 1698175906
transform 1 0 151872 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1348
timestamp 1698175906
transform 1 0 152320 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1357
timestamp 1698175906
transform 1 0 153328 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1359
timestamp 1698175906
transform 1 0 153552 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1362
timestamp 1698175906
transform 1 0 153888 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1378
timestamp 1698175906
transform 1 0 155680 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1386
timestamp 1698175906
transform 1 0 156576 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1390
timestamp 1698175906
transform 1 0 157024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1396
timestamp 1698175906
transform 1 0 157696 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1398
timestamp 1698175906
transform 1 0 157920 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1405
timestamp 1698175906
transform 1 0 158704 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1421
timestamp 1698175906
transform 1 0 160496 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1425
timestamp 1698175906
transform 1 0 160944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1427
timestamp 1698175906
transform 1 0 161168 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1430
timestamp 1698175906
transform 1 0 161504 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1438
timestamp 1698175906
transform 1 0 162400 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1442
timestamp 1698175906
transform 1 0 162848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1444
timestamp 1698175906
transform 1 0 163072 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1453
timestamp 1698175906
transform 1 0 164080 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1461
timestamp 1698175906
transform 1 0 164976 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1464
timestamp 1698175906
transform 1 0 165312 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1480
timestamp 1698175906
transform 1 0 167104 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1488
timestamp 1698175906
transform 1 0 168000 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1492
timestamp 1698175906
transform 1 0 168448 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1504
timestamp 1698175906
transform 1 0 169792 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1520
timestamp 1698175906
transform 1 0 171584 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1528
timestamp 1698175906
transform 1 0 172480 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1532
timestamp 1698175906
transform 1 0 172928 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1540
timestamp 1698175906
transform 1 0 173824 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1549
timestamp 1698175906
transform 1 0 174832 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1557
timestamp 1698175906
transform 1 0 175728 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1561
timestamp 1698175906
transform 1 0 176176 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1563
timestamp 1698175906
transform 1 0 176400 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1566
timestamp 1698175906
transform 1 0 176736 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1582
timestamp 1698175906
transform 1 0 178528 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1586
timestamp 1698175906
transform 1 0 178976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1588
timestamp 1698175906
transform 1 0 179200 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1597
timestamp 1698175906
transform 1 0 180208 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_1600
timestamp 1698175906
transform 1 0 180544 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1634
timestamp 1698175906
transform 1 0 184352 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1636
timestamp 1698175906
transform 1 0 184576 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1645
timestamp 1698175906
transform 1 0 185584 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1661
timestamp 1698175906
transform 1 0 187376 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1663
timestamp 1698175906
transform 1 0 187600 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1702
timestamp 1698175906
transform 1 0 191968 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1706
timestamp 1698175906
transform 1 0 192416 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1722
timestamp 1698175906
transform 1 0 194208 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1730
timestamp 1698175906
transform 1 0 195104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1742
timestamp 1698175906
transform 1 0 196448 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1758
timestamp 1698175906
transform 1 0 198240 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1766
timestamp 1698175906
transform 1 0 199136 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1770
timestamp 1698175906
transform 1 0 199584 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1774
timestamp 1698175906
transform 1 0 200032 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1804
timestamp 1698175906
transform 1 0 203392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1808
timestamp 1698175906
transform 1 0 203840 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1824
timestamp 1698175906
transform 1 0 205632 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1832
timestamp 1698175906
transform 1 0 206528 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1864
timestamp 1698175906
transform 1 0 210112 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1868
timestamp 1698175906
transform 1 0 210560 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1872
timestamp 1698175906
transform 1 0 211008 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1876
timestamp 1698175906
transform 1 0 211456 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1885
timestamp 1698175906
transform 1 0 212464 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1901
timestamp 1698175906
transform 1 0 214256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1903
timestamp 1698175906
transform 1 0 214480 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1906
timestamp 1698175906
transform 1 0 214816 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1922
timestamp 1698175906
transform 1 0 216608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1924
timestamp 1698175906
transform 1 0 216832 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1933
timestamp 1698175906
transform 1 0 217840 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1937
timestamp 1698175906
transform 1 0 218288 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1940
timestamp 1698175906
transform 1 0 218624 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1956
timestamp 1698175906
transform 1 0 220416 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1964
timestamp 1698175906
transform 1 0 221312 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1968
timestamp 1698175906
transform 1 0 221760 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1974
timestamp 1698175906
transform 1 0 222432 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_1981
timestamp 1698175906
transform 1 0 223216 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_1997
timestamp 1698175906
transform 1 0 225008 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2005
timestamp 1698175906
transform 1 0 225904 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2008
timestamp 1698175906
transform 1 0 226240 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2016
timestamp 1698175906
transform 1 0 227136 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2020
timestamp 1698175906
transform 1 0 227584 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2029
timestamp 1698175906
transform 1 0 228592 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2037
timestamp 1698175906
transform 1 0 229488 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2039
timestamp 1698175906
transform 1 0 229712 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2042
timestamp 1698175906
transform 1 0 230048 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2058
timestamp 1698175906
transform 1 0 231840 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2066
timestamp 1698175906
transform 1 0 232736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2070
timestamp 1698175906
transform 1 0 233184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2082
timestamp 1698175906
transform 1 0 234528 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2098
timestamp 1698175906
transform 1 0 236320 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2106
timestamp 1698175906
transform 1 0 237216 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2110
timestamp 1698175906
transform 1 0 237664 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2114
timestamp 1698175906
transform 1 0 238112 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2116
timestamp 1698175906
transform 1 0 238336 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2127
timestamp 1698175906
transform 1 0 239568 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2135
timestamp 1698175906
transform 1 0 240464 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2139
timestamp 1698175906
transform 1 0 240912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2141
timestamp 1698175906
transform 1 0 241136 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2144
timestamp 1698175906
transform 1 0 241472 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2160
timestamp 1698175906
transform 1 0 243264 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2164
timestamp 1698175906
transform 1 0 243712 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2175
timestamp 1698175906
transform 1 0 244944 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2178
timestamp 1698175906
transform 1 0 245280 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2194
timestamp 1698175906
transform 1 0 247072 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2202
timestamp 1698175906
transform 1 0 247968 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2206
timestamp 1698175906
transform 1 0 248416 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2212
timestamp 1698175906
transform 1 0 249088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2214
timestamp 1698175906
transform 1 0 249312 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2223
timestamp 1698175906
transform 1 0 250320 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2239
timestamp 1698175906
transform 1 0 252112 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2243
timestamp 1698175906
transform 1 0 252560 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2246
timestamp 1698175906
transform 1 0 252896 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2254
timestamp 1698175906
transform 1 0 253792 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2258
timestamp 1698175906
transform 1 0 254240 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2260
timestamp 1698175906
transform 1 0 254464 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2277
timestamp 1698175906
transform 1 0 256368 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2280
timestamp 1698175906
transform 1 0 256704 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2296
timestamp 1698175906
transform 1 0 258496 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2304
timestamp 1698175906
transform 1 0 259392 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2308
timestamp 1698175906
transform 1 0 259840 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2328
timestamp 1698175906
transform 1 0 262080 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2344
timestamp 1698175906
transform 1 0 263872 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2348
timestamp 1698175906
transform 1 0 264320 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2356
timestamp 1698175906
transform 1 0 265216 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2373
timestamp 1698175906
transform 1 0 267120 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2377
timestamp 1698175906
transform 1 0 267568 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2379
timestamp 1698175906
transform 1 0 267792 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2382
timestamp 1698175906
transform 1 0 268128 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2398
timestamp 1698175906
transform 1 0 269920 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2406
timestamp 1698175906
transform 1 0 270816 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2410
timestamp 1698175906
transform 1 0 271264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2430
timestamp 1698175906
transform 1 0 273504 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2446
timestamp 1698175906
transform 1 0 275296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2450
timestamp 1698175906
transform 1 0 275744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2452
timestamp 1698175906
transform 1 0 275968 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2469
timestamp 1698175906
transform 1 0 277872 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2477
timestamp 1698175906
transform 1 0 278768 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2481
timestamp 1698175906
transform 1 0 279216 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2484
timestamp 1698175906
transform 1 0 279552 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2500
timestamp 1698175906
transform 1 0 281344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2518
timestamp 1698175906
transform 1 0 283360 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2522
timestamp 1698175906
transform 1 0 283808 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2538
timestamp 1698175906
transform 1 0 285600 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2546
timestamp 1698175906
transform 1 0 286496 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2562
timestamp 1698175906
transform 1 0 288288 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2578
timestamp 1698175906
transform 1 0 290080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2582
timestamp 1698175906
transform 1 0 290528 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2586
timestamp 1698175906
transform 1 0 290976 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2594
timestamp 1698175906
transform 1 0 291872 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2596
timestamp 1698175906
transform 1 0 292096 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_2609
timestamp 1698175906
transform 1 0 293552 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_2617
timestamp 1698175906
transform 1 0 294448 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_2620
timestamp 1698175906
transform 1 0 294784 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698175906
transform 1 0 123424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2
timestamp 1698175906
transform 1 0 127232 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input3
timestamp 1698175906
transform 1 0 131040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698175906
transform 1 0 133840 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698175906
transform 1 0 137424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input6
timestamp 1698175906
transform 1 0 141008 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698175906
transform 1 0 144592 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698175906
transform 1 0 148176 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698175906
transform 1 0 151760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input10
timestamp 1698175906
transform 1 0 155344 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input11
timestamp 1698175906
transform 1 0 158928 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input12
timestamp 1698175906
transform 1 0 162512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input13
timestamp 1698175906
transform 1 0 166096 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input14
timestamp 1698175906
transform 1 0 169680 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698175906
transform 1 0 173264 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698175906
transform 1 0 176848 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input17
timestamp 1698175906
transform 1 0 180544 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input18
timestamp 1698175906
transform 1 0 183456 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input19
timestamp 1698175906
transform -1 0 188832 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input20
timestamp 1698175906
transform 1 0 191072 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input21
timestamp 1698175906
transform 1 0 195776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698175906
transform -1 0 199024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input23
timestamp 1698175906
transform -1 0 206416 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698175906
transform -1 0 207872 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698175906
transform -1 0 210336 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698175906
transform -1 0 213360 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698175906
transform -1 0 216944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698175906
transform 1 0 219408 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698175906
transform -1 0 224112 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698175906
transform -1 0 227696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698175906
transform -1 0 231280 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698175906
transform -1 0 234864 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698175906
transform -1 0 238448 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698175906
transform -1 0 242144 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698175906
transform -1 0 245952 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698175906
transform -1 0 249760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698175906
transform -1 0 253568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698175906
transform -1 0 256368 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input39
timestamp 1698175906
transform -1 0 259952 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input40
timestamp 1698175906
transform -1 0 263536 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input41
timestamp 1698175906
transform 1 0 266448 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input42
timestamp 1698175906
transform 1 0 270032 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input43
timestamp 1698175906
transform 1 0 273616 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input44
timestamp 1698175906
transform 1 0 277200 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input45
timestamp 1698175906
transform 1 0 280784 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input46
timestamp 1698175906
transform 1 0 284368 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input47
timestamp 1698175906
transform 1 0 287952 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input48
timestamp 1698175906
transform 1 0 291536 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input49
timestamp 1698175906
transform 1 0 211792 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input50
timestamp 1698175906
transform -1 0 217840 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input51
timestamp 1698175906
transform -1 0 223216 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input52
timestamp 1698175906
transform -1 0 228592 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input53
timestamp 1698175906
transform -1 0 234528 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input54
timestamp 1698175906
transform 1 0 238672 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input55
timestamp 1698175906
transform 1 0 244048 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input56
timestamp 1698175906
transform 1 0 249424 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input57
timestamp 1698175906
transform 1 0 254800 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input58
timestamp 1698175906
transform 1 0 260512 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input59
timestamp 1698175906
transform 1 0 265552 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input60
timestamp 1698175906
transform 1 0 271936 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input61
timestamp 1698175906
transform 1 0 276304 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input62
timestamp 1698175906
transform -1 0 283136 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  input63
timestamp 1698175906
transform 1 0 287168 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  input64
timestamp 1698175906
transform 1 0 292432 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  input65
timestamp 1698175906
transform 1 0 18256 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input66
timestamp 1698175906
transform 1 0 24416 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input67
timestamp 1698175906
transform 1 0 29008 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input68
timestamp 1698175906
transform 1 0 34384 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input69
timestamp 1698175906
transform 1 0 39760 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input70
timestamp 1698175906
transform 1 0 45136 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input71
timestamp 1698175906
transform 1 0 51072 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input72
timestamp 1698175906
transform 1 0 55888 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input73
timestamp 1698175906
transform 1 0 61264 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input74
timestamp 1698175906
transform 1 0 109648 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input75
timestamp 1698175906
transform 1 0 115808 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1698175906
transform -1 0 169792 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input77
timestamp 1698175906
transform -1 0 174832 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1698175906
transform 1 0 179536 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input79
timestamp 1698175906
transform -1 0 185584 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input80
timestamp 1698175906
transform -1 0 191744 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input81
timestamp 1698175906
transform -1 0 196448 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input82
timestamp 1698175906
transform 1 0 120400 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input83
timestamp 1698175906
transform 1 0 125776 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input84
timestamp 1698175906
transform 1 0 131152 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input85
timestamp 1698175906
transform -1 0 137200 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input86
timestamp 1698175906
transform -1 0 143136 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input87
timestamp 1698175906
transform -1 0 147952 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input88
timestamp 1698175906
transform 1 0 152656 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input89
timestamp 1698175906
transform -1 0 158704 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input90
timestamp 1698175906
transform -1 0 164080 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input91
timestamp 1698175906
transform -1 0 13664 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output92 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 43232 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output93
timestamp 1698175906
transform -1 0 47040 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output94
timestamp 1698175906
transform -1 0 50736 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output95
timestamp 1698175906
transform -1 0 54320 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output96
timestamp 1698175906
transform -1 0 57904 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output97
timestamp 1698175906
transform -1 0 61600 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output98
timestamp 1698175906
transform -1 0 65408 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output99
timestamp 1698175906
transform -1 0 69216 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output100
timestamp 1698175906
transform -1 0 73024 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output101
timestamp 1698175906
transform -1 0 12096 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output102
timestamp 1698175906
transform 1 0 73920 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output103
timestamp 1698175906
transform 1 0 76496 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output104
timestamp 1698175906
transform 1 0 80080 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output105
timestamp 1698175906
transform 1 0 83664 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output106
timestamp 1698175906
transform 1 0 87808 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output107
timestamp 1698175906
transform 1 0 90832 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output108
timestamp 1698175906
transform 1 0 93632 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output109
timestamp 1698175906
transform 1 0 97440 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output110
timestamp 1698175906
transform -1 0 104160 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output111
timestamp 1698175906
transform -1 0 107968 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output112
timestamp 1698175906
transform -1 0 111664 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output113
timestamp 1698175906
transform -1 0 115248 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output114
timestamp 1698175906
transform -1 0 118832 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output115
timestamp 1698175906
transform -1 0 122528 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output116
timestamp 1698175906
transform -1 0 203168 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output117
timestamp 1698175906
transform 1 0 207200 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output118
timestamp 1698175906
transform -1 0 69552 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output119
timestamp 1698175906
transform -1 0 74928 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output120
timestamp 1698175906
transform -1 0 80640 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output121
timestamp 1698175906
transform -1 0 85120 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output122
timestamp 1698175906
transform -1 0 92064 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output123
timestamp 1698175906
transform -1 0 96432 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output124
timestamp 1698175906
transform -1 0 102480 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output125
timestamp 1698175906
transform -1 0 107296 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 298592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 298592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 298592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 298592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 298592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 298592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 298592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 298592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 298592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 298592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 298592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 298592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 298592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 298592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 298592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 298592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 298592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 298592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 298592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 298592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 298592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 298592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 298592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 298592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 298592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 298592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 298592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 298592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 298592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 298592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 298592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 298592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 298592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 298592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 298592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 298592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 298592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 298592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 298592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 298592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 298592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 298592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 298592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 298592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 298592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698175906
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698175906
transform -1 0 298592 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698175906
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698175906
transform -1 0 298592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698175906
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698175906
transform -1 0 298592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698175906
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698175906
transform -1 0 298592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698175906
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698175906
transform -1 0 298592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698175906
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698175906
transform -1 0 298592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698175906
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698175906
transform -1 0 298592 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698175906
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698175906
transform -1 0 298592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698175906
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698175906
transform -1 0 298592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698175906
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698175906
transform -1 0 298592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698175906
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698175906
transform -1 0 298592 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698175906
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698175906
transform -1 0 298592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698175906
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698175906
transform -1 0 298592 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698175906
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698175906
transform -1 0 298592 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698175906
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698175906
transform -1 0 298592 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698175906
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698175906
transform -1 0 298592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698175906
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698175906
transform -1 0 298592 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698175906
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698175906
transform -1 0 298592 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698175906
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698175906
transform -1 0 298592 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698175906
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698175906
transform -1 0 298592 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698175906
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698175906
transform -1 0 298592 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698175906
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698175906
transform -1 0 298592 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698175906
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698175906
transform -1 0 298592 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_126 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12544 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_127
timestamp 1698175906
transform -1 0 16016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_128
timestamp 1698175906
transform -1 0 19600 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_129
timestamp 1698175906
transform -1 0 23184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_130
timestamp 1698175906
transform -1 0 26768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_131
timestamp 1698175906
transform -1 0 30352 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_132
timestamp 1698175906
transform -1 0 33936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_133
timestamp 1698175906
transform -1 0 37520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698175906
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698175906
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698175906
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698175906
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_150
timestamp 1698175906
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_151
timestamp 1698175906
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_152
timestamp 1698175906
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_153
timestamp 1698175906
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_154
timestamp 1698175906
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_155
timestamp 1698175906
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_156
timestamp 1698175906
transform 1 0 81312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_157
timestamp 1698175906
transform 1 0 85120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_158
timestamp 1698175906
transform 1 0 88928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_159
timestamp 1698175906
transform 1 0 92736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_160
timestamp 1698175906
transform 1 0 96544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_161
timestamp 1698175906
transform 1 0 100352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_162
timestamp 1698175906
transform 1 0 104160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_163
timestamp 1698175906
transform 1 0 107968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_164
timestamp 1698175906
transform 1 0 111776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_165
timestamp 1698175906
transform 1 0 115584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_166
timestamp 1698175906
transform 1 0 119392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_167
timestamp 1698175906
transform 1 0 123200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_168
timestamp 1698175906
transform 1 0 127008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_169
timestamp 1698175906
transform 1 0 130816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_170
timestamp 1698175906
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_171
timestamp 1698175906
transform 1 0 138432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_172
timestamp 1698175906
transform 1 0 142240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_173
timestamp 1698175906
transform 1 0 146048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_174
timestamp 1698175906
transform 1 0 149856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_175
timestamp 1698175906
transform 1 0 153664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_176
timestamp 1698175906
transform 1 0 157472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_177
timestamp 1698175906
transform 1 0 161280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_178
timestamp 1698175906
transform 1 0 165088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_179
timestamp 1698175906
transform 1 0 168896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_180
timestamp 1698175906
transform 1 0 172704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_181
timestamp 1698175906
transform 1 0 176512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_182
timestamp 1698175906
transform 1 0 180320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_183
timestamp 1698175906
transform 1 0 184128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_184
timestamp 1698175906
transform 1 0 187936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_185
timestamp 1698175906
transform 1 0 191744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_186
timestamp 1698175906
transform 1 0 195552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_187
timestamp 1698175906
transform 1 0 199360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_188
timestamp 1698175906
transform 1 0 203168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_189
timestamp 1698175906
transform 1 0 206976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_190
timestamp 1698175906
transform 1 0 210784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_191
timestamp 1698175906
transform 1 0 214592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_192
timestamp 1698175906
transform 1 0 218400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_193
timestamp 1698175906
transform 1 0 222208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_194
timestamp 1698175906
transform 1 0 226016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_195
timestamp 1698175906
transform 1 0 229824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_196
timestamp 1698175906
transform 1 0 233632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_197
timestamp 1698175906
transform 1 0 237440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_198
timestamp 1698175906
transform 1 0 241248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_199
timestamp 1698175906
transform 1 0 245056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_200
timestamp 1698175906
transform 1 0 248864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_201
timestamp 1698175906
transform 1 0 252672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_202
timestamp 1698175906
transform 1 0 256480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_203
timestamp 1698175906
transform 1 0 260288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_204
timestamp 1698175906
transform 1 0 264096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_205
timestamp 1698175906
transform 1 0 267904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_206
timestamp 1698175906
transform 1 0 271712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_207
timestamp 1698175906
transform 1 0 275520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_208
timestamp 1698175906
transform 1 0 279328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_209
timestamp 1698175906
transform 1 0 283136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_210
timestamp 1698175906
transform 1 0 286944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_211
timestamp 1698175906
transform 1 0 290752 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_212
timestamp 1698175906
transform 1 0 294560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_213
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_214
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_215
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_216
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_217
timestamp 1698175906
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_218
timestamp 1698175906
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_219
timestamp 1698175906
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_220
timestamp 1698175906
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_221
timestamp 1698175906
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_222
timestamp 1698175906
transform 1 0 79744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_223
timestamp 1698175906
transform 1 0 87584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_224
timestamp 1698175906
transform 1 0 95424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_225
timestamp 1698175906
transform 1 0 103264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_226
timestamp 1698175906
transform 1 0 111104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_227
timestamp 1698175906
transform 1 0 118944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_228
timestamp 1698175906
transform 1 0 126784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_229
timestamp 1698175906
transform 1 0 134624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_230
timestamp 1698175906
transform 1 0 142464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_231
timestamp 1698175906
transform 1 0 150304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_232
timestamp 1698175906
transform 1 0 158144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_233
timestamp 1698175906
transform 1 0 165984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_234
timestamp 1698175906
transform 1 0 173824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_235
timestamp 1698175906
transform 1 0 181664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_236
timestamp 1698175906
transform 1 0 189504 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_237
timestamp 1698175906
transform 1 0 197344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_238
timestamp 1698175906
transform 1 0 205184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_239
timestamp 1698175906
transform 1 0 213024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_240
timestamp 1698175906
transform 1 0 220864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_241
timestamp 1698175906
transform 1 0 228704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_242
timestamp 1698175906
transform 1 0 236544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_243
timestamp 1698175906
transform 1 0 244384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_244
timestamp 1698175906
transform 1 0 252224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_245
timestamp 1698175906
transform 1 0 260064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_246
timestamp 1698175906
transform 1 0 267904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_247
timestamp 1698175906
transform 1 0 275744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_248
timestamp 1698175906
transform 1 0 283584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_249
timestamp 1698175906
transform 1 0 291424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_250
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_251
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_252
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_253
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_254
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_255
timestamp 1698175906
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_256
timestamp 1698175906
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_257
timestamp 1698175906
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_258
timestamp 1698175906
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_259
timestamp 1698175906
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_260
timestamp 1698175906
transform 1 0 83664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_261
timestamp 1698175906
transform 1 0 91504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_262
timestamp 1698175906
transform 1 0 99344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_263
timestamp 1698175906
transform 1 0 107184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_264
timestamp 1698175906
transform 1 0 115024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_265
timestamp 1698175906
transform 1 0 122864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_266
timestamp 1698175906
transform 1 0 130704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_267
timestamp 1698175906
transform 1 0 138544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_268
timestamp 1698175906
transform 1 0 146384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_269
timestamp 1698175906
transform 1 0 154224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_270
timestamp 1698175906
transform 1 0 162064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_271
timestamp 1698175906
transform 1 0 169904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_272
timestamp 1698175906
transform 1 0 177744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_273
timestamp 1698175906
transform 1 0 185584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_274
timestamp 1698175906
transform 1 0 193424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_275
timestamp 1698175906
transform 1 0 201264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_276
timestamp 1698175906
transform 1 0 209104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_277
timestamp 1698175906
transform 1 0 216944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_278
timestamp 1698175906
transform 1 0 224784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_279
timestamp 1698175906
transform 1 0 232624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_280
timestamp 1698175906
transform 1 0 240464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_281
timestamp 1698175906
transform 1 0 248304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_282
timestamp 1698175906
transform 1 0 256144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_283
timestamp 1698175906
transform 1 0 263984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_284
timestamp 1698175906
transform 1 0 271824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_285
timestamp 1698175906
transform 1 0 279664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_286
timestamp 1698175906
transform 1 0 287504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_287
timestamp 1698175906
transform 1 0 295344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_288
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_289
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_290
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_291
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_292
timestamp 1698175906
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_293
timestamp 1698175906
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_294
timestamp 1698175906
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_295
timestamp 1698175906
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_296
timestamp 1698175906
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_297
timestamp 1698175906
transform 1 0 79744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_298
timestamp 1698175906
transform 1 0 87584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_299
timestamp 1698175906
transform 1 0 95424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_300
timestamp 1698175906
transform 1 0 103264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_301
timestamp 1698175906
transform 1 0 111104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_302
timestamp 1698175906
transform 1 0 118944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_303
timestamp 1698175906
transform 1 0 126784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_304
timestamp 1698175906
transform 1 0 134624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_305
timestamp 1698175906
transform 1 0 142464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_306
timestamp 1698175906
transform 1 0 150304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_307
timestamp 1698175906
transform 1 0 158144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_308
timestamp 1698175906
transform 1 0 165984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_309
timestamp 1698175906
transform 1 0 173824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_310
timestamp 1698175906
transform 1 0 181664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_311
timestamp 1698175906
transform 1 0 189504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_312
timestamp 1698175906
transform 1 0 197344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_313
timestamp 1698175906
transform 1 0 205184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_314
timestamp 1698175906
transform 1 0 213024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_315
timestamp 1698175906
transform 1 0 220864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_316
timestamp 1698175906
transform 1 0 228704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_317
timestamp 1698175906
transform 1 0 236544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_318
timestamp 1698175906
transform 1 0 244384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_319
timestamp 1698175906
transform 1 0 252224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_320
timestamp 1698175906
transform 1 0 260064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_321
timestamp 1698175906
transform 1 0 267904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_322
timestamp 1698175906
transform 1 0 275744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_323
timestamp 1698175906
transform 1 0 283584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_324
timestamp 1698175906
transform 1 0 291424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_325
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_326
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_327
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_328
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_329
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_330
timestamp 1698175906
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_331
timestamp 1698175906
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_332
timestamp 1698175906
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_333
timestamp 1698175906
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_334
timestamp 1698175906
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_335
timestamp 1698175906
transform 1 0 83664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_336
timestamp 1698175906
transform 1 0 91504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_337
timestamp 1698175906
transform 1 0 99344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_338
timestamp 1698175906
transform 1 0 107184 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_339
timestamp 1698175906
transform 1 0 115024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_340
timestamp 1698175906
transform 1 0 122864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_341
timestamp 1698175906
transform 1 0 130704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_342
timestamp 1698175906
transform 1 0 138544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_343
timestamp 1698175906
transform 1 0 146384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_344
timestamp 1698175906
transform 1 0 154224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_345
timestamp 1698175906
transform 1 0 162064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_346
timestamp 1698175906
transform 1 0 169904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_347
timestamp 1698175906
transform 1 0 177744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_348
timestamp 1698175906
transform 1 0 185584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_349
timestamp 1698175906
transform 1 0 193424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_350
timestamp 1698175906
transform 1 0 201264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_351
timestamp 1698175906
transform 1 0 209104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_352
timestamp 1698175906
transform 1 0 216944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_353
timestamp 1698175906
transform 1 0 224784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_354
timestamp 1698175906
transform 1 0 232624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_355
timestamp 1698175906
transform 1 0 240464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_356
timestamp 1698175906
transform 1 0 248304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_357
timestamp 1698175906
transform 1 0 256144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_358
timestamp 1698175906
transform 1 0 263984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_359
timestamp 1698175906
transform 1 0 271824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_360
timestamp 1698175906
transform 1 0 279664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_361
timestamp 1698175906
transform 1 0 287504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_362
timestamp 1698175906
transform 1 0 295344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_363
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_364
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_365
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_366
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_367
timestamp 1698175906
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_368
timestamp 1698175906
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_369
timestamp 1698175906
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_370
timestamp 1698175906
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_371
timestamp 1698175906
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_372
timestamp 1698175906
transform 1 0 79744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_373
timestamp 1698175906
transform 1 0 87584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_374
timestamp 1698175906
transform 1 0 95424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_375
timestamp 1698175906
transform 1 0 103264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_376
timestamp 1698175906
transform 1 0 111104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_377
timestamp 1698175906
transform 1 0 118944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_378
timestamp 1698175906
transform 1 0 126784 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_379
timestamp 1698175906
transform 1 0 134624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_380
timestamp 1698175906
transform 1 0 142464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_381
timestamp 1698175906
transform 1 0 150304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_382
timestamp 1698175906
transform 1 0 158144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_383
timestamp 1698175906
transform 1 0 165984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_384
timestamp 1698175906
transform 1 0 173824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_385
timestamp 1698175906
transform 1 0 181664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_386
timestamp 1698175906
transform 1 0 189504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_387
timestamp 1698175906
transform 1 0 197344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_388
timestamp 1698175906
transform 1 0 205184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_389
timestamp 1698175906
transform 1 0 213024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_390
timestamp 1698175906
transform 1 0 220864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_391
timestamp 1698175906
transform 1 0 228704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_392
timestamp 1698175906
transform 1 0 236544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_393
timestamp 1698175906
transform 1 0 244384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_394
timestamp 1698175906
transform 1 0 252224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_395
timestamp 1698175906
transform 1 0 260064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_396
timestamp 1698175906
transform 1 0 267904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_397
timestamp 1698175906
transform 1 0 275744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_398
timestamp 1698175906
transform 1 0 283584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_399
timestamp 1698175906
transform 1 0 291424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_400
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_401
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_402
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_403
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_404
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_405
timestamp 1698175906
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_406
timestamp 1698175906
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_407
timestamp 1698175906
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_408
timestamp 1698175906
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_409
timestamp 1698175906
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_410
timestamp 1698175906
transform 1 0 83664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_411
timestamp 1698175906
transform 1 0 91504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_412
timestamp 1698175906
transform 1 0 99344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_413
timestamp 1698175906
transform 1 0 107184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_414
timestamp 1698175906
transform 1 0 115024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_415
timestamp 1698175906
transform 1 0 122864 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_416
timestamp 1698175906
transform 1 0 130704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_417
timestamp 1698175906
transform 1 0 138544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_418
timestamp 1698175906
transform 1 0 146384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_419
timestamp 1698175906
transform 1 0 154224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_420
timestamp 1698175906
transform 1 0 162064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_421
timestamp 1698175906
transform 1 0 169904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_422
timestamp 1698175906
transform 1 0 177744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_423
timestamp 1698175906
transform 1 0 185584 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_424
timestamp 1698175906
transform 1 0 193424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_425
timestamp 1698175906
transform 1 0 201264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_426
timestamp 1698175906
transform 1 0 209104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_427
timestamp 1698175906
transform 1 0 216944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_428
timestamp 1698175906
transform 1 0 224784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_429
timestamp 1698175906
transform 1 0 232624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_430
timestamp 1698175906
transform 1 0 240464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_431
timestamp 1698175906
transform 1 0 248304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_432
timestamp 1698175906
transform 1 0 256144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_433
timestamp 1698175906
transform 1 0 263984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_434
timestamp 1698175906
transform 1 0 271824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_435
timestamp 1698175906
transform 1 0 279664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_436
timestamp 1698175906
transform 1 0 287504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_437
timestamp 1698175906
transform 1 0 295344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_438
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_439
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_440
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_441
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_442
timestamp 1698175906
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_443
timestamp 1698175906
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_444
timestamp 1698175906
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_445
timestamp 1698175906
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_446
timestamp 1698175906
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_447
timestamp 1698175906
transform 1 0 79744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_448
timestamp 1698175906
transform 1 0 87584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_449
timestamp 1698175906
transform 1 0 95424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_450
timestamp 1698175906
transform 1 0 103264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_451
timestamp 1698175906
transform 1 0 111104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_452
timestamp 1698175906
transform 1 0 118944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_453
timestamp 1698175906
transform 1 0 126784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_454
timestamp 1698175906
transform 1 0 134624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_455
timestamp 1698175906
transform 1 0 142464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_456
timestamp 1698175906
transform 1 0 150304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_457
timestamp 1698175906
transform 1 0 158144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_458
timestamp 1698175906
transform 1 0 165984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_459
timestamp 1698175906
transform 1 0 173824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_460
timestamp 1698175906
transform 1 0 181664 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_461
timestamp 1698175906
transform 1 0 189504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_462
timestamp 1698175906
transform 1 0 197344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_463
timestamp 1698175906
transform 1 0 205184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_464
timestamp 1698175906
transform 1 0 213024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_465
timestamp 1698175906
transform 1 0 220864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_466
timestamp 1698175906
transform 1 0 228704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_467
timestamp 1698175906
transform 1 0 236544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_468
timestamp 1698175906
transform 1 0 244384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_469
timestamp 1698175906
transform 1 0 252224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_470
timestamp 1698175906
transform 1 0 260064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_471
timestamp 1698175906
transform 1 0 267904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_472
timestamp 1698175906
transform 1 0 275744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_473
timestamp 1698175906
transform 1 0 283584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_474
timestamp 1698175906
transform 1 0 291424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_475
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_476
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_477
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_478
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_479
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_480
timestamp 1698175906
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_481
timestamp 1698175906
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_482
timestamp 1698175906
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_483
timestamp 1698175906
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_484
timestamp 1698175906
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_485
timestamp 1698175906
transform 1 0 83664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_486
timestamp 1698175906
transform 1 0 91504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_487
timestamp 1698175906
transform 1 0 99344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_488
timestamp 1698175906
transform 1 0 107184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_489
timestamp 1698175906
transform 1 0 115024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_490
timestamp 1698175906
transform 1 0 122864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_491
timestamp 1698175906
transform 1 0 130704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_492
timestamp 1698175906
transform 1 0 138544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_493
timestamp 1698175906
transform 1 0 146384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_494
timestamp 1698175906
transform 1 0 154224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_495
timestamp 1698175906
transform 1 0 162064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_496
timestamp 1698175906
transform 1 0 169904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_497
timestamp 1698175906
transform 1 0 177744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_498
timestamp 1698175906
transform 1 0 185584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_499
timestamp 1698175906
transform 1 0 193424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_500
timestamp 1698175906
transform 1 0 201264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_501
timestamp 1698175906
transform 1 0 209104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_502
timestamp 1698175906
transform 1 0 216944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_503
timestamp 1698175906
transform 1 0 224784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_504
timestamp 1698175906
transform 1 0 232624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_505
timestamp 1698175906
transform 1 0 240464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_506
timestamp 1698175906
transform 1 0 248304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_507
timestamp 1698175906
transform 1 0 256144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_508
timestamp 1698175906
transform 1 0 263984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_509
timestamp 1698175906
transform 1 0 271824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_510
timestamp 1698175906
transform 1 0 279664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_511
timestamp 1698175906
transform 1 0 287504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_512
timestamp 1698175906
transform 1 0 295344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_513
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_514
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_515
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_516
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_517
timestamp 1698175906
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_518
timestamp 1698175906
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_519
timestamp 1698175906
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_520
timestamp 1698175906
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_521
timestamp 1698175906
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_522
timestamp 1698175906
transform 1 0 79744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_523
timestamp 1698175906
transform 1 0 87584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_524
timestamp 1698175906
transform 1 0 95424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_525
timestamp 1698175906
transform 1 0 103264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_526
timestamp 1698175906
transform 1 0 111104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_527
timestamp 1698175906
transform 1 0 118944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_528
timestamp 1698175906
transform 1 0 126784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_529
timestamp 1698175906
transform 1 0 134624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_530
timestamp 1698175906
transform 1 0 142464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_531
timestamp 1698175906
transform 1 0 150304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_532
timestamp 1698175906
transform 1 0 158144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_533
timestamp 1698175906
transform 1 0 165984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_534
timestamp 1698175906
transform 1 0 173824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_535
timestamp 1698175906
transform 1 0 181664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_536
timestamp 1698175906
transform 1 0 189504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_537
timestamp 1698175906
transform 1 0 197344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_538
timestamp 1698175906
transform 1 0 205184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_539
timestamp 1698175906
transform 1 0 213024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_540
timestamp 1698175906
transform 1 0 220864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_541
timestamp 1698175906
transform 1 0 228704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_542
timestamp 1698175906
transform 1 0 236544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_543
timestamp 1698175906
transform 1 0 244384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_544
timestamp 1698175906
transform 1 0 252224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_545
timestamp 1698175906
transform 1 0 260064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_546
timestamp 1698175906
transform 1 0 267904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_547
timestamp 1698175906
transform 1 0 275744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_548
timestamp 1698175906
transform 1 0 283584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_549
timestamp 1698175906
transform 1 0 291424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_550
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_551
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_552
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_553
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_554
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_555
timestamp 1698175906
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_556
timestamp 1698175906
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_557
timestamp 1698175906
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_558
timestamp 1698175906
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_559
timestamp 1698175906
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_560
timestamp 1698175906
transform 1 0 83664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_561
timestamp 1698175906
transform 1 0 91504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_562
timestamp 1698175906
transform 1 0 99344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_563
timestamp 1698175906
transform 1 0 107184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_564
timestamp 1698175906
transform 1 0 115024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_565
timestamp 1698175906
transform 1 0 122864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_566
timestamp 1698175906
transform 1 0 130704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_567
timestamp 1698175906
transform 1 0 138544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_568
timestamp 1698175906
transform 1 0 146384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_569
timestamp 1698175906
transform 1 0 154224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_570
timestamp 1698175906
transform 1 0 162064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_571
timestamp 1698175906
transform 1 0 169904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_572
timestamp 1698175906
transform 1 0 177744 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_573
timestamp 1698175906
transform 1 0 185584 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_574
timestamp 1698175906
transform 1 0 193424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_575
timestamp 1698175906
transform 1 0 201264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_576
timestamp 1698175906
transform 1 0 209104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_577
timestamp 1698175906
transform 1 0 216944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_578
timestamp 1698175906
transform 1 0 224784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_579
timestamp 1698175906
transform 1 0 232624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_580
timestamp 1698175906
transform 1 0 240464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_581
timestamp 1698175906
transform 1 0 248304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_582
timestamp 1698175906
transform 1 0 256144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_583
timestamp 1698175906
transform 1 0 263984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_584
timestamp 1698175906
transform 1 0 271824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_585
timestamp 1698175906
transform 1 0 279664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_586
timestamp 1698175906
transform 1 0 287504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_587
timestamp 1698175906
transform 1 0 295344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_588
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_589
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_590
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_591
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_592
timestamp 1698175906
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_593
timestamp 1698175906
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_594
timestamp 1698175906
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_595
timestamp 1698175906
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_596
timestamp 1698175906
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_597
timestamp 1698175906
transform 1 0 79744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_598
timestamp 1698175906
transform 1 0 87584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_599
timestamp 1698175906
transform 1 0 95424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_600
timestamp 1698175906
transform 1 0 103264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_601
timestamp 1698175906
transform 1 0 111104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_602
timestamp 1698175906
transform 1 0 118944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_603
timestamp 1698175906
transform 1 0 126784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_604
timestamp 1698175906
transform 1 0 134624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_605
timestamp 1698175906
transform 1 0 142464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_606
timestamp 1698175906
transform 1 0 150304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_607
timestamp 1698175906
transform 1 0 158144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_608
timestamp 1698175906
transform 1 0 165984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_609
timestamp 1698175906
transform 1 0 173824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_610
timestamp 1698175906
transform 1 0 181664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_611
timestamp 1698175906
transform 1 0 189504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_612
timestamp 1698175906
transform 1 0 197344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_613
timestamp 1698175906
transform 1 0 205184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_614
timestamp 1698175906
transform 1 0 213024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_615
timestamp 1698175906
transform 1 0 220864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_616
timestamp 1698175906
transform 1 0 228704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_617
timestamp 1698175906
transform 1 0 236544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_618
timestamp 1698175906
transform 1 0 244384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_619
timestamp 1698175906
transform 1 0 252224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_620
timestamp 1698175906
transform 1 0 260064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_621
timestamp 1698175906
transform 1 0 267904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_622
timestamp 1698175906
transform 1 0 275744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_623
timestamp 1698175906
transform 1 0 283584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_624
timestamp 1698175906
transform 1 0 291424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_625
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_626
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_627
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_628
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_629
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_630
timestamp 1698175906
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_631
timestamp 1698175906
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_632
timestamp 1698175906
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_633
timestamp 1698175906
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_634
timestamp 1698175906
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_635
timestamp 1698175906
transform 1 0 83664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_636
timestamp 1698175906
transform 1 0 91504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_637
timestamp 1698175906
transform 1 0 99344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_638
timestamp 1698175906
transform 1 0 107184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_639
timestamp 1698175906
transform 1 0 115024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_640
timestamp 1698175906
transform 1 0 122864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_641
timestamp 1698175906
transform 1 0 130704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_642
timestamp 1698175906
transform 1 0 138544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_643
timestamp 1698175906
transform 1 0 146384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_644
timestamp 1698175906
transform 1 0 154224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_645
timestamp 1698175906
transform 1 0 162064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_646
timestamp 1698175906
transform 1 0 169904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_647
timestamp 1698175906
transform 1 0 177744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_648
timestamp 1698175906
transform 1 0 185584 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_649
timestamp 1698175906
transform 1 0 193424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_650
timestamp 1698175906
transform 1 0 201264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_651
timestamp 1698175906
transform 1 0 209104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_652
timestamp 1698175906
transform 1 0 216944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_653
timestamp 1698175906
transform 1 0 224784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_654
timestamp 1698175906
transform 1 0 232624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_655
timestamp 1698175906
transform 1 0 240464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_656
timestamp 1698175906
transform 1 0 248304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_657
timestamp 1698175906
transform 1 0 256144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_658
timestamp 1698175906
transform 1 0 263984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_659
timestamp 1698175906
transform 1 0 271824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_660
timestamp 1698175906
transform 1 0 279664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_661
timestamp 1698175906
transform 1 0 287504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_662
timestamp 1698175906
transform 1 0 295344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_663
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_664
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_665
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_666
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_667
timestamp 1698175906
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_668
timestamp 1698175906
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_669
timestamp 1698175906
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_670
timestamp 1698175906
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_671
timestamp 1698175906
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_672
timestamp 1698175906
transform 1 0 79744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_673
timestamp 1698175906
transform 1 0 87584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_674
timestamp 1698175906
transform 1 0 95424 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_675
timestamp 1698175906
transform 1 0 103264 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_676
timestamp 1698175906
transform 1 0 111104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_677
timestamp 1698175906
transform 1 0 118944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_678
timestamp 1698175906
transform 1 0 126784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_679
timestamp 1698175906
transform 1 0 134624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_680
timestamp 1698175906
transform 1 0 142464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_681
timestamp 1698175906
transform 1 0 150304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_682
timestamp 1698175906
transform 1 0 158144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_683
timestamp 1698175906
transform 1 0 165984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_684
timestamp 1698175906
transform 1 0 173824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_685
timestamp 1698175906
transform 1 0 181664 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_686
timestamp 1698175906
transform 1 0 189504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_687
timestamp 1698175906
transform 1 0 197344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_688
timestamp 1698175906
transform 1 0 205184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_689
timestamp 1698175906
transform 1 0 213024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_690
timestamp 1698175906
transform 1 0 220864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_691
timestamp 1698175906
transform 1 0 228704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_692
timestamp 1698175906
transform 1 0 236544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_693
timestamp 1698175906
transform 1 0 244384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_694
timestamp 1698175906
transform 1 0 252224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_695
timestamp 1698175906
transform 1 0 260064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_696
timestamp 1698175906
transform 1 0 267904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_697
timestamp 1698175906
transform 1 0 275744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_698
timestamp 1698175906
transform 1 0 283584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_699
timestamp 1698175906
transform 1 0 291424 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_700
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_701
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_702
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_703
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_704
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_705
timestamp 1698175906
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_706
timestamp 1698175906
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_707
timestamp 1698175906
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_708
timestamp 1698175906
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_709
timestamp 1698175906
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_710
timestamp 1698175906
transform 1 0 83664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_711
timestamp 1698175906
transform 1 0 91504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_712
timestamp 1698175906
transform 1 0 99344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_713
timestamp 1698175906
transform 1 0 107184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_714
timestamp 1698175906
transform 1 0 115024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_715
timestamp 1698175906
transform 1 0 122864 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_716
timestamp 1698175906
transform 1 0 130704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_717
timestamp 1698175906
transform 1 0 138544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_718
timestamp 1698175906
transform 1 0 146384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_719
timestamp 1698175906
transform 1 0 154224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_720
timestamp 1698175906
transform 1 0 162064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_721
timestamp 1698175906
transform 1 0 169904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_722
timestamp 1698175906
transform 1 0 177744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_723
timestamp 1698175906
transform 1 0 185584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_724
timestamp 1698175906
transform 1 0 193424 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_725
timestamp 1698175906
transform 1 0 201264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_726
timestamp 1698175906
transform 1 0 209104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_727
timestamp 1698175906
transform 1 0 216944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_728
timestamp 1698175906
transform 1 0 224784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_729
timestamp 1698175906
transform 1 0 232624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_730
timestamp 1698175906
transform 1 0 240464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_731
timestamp 1698175906
transform 1 0 248304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_732
timestamp 1698175906
transform 1 0 256144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_733
timestamp 1698175906
transform 1 0 263984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_734
timestamp 1698175906
transform 1 0 271824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_735
timestamp 1698175906
transform 1 0 279664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_736
timestamp 1698175906
transform 1 0 287504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_737
timestamp 1698175906
transform 1 0 295344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_738
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_739
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_740
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_741
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_742
timestamp 1698175906
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_743
timestamp 1698175906
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_744
timestamp 1698175906
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_745
timestamp 1698175906
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_746
timestamp 1698175906
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_747
timestamp 1698175906
transform 1 0 79744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_748
timestamp 1698175906
transform 1 0 87584 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_749
timestamp 1698175906
transform 1 0 95424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_750
timestamp 1698175906
transform 1 0 103264 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_751
timestamp 1698175906
transform 1 0 111104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_752
timestamp 1698175906
transform 1 0 118944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_753
timestamp 1698175906
transform 1 0 126784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_754
timestamp 1698175906
transform 1 0 134624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_755
timestamp 1698175906
transform 1 0 142464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_756
timestamp 1698175906
transform 1 0 150304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_757
timestamp 1698175906
transform 1 0 158144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_758
timestamp 1698175906
transform 1 0 165984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_759
timestamp 1698175906
transform 1 0 173824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_760
timestamp 1698175906
transform 1 0 181664 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_761
timestamp 1698175906
transform 1 0 189504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_762
timestamp 1698175906
transform 1 0 197344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_763
timestamp 1698175906
transform 1 0 205184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_764
timestamp 1698175906
transform 1 0 213024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_765
timestamp 1698175906
transform 1 0 220864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_766
timestamp 1698175906
transform 1 0 228704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_767
timestamp 1698175906
transform 1 0 236544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_768
timestamp 1698175906
transform 1 0 244384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_769
timestamp 1698175906
transform 1 0 252224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_770
timestamp 1698175906
transform 1 0 260064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_771
timestamp 1698175906
transform 1 0 267904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_772
timestamp 1698175906
transform 1 0 275744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_773
timestamp 1698175906
transform 1 0 283584 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_774
timestamp 1698175906
transform 1 0 291424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_775
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_776
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_777
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_778
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_779
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_780
timestamp 1698175906
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_781
timestamp 1698175906
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_782
timestamp 1698175906
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_783
timestamp 1698175906
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_784
timestamp 1698175906
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_785
timestamp 1698175906
transform 1 0 83664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_786
timestamp 1698175906
transform 1 0 91504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_787
timestamp 1698175906
transform 1 0 99344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_788
timestamp 1698175906
transform 1 0 107184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_789
timestamp 1698175906
transform 1 0 115024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_790
timestamp 1698175906
transform 1 0 122864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_791
timestamp 1698175906
transform 1 0 130704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_792
timestamp 1698175906
transform 1 0 138544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_793
timestamp 1698175906
transform 1 0 146384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_794
timestamp 1698175906
transform 1 0 154224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_795
timestamp 1698175906
transform 1 0 162064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_796
timestamp 1698175906
transform 1 0 169904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_797
timestamp 1698175906
transform 1 0 177744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_798
timestamp 1698175906
transform 1 0 185584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_799
timestamp 1698175906
transform 1 0 193424 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_800
timestamp 1698175906
transform 1 0 201264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_801
timestamp 1698175906
transform 1 0 209104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_802
timestamp 1698175906
transform 1 0 216944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_803
timestamp 1698175906
transform 1 0 224784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_804
timestamp 1698175906
transform 1 0 232624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_805
timestamp 1698175906
transform 1 0 240464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_806
timestamp 1698175906
transform 1 0 248304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_807
timestamp 1698175906
transform 1 0 256144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_808
timestamp 1698175906
transform 1 0 263984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_809
timestamp 1698175906
transform 1 0 271824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_810
timestamp 1698175906
transform 1 0 279664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_811
timestamp 1698175906
transform 1 0 287504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_812
timestamp 1698175906
transform 1 0 295344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_813
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_814
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_815
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_816
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_817
timestamp 1698175906
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_818
timestamp 1698175906
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_819
timestamp 1698175906
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_820
timestamp 1698175906
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_821
timestamp 1698175906
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_822
timestamp 1698175906
transform 1 0 79744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_823
timestamp 1698175906
transform 1 0 87584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_824
timestamp 1698175906
transform 1 0 95424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_825
timestamp 1698175906
transform 1 0 103264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_826
timestamp 1698175906
transform 1 0 111104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_827
timestamp 1698175906
transform 1 0 118944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_828
timestamp 1698175906
transform 1 0 126784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_829
timestamp 1698175906
transform 1 0 134624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_830
timestamp 1698175906
transform 1 0 142464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_831
timestamp 1698175906
transform 1 0 150304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_832
timestamp 1698175906
transform 1 0 158144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_833
timestamp 1698175906
transform 1 0 165984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_834
timestamp 1698175906
transform 1 0 173824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_835
timestamp 1698175906
transform 1 0 181664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_836
timestamp 1698175906
transform 1 0 189504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_837
timestamp 1698175906
transform 1 0 197344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_838
timestamp 1698175906
transform 1 0 205184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_839
timestamp 1698175906
transform 1 0 213024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_840
timestamp 1698175906
transform 1 0 220864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_841
timestamp 1698175906
transform 1 0 228704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_842
timestamp 1698175906
transform 1 0 236544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_843
timestamp 1698175906
transform 1 0 244384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_844
timestamp 1698175906
transform 1 0 252224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_845
timestamp 1698175906
transform 1 0 260064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_846
timestamp 1698175906
transform 1 0 267904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_847
timestamp 1698175906
transform 1 0 275744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_848
timestamp 1698175906
transform 1 0 283584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_849
timestamp 1698175906
transform 1 0 291424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_850
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_851
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_852
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_853
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_854
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_855
timestamp 1698175906
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_856
timestamp 1698175906
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_857
timestamp 1698175906
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_858
timestamp 1698175906
transform 1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_859
timestamp 1698175906
transform 1 0 75824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_860
timestamp 1698175906
transform 1 0 83664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_861
timestamp 1698175906
transform 1 0 91504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_862
timestamp 1698175906
transform 1 0 99344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_863
timestamp 1698175906
transform 1 0 107184 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_864
timestamp 1698175906
transform 1 0 115024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_865
timestamp 1698175906
transform 1 0 122864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_866
timestamp 1698175906
transform 1 0 130704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_867
timestamp 1698175906
transform 1 0 138544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_868
timestamp 1698175906
transform 1 0 146384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_869
timestamp 1698175906
transform 1 0 154224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_870
timestamp 1698175906
transform 1 0 162064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_871
timestamp 1698175906
transform 1 0 169904 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_872
timestamp 1698175906
transform 1 0 177744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_873
timestamp 1698175906
transform 1 0 185584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_874
timestamp 1698175906
transform 1 0 193424 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_875
timestamp 1698175906
transform 1 0 201264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_876
timestamp 1698175906
transform 1 0 209104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_877
timestamp 1698175906
transform 1 0 216944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_878
timestamp 1698175906
transform 1 0 224784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_879
timestamp 1698175906
transform 1 0 232624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_880
timestamp 1698175906
transform 1 0 240464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_881
timestamp 1698175906
transform 1 0 248304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_882
timestamp 1698175906
transform 1 0 256144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_883
timestamp 1698175906
transform 1 0 263984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_884
timestamp 1698175906
transform 1 0 271824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_885
timestamp 1698175906
transform 1 0 279664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_886
timestamp 1698175906
transform 1 0 287504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_887
timestamp 1698175906
transform 1 0 295344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_888
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_889
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_890
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_891
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_892
timestamp 1698175906
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_893
timestamp 1698175906
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_894
timestamp 1698175906
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_895
timestamp 1698175906
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_896
timestamp 1698175906
transform 1 0 71904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_897
timestamp 1698175906
transform 1 0 79744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_898
timestamp 1698175906
transform 1 0 87584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_899
timestamp 1698175906
transform 1 0 95424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_900
timestamp 1698175906
transform 1 0 103264 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_901
timestamp 1698175906
transform 1 0 111104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_902
timestamp 1698175906
transform 1 0 118944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_903
timestamp 1698175906
transform 1 0 126784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_904
timestamp 1698175906
transform 1 0 134624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_905
timestamp 1698175906
transform 1 0 142464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_906
timestamp 1698175906
transform 1 0 150304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_907
timestamp 1698175906
transform 1 0 158144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_908
timestamp 1698175906
transform 1 0 165984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_909
timestamp 1698175906
transform 1 0 173824 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_910
timestamp 1698175906
transform 1 0 181664 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_911
timestamp 1698175906
transform 1 0 189504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_912
timestamp 1698175906
transform 1 0 197344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_913
timestamp 1698175906
transform 1 0 205184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_914
timestamp 1698175906
transform 1 0 213024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_915
timestamp 1698175906
transform 1 0 220864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_916
timestamp 1698175906
transform 1 0 228704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_917
timestamp 1698175906
transform 1 0 236544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_918
timestamp 1698175906
transform 1 0 244384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_919
timestamp 1698175906
transform 1 0 252224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_920
timestamp 1698175906
transform 1 0 260064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_921
timestamp 1698175906
transform 1 0 267904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_922
timestamp 1698175906
transform 1 0 275744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_923
timestamp 1698175906
transform 1 0 283584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_924
timestamp 1698175906
transform 1 0 291424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_925
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_926
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_927
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_928
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_929
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_930
timestamp 1698175906
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_931
timestamp 1698175906
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_932
timestamp 1698175906
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_933
timestamp 1698175906
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_934
timestamp 1698175906
transform 1 0 75824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_935
timestamp 1698175906
transform 1 0 83664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_936
timestamp 1698175906
transform 1 0 91504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_937
timestamp 1698175906
transform 1 0 99344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_938
timestamp 1698175906
transform 1 0 107184 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_939
timestamp 1698175906
transform 1 0 115024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_940
timestamp 1698175906
transform 1 0 122864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_941
timestamp 1698175906
transform 1 0 130704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_942
timestamp 1698175906
transform 1 0 138544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_943
timestamp 1698175906
transform 1 0 146384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_944
timestamp 1698175906
transform 1 0 154224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_945
timestamp 1698175906
transform 1 0 162064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_946
timestamp 1698175906
transform 1 0 169904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_947
timestamp 1698175906
transform 1 0 177744 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_948
timestamp 1698175906
transform 1 0 185584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_949
timestamp 1698175906
transform 1 0 193424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_950
timestamp 1698175906
transform 1 0 201264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_951
timestamp 1698175906
transform 1 0 209104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_952
timestamp 1698175906
transform 1 0 216944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_953
timestamp 1698175906
transform 1 0 224784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_954
timestamp 1698175906
transform 1 0 232624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_955
timestamp 1698175906
transform 1 0 240464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_956
timestamp 1698175906
transform 1 0 248304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_957
timestamp 1698175906
transform 1 0 256144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_958
timestamp 1698175906
transform 1 0 263984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_959
timestamp 1698175906
transform 1 0 271824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_960
timestamp 1698175906
transform 1 0 279664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_961
timestamp 1698175906
transform 1 0 287504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_962
timestamp 1698175906
transform 1 0 295344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_963
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_964
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_965
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_966
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_967
timestamp 1698175906
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_968
timestamp 1698175906
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_969
timestamp 1698175906
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_970
timestamp 1698175906
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_971
timestamp 1698175906
transform 1 0 71904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_972
timestamp 1698175906
transform 1 0 79744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_973
timestamp 1698175906
transform 1 0 87584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_974
timestamp 1698175906
transform 1 0 95424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_975
timestamp 1698175906
transform 1 0 103264 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_976
timestamp 1698175906
transform 1 0 111104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_977
timestamp 1698175906
transform 1 0 118944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_978
timestamp 1698175906
transform 1 0 126784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_979
timestamp 1698175906
transform 1 0 134624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_980
timestamp 1698175906
transform 1 0 142464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_981
timestamp 1698175906
transform 1 0 150304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_982
timestamp 1698175906
transform 1 0 158144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_983
timestamp 1698175906
transform 1 0 165984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_984
timestamp 1698175906
transform 1 0 173824 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_985
timestamp 1698175906
transform 1 0 181664 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_986
timestamp 1698175906
transform 1 0 189504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_987
timestamp 1698175906
transform 1 0 197344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_988
timestamp 1698175906
transform 1 0 205184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_989
timestamp 1698175906
transform 1 0 213024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_990
timestamp 1698175906
transform 1 0 220864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_991
timestamp 1698175906
transform 1 0 228704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_992
timestamp 1698175906
transform 1 0 236544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_993
timestamp 1698175906
transform 1 0 244384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_994
timestamp 1698175906
transform 1 0 252224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_995
timestamp 1698175906
transform 1 0 260064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_996
timestamp 1698175906
transform 1 0 267904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_997
timestamp 1698175906
transform 1 0 275744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_998
timestamp 1698175906
transform 1 0 283584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_999
timestamp 1698175906
transform 1 0 291424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1000
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1001
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1002
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1003
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1004
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1005
timestamp 1698175906
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1006
timestamp 1698175906
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1007
timestamp 1698175906
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1008
timestamp 1698175906
transform 1 0 67984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1009
timestamp 1698175906
transform 1 0 75824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1010
timestamp 1698175906
transform 1 0 83664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1011
timestamp 1698175906
transform 1 0 91504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1012
timestamp 1698175906
transform 1 0 99344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1013
timestamp 1698175906
transform 1 0 107184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1014
timestamp 1698175906
transform 1 0 115024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1015
timestamp 1698175906
transform 1 0 122864 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1016
timestamp 1698175906
transform 1 0 130704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1017
timestamp 1698175906
transform 1 0 138544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1018
timestamp 1698175906
transform 1 0 146384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1019
timestamp 1698175906
transform 1 0 154224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1020
timestamp 1698175906
transform 1 0 162064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1021
timestamp 1698175906
transform 1 0 169904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1022
timestamp 1698175906
transform 1 0 177744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1023
timestamp 1698175906
transform 1 0 185584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1024
timestamp 1698175906
transform 1 0 193424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1025
timestamp 1698175906
transform 1 0 201264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1026
timestamp 1698175906
transform 1 0 209104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1027
timestamp 1698175906
transform 1 0 216944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1028
timestamp 1698175906
transform 1 0 224784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1029
timestamp 1698175906
transform 1 0 232624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1030
timestamp 1698175906
transform 1 0 240464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1031
timestamp 1698175906
transform 1 0 248304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1032
timestamp 1698175906
transform 1 0 256144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1033
timestamp 1698175906
transform 1 0 263984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1034
timestamp 1698175906
transform 1 0 271824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1035
timestamp 1698175906
transform 1 0 279664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1036
timestamp 1698175906
transform 1 0 287504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1037
timestamp 1698175906
transform 1 0 295344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1038
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1039
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1040
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1041
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1042
timestamp 1698175906
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1043
timestamp 1698175906
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1044
timestamp 1698175906
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1045
timestamp 1698175906
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1046
timestamp 1698175906
transform 1 0 71904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1047
timestamp 1698175906
transform 1 0 79744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1048
timestamp 1698175906
transform 1 0 87584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1049
timestamp 1698175906
transform 1 0 95424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1050
timestamp 1698175906
transform 1 0 103264 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1051
timestamp 1698175906
transform 1 0 111104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1052
timestamp 1698175906
transform 1 0 118944 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1053
timestamp 1698175906
transform 1 0 126784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1054
timestamp 1698175906
transform 1 0 134624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1055
timestamp 1698175906
transform 1 0 142464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1056
timestamp 1698175906
transform 1 0 150304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1057
timestamp 1698175906
transform 1 0 158144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1058
timestamp 1698175906
transform 1 0 165984 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1059
timestamp 1698175906
transform 1 0 173824 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1060
timestamp 1698175906
transform 1 0 181664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1061
timestamp 1698175906
transform 1 0 189504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1062
timestamp 1698175906
transform 1 0 197344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1063
timestamp 1698175906
transform 1 0 205184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1064
timestamp 1698175906
transform 1 0 213024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1065
timestamp 1698175906
transform 1 0 220864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1066
timestamp 1698175906
transform 1 0 228704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1067
timestamp 1698175906
transform 1 0 236544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1068
timestamp 1698175906
transform 1 0 244384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1069
timestamp 1698175906
transform 1 0 252224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1070
timestamp 1698175906
transform 1 0 260064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1071
timestamp 1698175906
transform 1 0 267904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1072
timestamp 1698175906
transform 1 0 275744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1073
timestamp 1698175906
transform 1 0 283584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1074
timestamp 1698175906
transform 1 0 291424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1075
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1076
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1077
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1078
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1079
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1080
timestamp 1698175906
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1081
timestamp 1698175906
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1082
timestamp 1698175906
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1083
timestamp 1698175906
transform 1 0 67984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1084
timestamp 1698175906
transform 1 0 75824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1085
timestamp 1698175906
transform 1 0 83664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1086
timestamp 1698175906
transform 1 0 91504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1087
timestamp 1698175906
transform 1 0 99344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1088
timestamp 1698175906
transform 1 0 107184 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1089
timestamp 1698175906
transform 1 0 115024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1090
timestamp 1698175906
transform 1 0 122864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1091
timestamp 1698175906
transform 1 0 130704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1092
timestamp 1698175906
transform 1 0 138544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1093
timestamp 1698175906
transform 1 0 146384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1094
timestamp 1698175906
transform 1 0 154224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1095
timestamp 1698175906
transform 1 0 162064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1096
timestamp 1698175906
transform 1 0 169904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1097
timestamp 1698175906
transform 1 0 177744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1098
timestamp 1698175906
transform 1 0 185584 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1099
timestamp 1698175906
transform 1 0 193424 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1100
timestamp 1698175906
transform 1 0 201264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1101
timestamp 1698175906
transform 1 0 209104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1102
timestamp 1698175906
transform 1 0 216944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1103
timestamp 1698175906
transform 1 0 224784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1104
timestamp 1698175906
transform 1 0 232624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1105
timestamp 1698175906
transform 1 0 240464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1106
timestamp 1698175906
transform 1 0 248304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1107
timestamp 1698175906
transform 1 0 256144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1108
timestamp 1698175906
transform 1 0 263984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1109
timestamp 1698175906
transform 1 0 271824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1110
timestamp 1698175906
transform 1 0 279664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1111
timestamp 1698175906
transform 1 0 287504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1112
timestamp 1698175906
transform 1 0 295344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1113
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1114
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1115
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1116
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1117
timestamp 1698175906
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1118
timestamp 1698175906
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1119
timestamp 1698175906
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1120
timestamp 1698175906
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1121
timestamp 1698175906
transform 1 0 71904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1122
timestamp 1698175906
transform 1 0 79744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1123
timestamp 1698175906
transform 1 0 87584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1124
timestamp 1698175906
transform 1 0 95424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1125
timestamp 1698175906
transform 1 0 103264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1126
timestamp 1698175906
transform 1 0 111104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1127
timestamp 1698175906
transform 1 0 118944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1128
timestamp 1698175906
transform 1 0 126784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1129
timestamp 1698175906
transform 1 0 134624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1130
timestamp 1698175906
transform 1 0 142464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1131
timestamp 1698175906
transform 1 0 150304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1132
timestamp 1698175906
transform 1 0 158144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1133
timestamp 1698175906
transform 1 0 165984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1134
timestamp 1698175906
transform 1 0 173824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1135
timestamp 1698175906
transform 1 0 181664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1136
timestamp 1698175906
transform 1 0 189504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1137
timestamp 1698175906
transform 1 0 197344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1138
timestamp 1698175906
transform 1 0 205184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1139
timestamp 1698175906
transform 1 0 213024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1140
timestamp 1698175906
transform 1 0 220864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1141
timestamp 1698175906
transform 1 0 228704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1142
timestamp 1698175906
transform 1 0 236544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1143
timestamp 1698175906
transform 1 0 244384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1144
timestamp 1698175906
transform 1 0 252224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1145
timestamp 1698175906
transform 1 0 260064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1146
timestamp 1698175906
transform 1 0 267904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1147
timestamp 1698175906
transform 1 0 275744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1148
timestamp 1698175906
transform 1 0 283584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1149
timestamp 1698175906
transform 1 0 291424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1150
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1151
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1152
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1153
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1154
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1155
timestamp 1698175906
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1156
timestamp 1698175906
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1157
timestamp 1698175906
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1158
timestamp 1698175906
transform 1 0 67984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1159
timestamp 1698175906
transform 1 0 75824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1160
timestamp 1698175906
transform 1 0 83664 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1161
timestamp 1698175906
transform 1 0 91504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1162
timestamp 1698175906
transform 1 0 99344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1163
timestamp 1698175906
transform 1 0 107184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1164
timestamp 1698175906
transform 1 0 115024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1165
timestamp 1698175906
transform 1 0 122864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1166
timestamp 1698175906
transform 1 0 130704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1167
timestamp 1698175906
transform 1 0 138544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1168
timestamp 1698175906
transform 1 0 146384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1169
timestamp 1698175906
transform 1 0 154224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1170
timestamp 1698175906
transform 1 0 162064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1171
timestamp 1698175906
transform 1 0 169904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1172
timestamp 1698175906
transform 1 0 177744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1173
timestamp 1698175906
transform 1 0 185584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1174
timestamp 1698175906
transform 1 0 193424 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1175
timestamp 1698175906
transform 1 0 201264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1176
timestamp 1698175906
transform 1 0 209104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1177
timestamp 1698175906
transform 1 0 216944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1178
timestamp 1698175906
transform 1 0 224784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1179
timestamp 1698175906
transform 1 0 232624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1180
timestamp 1698175906
transform 1 0 240464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1181
timestamp 1698175906
transform 1 0 248304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1182
timestamp 1698175906
transform 1 0 256144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1183
timestamp 1698175906
transform 1 0 263984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1184
timestamp 1698175906
transform 1 0 271824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1185
timestamp 1698175906
transform 1 0 279664 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1186
timestamp 1698175906
transform 1 0 287504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1187
timestamp 1698175906
transform 1 0 295344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1188
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1189
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1190
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1191
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1192
timestamp 1698175906
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1193
timestamp 1698175906
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1194
timestamp 1698175906
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1195
timestamp 1698175906
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1196
timestamp 1698175906
transform 1 0 71904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1197
timestamp 1698175906
transform 1 0 79744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1198
timestamp 1698175906
transform 1 0 87584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1199
timestamp 1698175906
transform 1 0 95424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1200
timestamp 1698175906
transform 1 0 103264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1201
timestamp 1698175906
transform 1 0 111104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1202
timestamp 1698175906
transform 1 0 118944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1203
timestamp 1698175906
transform 1 0 126784 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1204
timestamp 1698175906
transform 1 0 134624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1205
timestamp 1698175906
transform 1 0 142464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1206
timestamp 1698175906
transform 1 0 150304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1207
timestamp 1698175906
transform 1 0 158144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1208
timestamp 1698175906
transform 1 0 165984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1209
timestamp 1698175906
transform 1 0 173824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1210
timestamp 1698175906
transform 1 0 181664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1211
timestamp 1698175906
transform 1 0 189504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1212
timestamp 1698175906
transform 1 0 197344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1213
timestamp 1698175906
transform 1 0 205184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1214
timestamp 1698175906
transform 1 0 213024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1215
timestamp 1698175906
transform 1 0 220864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1216
timestamp 1698175906
transform 1 0 228704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1217
timestamp 1698175906
transform 1 0 236544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1218
timestamp 1698175906
transform 1 0 244384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1219
timestamp 1698175906
transform 1 0 252224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1220
timestamp 1698175906
transform 1 0 260064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1221
timestamp 1698175906
transform 1 0 267904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1222
timestamp 1698175906
transform 1 0 275744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1223
timestamp 1698175906
transform 1 0 283584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1224
timestamp 1698175906
transform 1 0 291424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1225
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1226
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1227
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1228
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1229
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1230
timestamp 1698175906
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1231
timestamp 1698175906
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1232
timestamp 1698175906
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1233
timestamp 1698175906
transform 1 0 67984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1234
timestamp 1698175906
transform 1 0 75824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1235
timestamp 1698175906
transform 1 0 83664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1236
timestamp 1698175906
transform 1 0 91504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1237
timestamp 1698175906
transform 1 0 99344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1238
timestamp 1698175906
transform 1 0 107184 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1239
timestamp 1698175906
transform 1 0 115024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1240
timestamp 1698175906
transform 1 0 122864 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1241
timestamp 1698175906
transform 1 0 130704 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1242
timestamp 1698175906
transform 1 0 138544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1243
timestamp 1698175906
transform 1 0 146384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1244
timestamp 1698175906
transform 1 0 154224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1245
timestamp 1698175906
transform 1 0 162064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1246
timestamp 1698175906
transform 1 0 169904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1247
timestamp 1698175906
transform 1 0 177744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1248
timestamp 1698175906
transform 1 0 185584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1249
timestamp 1698175906
transform 1 0 193424 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1250
timestamp 1698175906
transform 1 0 201264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1251
timestamp 1698175906
transform 1 0 209104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1252
timestamp 1698175906
transform 1 0 216944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1253
timestamp 1698175906
transform 1 0 224784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1254
timestamp 1698175906
transform 1 0 232624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1255
timestamp 1698175906
transform 1 0 240464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1256
timestamp 1698175906
transform 1 0 248304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1257
timestamp 1698175906
transform 1 0 256144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1258
timestamp 1698175906
transform 1 0 263984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1259
timestamp 1698175906
transform 1 0 271824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1260
timestamp 1698175906
transform 1 0 279664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1261
timestamp 1698175906
transform 1 0 287504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1262
timestamp 1698175906
transform 1 0 295344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1263
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1264
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1265
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1266
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1267
timestamp 1698175906
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1268
timestamp 1698175906
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1269
timestamp 1698175906
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1270
timestamp 1698175906
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1271
timestamp 1698175906
transform 1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1272
timestamp 1698175906
transform 1 0 79744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1273
timestamp 1698175906
transform 1 0 87584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1274
timestamp 1698175906
transform 1 0 95424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1275
timestamp 1698175906
transform 1 0 103264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1276
timestamp 1698175906
transform 1 0 111104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1277
timestamp 1698175906
transform 1 0 118944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1278
timestamp 1698175906
transform 1 0 126784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1279
timestamp 1698175906
transform 1 0 134624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1280
timestamp 1698175906
transform 1 0 142464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1281
timestamp 1698175906
transform 1 0 150304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1282
timestamp 1698175906
transform 1 0 158144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1283
timestamp 1698175906
transform 1 0 165984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1284
timestamp 1698175906
transform 1 0 173824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1285
timestamp 1698175906
transform 1 0 181664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1286
timestamp 1698175906
transform 1 0 189504 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1287
timestamp 1698175906
transform 1 0 197344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1288
timestamp 1698175906
transform 1 0 205184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1289
timestamp 1698175906
transform 1 0 213024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1290
timestamp 1698175906
transform 1 0 220864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1291
timestamp 1698175906
transform 1 0 228704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1292
timestamp 1698175906
transform 1 0 236544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1293
timestamp 1698175906
transform 1 0 244384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1294
timestamp 1698175906
transform 1 0 252224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1295
timestamp 1698175906
transform 1 0 260064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1296
timestamp 1698175906
transform 1 0 267904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1297
timestamp 1698175906
transform 1 0 275744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1298
timestamp 1698175906
transform 1 0 283584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1299
timestamp 1698175906
transform 1 0 291424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1300
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1301
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1302
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1303
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1304
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1305
timestamp 1698175906
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1306
timestamp 1698175906
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1307
timestamp 1698175906
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1308
timestamp 1698175906
transform 1 0 67984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1309
timestamp 1698175906
transform 1 0 75824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1310
timestamp 1698175906
transform 1 0 83664 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1311
timestamp 1698175906
transform 1 0 91504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1312
timestamp 1698175906
transform 1 0 99344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1313
timestamp 1698175906
transform 1 0 107184 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1314
timestamp 1698175906
transform 1 0 115024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1315
timestamp 1698175906
transform 1 0 122864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1316
timestamp 1698175906
transform 1 0 130704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1317
timestamp 1698175906
transform 1 0 138544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1318
timestamp 1698175906
transform 1 0 146384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1319
timestamp 1698175906
transform 1 0 154224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1320
timestamp 1698175906
transform 1 0 162064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1321
timestamp 1698175906
transform 1 0 169904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1322
timestamp 1698175906
transform 1 0 177744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1323
timestamp 1698175906
transform 1 0 185584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1324
timestamp 1698175906
transform 1 0 193424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1325
timestamp 1698175906
transform 1 0 201264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1326
timestamp 1698175906
transform 1 0 209104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1327
timestamp 1698175906
transform 1 0 216944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1328
timestamp 1698175906
transform 1 0 224784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1329
timestamp 1698175906
transform 1 0 232624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1330
timestamp 1698175906
transform 1 0 240464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1331
timestamp 1698175906
transform 1 0 248304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1332
timestamp 1698175906
transform 1 0 256144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1333
timestamp 1698175906
transform 1 0 263984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1334
timestamp 1698175906
transform 1 0 271824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1335
timestamp 1698175906
transform 1 0 279664 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1336
timestamp 1698175906
transform 1 0 287504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1337
timestamp 1698175906
transform 1 0 295344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1338
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1339
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1340
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1341
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1342
timestamp 1698175906
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1343
timestamp 1698175906
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1344
timestamp 1698175906
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1345
timestamp 1698175906
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1346
timestamp 1698175906
transform 1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1347
timestamp 1698175906
transform 1 0 79744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1348
timestamp 1698175906
transform 1 0 87584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1349
timestamp 1698175906
transform 1 0 95424 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1350
timestamp 1698175906
transform 1 0 103264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1351
timestamp 1698175906
transform 1 0 111104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1352
timestamp 1698175906
transform 1 0 118944 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1353
timestamp 1698175906
transform 1 0 126784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1354
timestamp 1698175906
transform 1 0 134624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1355
timestamp 1698175906
transform 1 0 142464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1356
timestamp 1698175906
transform 1 0 150304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1357
timestamp 1698175906
transform 1 0 158144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1358
timestamp 1698175906
transform 1 0 165984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1359
timestamp 1698175906
transform 1 0 173824 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1360
timestamp 1698175906
transform 1 0 181664 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1361
timestamp 1698175906
transform 1 0 189504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1362
timestamp 1698175906
transform 1 0 197344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1363
timestamp 1698175906
transform 1 0 205184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1364
timestamp 1698175906
transform 1 0 213024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1365
timestamp 1698175906
transform 1 0 220864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1366
timestamp 1698175906
transform 1 0 228704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1367
timestamp 1698175906
transform 1 0 236544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1368
timestamp 1698175906
transform 1 0 244384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1369
timestamp 1698175906
transform 1 0 252224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1370
timestamp 1698175906
transform 1 0 260064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1371
timestamp 1698175906
transform 1 0 267904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1372
timestamp 1698175906
transform 1 0 275744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1373
timestamp 1698175906
transform 1 0 283584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1374
timestamp 1698175906
transform 1 0 291424 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1375
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1376
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1377
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1378
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1379
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1380
timestamp 1698175906
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1381
timestamp 1698175906
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1382
timestamp 1698175906
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1383
timestamp 1698175906
transform 1 0 67984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1384
timestamp 1698175906
transform 1 0 75824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1385
timestamp 1698175906
transform 1 0 83664 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1386
timestamp 1698175906
transform 1 0 91504 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1387
timestamp 1698175906
transform 1 0 99344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1388
timestamp 1698175906
transform 1 0 107184 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1389
timestamp 1698175906
transform 1 0 115024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1390
timestamp 1698175906
transform 1 0 122864 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1391
timestamp 1698175906
transform 1 0 130704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1392
timestamp 1698175906
transform 1 0 138544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1393
timestamp 1698175906
transform 1 0 146384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1394
timestamp 1698175906
transform 1 0 154224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1395
timestamp 1698175906
transform 1 0 162064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1396
timestamp 1698175906
transform 1 0 169904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1397
timestamp 1698175906
transform 1 0 177744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1398
timestamp 1698175906
transform 1 0 185584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1399
timestamp 1698175906
transform 1 0 193424 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1400
timestamp 1698175906
transform 1 0 201264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1401
timestamp 1698175906
transform 1 0 209104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1402
timestamp 1698175906
transform 1 0 216944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1403
timestamp 1698175906
transform 1 0 224784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1404
timestamp 1698175906
transform 1 0 232624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1405
timestamp 1698175906
transform 1 0 240464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1406
timestamp 1698175906
transform 1 0 248304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1407
timestamp 1698175906
transform 1 0 256144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1408
timestamp 1698175906
transform 1 0 263984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1409
timestamp 1698175906
transform 1 0 271824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1410
timestamp 1698175906
transform 1 0 279664 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1411
timestamp 1698175906
transform 1 0 287504 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1412
timestamp 1698175906
transform 1 0 295344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1413
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1414
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1415
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1416
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1417
timestamp 1698175906
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1418
timestamp 1698175906
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1419
timestamp 1698175906
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1420
timestamp 1698175906
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1421
timestamp 1698175906
transform 1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1422
timestamp 1698175906
transform 1 0 79744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1423
timestamp 1698175906
transform 1 0 87584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1424
timestamp 1698175906
transform 1 0 95424 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1425
timestamp 1698175906
transform 1 0 103264 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1426
timestamp 1698175906
transform 1 0 111104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1427
timestamp 1698175906
transform 1 0 118944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1428
timestamp 1698175906
transform 1 0 126784 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1429
timestamp 1698175906
transform 1 0 134624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1430
timestamp 1698175906
transform 1 0 142464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1431
timestamp 1698175906
transform 1 0 150304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1432
timestamp 1698175906
transform 1 0 158144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1433
timestamp 1698175906
transform 1 0 165984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1434
timestamp 1698175906
transform 1 0 173824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1435
timestamp 1698175906
transform 1 0 181664 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1436
timestamp 1698175906
transform 1 0 189504 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1437
timestamp 1698175906
transform 1 0 197344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1438
timestamp 1698175906
transform 1 0 205184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1439
timestamp 1698175906
transform 1 0 213024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1440
timestamp 1698175906
transform 1 0 220864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1441
timestamp 1698175906
transform 1 0 228704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1442
timestamp 1698175906
transform 1 0 236544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1443
timestamp 1698175906
transform 1 0 244384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1444
timestamp 1698175906
transform 1 0 252224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1445
timestamp 1698175906
transform 1 0 260064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1446
timestamp 1698175906
transform 1 0 267904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1447
timestamp 1698175906
transform 1 0 275744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1448
timestamp 1698175906
transform 1 0 283584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1449
timestamp 1698175906
transform 1 0 291424 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1450
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1451
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1452
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1453
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1454
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1455
timestamp 1698175906
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1456
timestamp 1698175906
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1457
timestamp 1698175906
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1458
timestamp 1698175906
transform 1 0 67984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1459
timestamp 1698175906
transform 1 0 75824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1460
timestamp 1698175906
transform 1 0 83664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1461
timestamp 1698175906
transform 1 0 91504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1462
timestamp 1698175906
transform 1 0 99344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1463
timestamp 1698175906
transform 1 0 107184 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1464
timestamp 1698175906
transform 1 0 115024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1465
timestamp 1698175906
transform 1 0 122864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1466
timestamp 1698175906
transform 1 0 130704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1467
timestamp 1698175906
transform 1 0 138544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1468
timestamp 1698175906
transform 1 0 146384 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1469
timestamp 1698175906
transform 1 0 154224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1470
timestamp 1698175906
transform 1 0 162064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1471
timestamp 1698175906
transform 1 0 169904 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1472
timestamp 1698175906
transform 1 0 177744 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1473
timestamp 1698175906
transform 1 0 185584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1474
timestamp 1698175906
transform 1 0 193424 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1475
timestamp 1698175906
transform 1 0 201264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1476
timestamp 1698175906
transform 1 0 209104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1477
timestamp 1698175906
transform 1 0 216944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1478
timestamp 1698175906
transform 1 0 224784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1479
timestamp 1698175906
transform 1 0 232624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1480
timestamp 1698175906
transform 1 0 240464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1481
timestamp 1698175906
transform 1 0 248304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1482
timestamp 1698175906
transform 1 0 256144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1483
timestamp 1698175906
transform 1 0 263984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1484
timestamp 1698175906
transform 1 0 271824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1485
timestamp 1698175906
transform 1 0 279664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1486
timestamp 1698175906
transform 1 0 287504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1487
timestamp 1698175906
transform 1 0 295344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1488
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1489
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1490
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1491
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1492
timestamp 1698175906
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1493
timestamp 1698175906
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1494
timestamp 1698175906
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1495
timestamp 1698175906
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1496
timestamp 1698175906
transform 1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1497
timestamp 1698175906
transform 1 0 79744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1498
timestamp 1698175906
transform 1 0 87584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1499
timestamp 1698175906
transform 1 0 95424 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1500
timestamp 1698175906
transform 1 0 103264 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1501
timestamp 1698175906
transform 1 0 111104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1502
timestamp 1698175906
transform 1 0 118944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1503
timestamp 1698175906
transform 1 0 126784 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1504
timestamp 1698175906
transform 1 0 134624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1505
timestamp 1698175906
transform 1 0 142464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1506
timestamp 1698175906
transform 1 0 150304 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1507
timestamp 1698175906
transform 1 0 158144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1508
timestamp 1698175906
transform 1 0 165984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1509
timestamp 1698175906
transform 1 0 173824 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1510
timestamp 1698175906
transform 1 0 181664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1511
timestamp 1698175906
transform 1 0 189504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1512
timestamp 1698175906
transform 1 0 197344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1513
timestamp 1698175906
transform 1 0 205184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1514
timestamp 1698175906
transform 1 0 213024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1515
timestamp 1698175906
transform 1 0 220864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1516
timestamp 1698175906
transform 1 0 228704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1517
timestamp 1698175906
transform 1 0 236544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1518
timestamp 1698175906
transform 1 0 244384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1519
timestamp 1698175906
transform 1 0 252224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1520
timestamp 1698175906
transform 1 0 260064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1521
timestamp 1698175906
transform 1 0 267904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1522
timestamp 1698175906
transform 1 0 275744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1523
timestamp 1698175906
transform 1 0 283584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1524
timestamp 1698175906
transform 1 0 291424 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1525
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1526
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1527
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1528
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1529
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1530
timestamp 1698175906
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1531
timestamp 1698175906
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1532
timestamp 1698175906
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1533
timestamp 1698175906
transform 1 0 67984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1534
timestamp 1698175906
transform 1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1535
timestamp 1698175906
transform 1 0 83664 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1536
timestamp 1698175906
transform 1 0 91504 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1537
timestamp 1698175906
transform 1 0 99344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1538
timestamp 1698175906
transform 1 0 107184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1539
timestamp 1698175906
transform 1 0 115024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1540
timestamp 1698175906
transform 1 0 122864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1541
timestamp 1698175906
transform 1 0 130704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1542
timestamp 1698175906
transform 1 0 138544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1543
timestamp 1698175906
transform 1 0 146384 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1544
timestamp 1698175906
transform 1 0 154224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1545
timestamp 1698175906
transform 1 0 162064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1546
timestamp 1698175906
transform 1 0 169904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1547
timestamp 1698175906
transform 1 0 177744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1548
timestamp 1698175906
transform 1 0 185584 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1549
timestamp 1698175906
transform 1 0 193424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1550
timestamp 1698175906
transform 1 0 201264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1551
timestamp 1698175906
transform 1 0 209104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1552
timestamp 1698175906
transform 1 0 216944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1553
timestamp 1698175906
transform 1 0 224784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1554
timestamp 1698175906
transform 1 0 232624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1555
timestamp 1698175906
transform 1 0 240464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1556
timestamp 1698175906
transform 1 0 248304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1557
timestamp 1698175906
transform 1 0 256144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1558
timestamp 1698175906
transform 1 0 263984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1559
timestamp 1698175906
transform 1 0 271824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1560
timestamp 1698175906
transform 1 0 279664 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1561
timestamp 1698175906
transform 1 0 287504 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1562
timestamp 1698175906
transform 1 0 295344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1563
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1564
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1565
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1566
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1567
timestamp 1698175906
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1568
timestamp 1698175906
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1569
timestamp 1698175906
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1570
timestamp 1698175906
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1571
timestamp 1698175906
transform 1 0 71904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1572
timestamp 1698175906
transform 1 0 79744 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1573
timestamp 1698175906
transform 1 0 87584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1574
timestamp 1698175906
transform 1 0 95424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1575
timestamp 1698175906
transform 1 0 103264 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1576
timestamp 1698175906
transform 1 0 111104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1577
timestamp 1698175906
transform 1 0 118944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1578
timestamp 1698175906
transform 1 0 126784 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1579
timestamp 1698175906
transform 1 0 134624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1580
timestamp 1698175906
transform 1 0 142464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1581
timestamp 1698175906
transform 1 0 150304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1582
timestamp 1698175906
transform 1 0 158144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1583
timestamp 1698175906
transform 1 0 165984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1584
timestamp 1698175906
transform 1 0 173824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1585
timestamp 1698175906
transform 1 0 181664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1586
timestamp 1698175906
transform 1 0 189504 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1587
timestamp 1698175906
transform 1 0 197344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1588
timestamp 1698175906
transform 1 0 205184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1589
timestamp 1698175906
transform 1 0 213024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1590
timestamp 1698175906
transform 1 0 220864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1591
timestamp 1698175906
transform 1 0 228704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1592
timestamp 1698175906
transform 1 0 236544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1593
timestamp 1698175906
transform 1 0 244384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1594
timestamp 1698175906
transform 1 0 252224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1595
timestamp 1698175906
transform 1 0 260064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1596
timestamp 1698175906
transform 1 0 267904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1597
timestamp 1698175906
transform 1 0 275744 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1598
timestamp 1698175906
transform 1 0 283584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1599
timestamp 1698175906
transform 1 0 291424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1600
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1601
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1602
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1603
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1604
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1605
timestamp 1698175906
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1606
timestamp 1698175906
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1607
timestamp 1698175906
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1608
timestamp 1698175906
transform 1 0 67984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1609
timestamp 1698175906
transform 1 0 75824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1610
timestamp 1698175906
transform 1 0 83664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1611
timestamp 1698175906
transform 1 0 91504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1612
timestamp 1698175906
transform 1 0 99344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1613
timestamp 1698175906
transform 1 0 107184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1614
timestamp 1698175906
transform 1 0 115024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1615
timestamp 1698175906
transform 1 0 122864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1616
timestamp 1698175906
transform 1 0 130704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1617
timestamp 1698175906
transform 1 0 138544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1618
timestamp 1698175906
transform 1 0 146384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1619
timestamp 1698175906
transform 1 0 154224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1620
timestamp 1698175906
transform 1 0 162064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1621
timestamp 1698175906
transform 1 0 169904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1622
timestamp 1698175906
transform 1 0 177744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1623
timestamp 1698175906
transform 1 0 185584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1624
timestamp 1698175906
transform 1 0 193424 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1625
timestamp 1698175906
transform 1 0 201264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1626
timestamp 1698175906
transform 1 0 209104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1627
timestamp 1698175906
transform 1 0 216944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1628
timestamp 1698175906
transform 1 0 224784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1629
timestamp 1698175906
transform 1 0 232624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1630
timestamp 1698175906
transform 1 0 240464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1631
timestamp 1698175906
transform 1 0 248304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1632
timestamp 1698175906
transform 1 0 256144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1633
timestamp 1698175906
transform 1 0 263984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1634
timestamp 1698175906
transform 1 0 271824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1635
timestamp 1698175906
transform 1 0 279664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1636
timestamp 1698175906
transform 1 0 287504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1637
timestamp 1698175906
transform 1 0 295344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1638
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1639
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1640
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1641
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1642
timestamp 1698175906
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1643
timestamp 1698175906
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1644
timestamp 1698175906
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1645
timestamp 1698175906
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1646
timestamp 1698175906
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1647
timestamp 1698175906
transform 1 0 79744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1648
timestamp 1698175906
transform 1 0 87584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1649
timestamp 1698175906
transform 1 0 95424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1650
timestamp 1698175906
transform 1 0 103264 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1651
timestamp 1698175906
transform 1 0 111104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1652
timestamp 1698175906
transform 1 0 118944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1653
timestamp 1698175906
transform 1 0 126784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1654
timestamp 1698175906
transform 1 0 134624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1655
timestamp 1698175906
transform 1 0 142464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1656
timestamp 1698175906
transform 1 0 150304 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1657
timestamp 1698175906
transform 1 0 158144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1658
timestamp 1698175906
transform 1 0 165984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1659
timestamp 1698175906
transform 1 0 173824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1660
timestamp 1698175906
transform 1 0 181664 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1661
timestamp 1698175906
transform 1 0 189504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1662
timestamp 1698175906
transform 1 0 197344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1663
timestamp 1698175906
transform 1 0 205184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1664
timestamp 1698175906
transform 1 0 213024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1665
timestamp 1698175906
transform 1 0 220864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1666
timestamp 1698175906
transform 1 0 228704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1667
timestamp 1698175906
transform 1 0 236544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1668
timestamp 1698175906
transform 1 0 244384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1669
timestamp 1698175906
transform 1 0 252224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1670
timestamp 1698175906
transform 1 0 260064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1671
timestamp 1698175906
transform 1 0 267904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1672
timestamp 1698175906
transform 1 0 275744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1673
timestamp 1698175906
transform 1 0 283584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1674
timestamp 1698175906
transform 1 0 291424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1675
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1676
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1677
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1678
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1679
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1680
timestamp 1698175906
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1681
timestamp 1698175906
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1682
timestamp 1698175906
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1683
timestamp 1698175906
transform 1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1684
timestamp 1698175906
transform 1 0 75824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1685
timestamp 1698175906
transform 1 0 83664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1686
timestamp 1698175906
transform 1 0 91504 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1687
timestamp 1698175906
transform 1 0 99344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1688
timestamp 1698175906
transform 1 0 107184 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1689
timestamp 1698175906
transform 1 0 115024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1690
timestamp 1698175906
transform 1 0 122864 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1691
timestamp 1698175906
transform 1 0 130704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1692
timestamp 1698175906
transform 1 0 138544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1693
timestamp 1698175906
transform 1 0 146384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1694
timestamp 1698175906
transform 1 0 154224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1695
timestamp 1698175906
transform 1 0 162064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1696
timestamp 1698175906
transform 1 0 169904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1697
timestamp 1698175906
transform 1 0 177744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1698
timestamp 1698175906
transform 1 0 185584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1699
timestamp 1698175906
transform 1 0 193424 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1700
timestamp 1698175906
transform 1 0 201264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1701
timestamp 1698175906
transform 1 0 209104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1702
timestamp 1698175906
transform 1 0 216944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1703
timestamp 1698175906
transform 1 0 224784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1704
timestamp 1698175906
transform 1 0 232624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1705
timestamp 1698175906
transform 1 0 240464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1706
timestamp 1698175906
transform 1 0 248304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1707
timestamp 1698175906
transform 1 0 256144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1708
timestamp 1698175906
transform 1 0 263984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1709
timestamp 1698175906
transform 1 0 271824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1710
timestamp 1698175906
transform 1 0 279664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1711
timestamp 1698175906
transform 1 0 287504 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1712
timestamp 1698175906
transform 1 0 295344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1713
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1714
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1715
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1716
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1717
timestamp 1698175906
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1718
timestamp 1698175906
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1719
timestamp 1698175906
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1720
timestamp 1698175906
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1721
timestamp 1698175906
transform 1 0 71904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1722
timestamp 1698175906
transform 1 0 79744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1723
timestamp 1698175906
transform 1 0 87584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1724
timestamp 1698175906
transform 1 0 95424 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1725
timestamp 1698175906
transform 1 0 103264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1726
timestamp 1698175906
transform 1 0 111104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1727
timestamp 1698175906
transform 1 0 118944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1728
timestamp 1698175906
transform 1 0 126784 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1729
timestamp 1698175906
transform 1 0 134624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1730
timestamp 1698175906
transform 1 0 142464 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1731
timestamp 1698175906
transform 1 0 150304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1732
timestamp 1698175906
transform 1 0 158144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1733
timestamp 1698175906
transform 1 0 165984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1734
timestamp 1698175906
transform 1 0 173824 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1735
timestamp 1698175906
transform 1 0 181664 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1736
timestamp 1698175906
transform 1 0 189504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1737
timestamp 1698175906
transform 1 0 197344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1738
timestamp 1698175906
transform 1 0 205184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1739
timestamp 1698175906
transform 1 0 213024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1740
timestamp 1698175906
transform 1 0 220864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1741
timestamp 1698175906
transform 1 0 228704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1742
timestamp 1698175906
transform 1 0 236544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1743
timestamp 1698175906
transform 1 0 244384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1744
timestamp 1698175906
transform 1 0 252224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1745
timestamp 1698175906
transform 1 0 260064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1746
timestamp 1698175906
transform 1 0 267904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1747
timestamp 1698175906
transform 1 0 275744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1748
timestamp 1698175906
transform 1 0 283584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1749
timestamp 1698175906
transform 1 0 291424 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1750
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1751
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1752
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1753
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1754
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1755
timestamp 1698175906
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1756
timestamp 1698175906
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1757
timestamp 1698175906
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1758
timestamp 1698175906
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1759
timestamp 1698175906
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1760
timestamp 1698175906
transform 1 0 83664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1761
timestamp 1698175906
transform 1 0 91504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1762
timestamp 1698175906
transform 1 0 99344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1763
timestamp 1698175906
transform 1 0 107184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1764
timestamp 1698175906
transform 1 0 115024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1765
timestamp 1698175906
transform 1 0 122864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1766
timestamp 1698175906
transform 1 0 130704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1767
timestamp 1698175906
transform 1 0 138544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1768
timestamp 1698175906
transform 1 0 146384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1769
timestamp 1698175906
transform 1 0 154224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1770
timestamp 1698175906
transform 1 0 162064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1771
timestamp 1698175906
transform 1 0 169904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1772
timestamp 1698175906
transform 1 0 177744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1773
timestamp 1698175906
transform 1 0 185584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1774
timestamp 1698175906
transform 1 0 193424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1775
timestamp 1698175906
transform 1 0 201264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1776
timestamp 1698175906
transform 1 0 209104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1777
timestamp 1698175906
transform 1 0 216944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1778
timestamp 1698175906
transform 1 0 224784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1779
timestamp 1698175906
transform 1 0 232624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1780
timestamp 1698175906
transform 1 0 240464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1781
timestamp 1698175906
transform 1 0 248304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1782
timestamp 1698175906
transform 1 0 256144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1783
timestamp 1698175906
transform 1 0 263984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1784
timestamp 1698175906
transform 1 0 271824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1785
timestamp 1698175906
transform 1 0 279664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1786
timestamp 1698175906
transform 1 0 287504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1787
timestamp 1698175906
transform 1 0 295344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1788
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1789
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1790
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1791
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1792
timestamp 1698175906
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1793
timestamp 1698175906
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1794
timestamp 1698175906
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1795
timestamp 1698175906
transform 1 0 64064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1796
timestamp 1698175906
transform 1 0 71904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1797
timestamp 1698175906
transform 1 0 79744 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1798
timestamp 1698175906
transform 1 0 87584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1799
timestamp 1698175906
transform 1 0 95424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1800
timestamp 1698175906
transform 1 0 103264 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1801
timestamp 1698175906
transform 1 0 111104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1802
timestamp 1698175906
transform 1 0 118944 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1803
timestamp 1698175906
transform 1 0 126784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1804
timestamp 1698175906
transform 1 0 134624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1805
timestamp 1698175906
transform 1 0 142464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1806
timestamp 1698175906
transform 1 0 150304 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1807
timestamp 1698175906
transform 1 0 158144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1808
timestamp 1698175906
transform 1 0 165984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1809
timestamp 1698175906
transform 1 0 173824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1810
timestamp 1698175906
transform 1 0 181664 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1811
timestamp 1698175906
transform 1 0 189504 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1812
timestamp 1698175906
transform 1 0 197344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1813
timestamp 1698175906
transform 1 0 205184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1814
timestamp 1698175906
transform 1 0 213024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1815
timestamp 1698175906
transform 1 0 220864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1816
timestamp 1698175906
transform 1 0 228704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1817
timestamp 1698175906
transform 1 0 236544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1818
timestamp 1698175906
transform 1 0 244384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1819
timestamp 1698175906
transform 1 0 252224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1820
timestamp 1698175906
transform 1 0 260064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1821
timestamp 1698175906
transform 1 0 267904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1822
timestamp 1698175906
transform 1 0 275744 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1823
timestamp 1698175906
transform 1 0 283584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1824
timestamp 1698175906
transform 1 0 291424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1825
timestamp 1698175906
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1826
timestamp 1698175906
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1827
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1828
timestamp 1698175906
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1829
timestamp 1698175906
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1830
timestamp 1698175906
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1831
timestamp 1698175906
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1832
timestamp 1698175906
transform 1 0 60144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1833
timestamp 1698175906
transform 1 0 67984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1834
timestamp 1698175906
transform 1 0 75824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1835
timestamp 1698175906
transform 1 0 83664 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1836
timestamp 1698175906
transform 1 0 91504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1837
timestamp 1698175906
transform 1 0 99344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1838
timestamp 1698175906
transform 1 0 107184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1839
timestamp 1698175906
transform 1 0 115024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1840
timestamp 1698175906
transform 1 0 122864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1841
timestamp 1698175906
transform 1 0 130704 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1842
timestamp 1698175906
transform 1 0 138544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1843
timestamp 1698175906
transform 1 0 146384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1844
timestamp 1698175906
transform 1 0 154224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1845
timestamp 1698175906
transform 1 0 162064 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1846
timestamp 1698175906
transform 1 0 169904 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1847
timestamp 1698175906
transform 1 0 177744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1848
timestamp 1698175906
transform 1 0 185584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1849
timestamp 1698175906
transform 1 0 193424 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1850
timestamp 1698175906
transform 1 0 201264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1851
timestamp 1698175906
transform 1 0 209104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1852
timestamp 1698175906
transform 1 0 216944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1853
timestamp 1698175906
transform 1 0 224784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1854
timestamp 1698175906
transform 1 0 232624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1855
timestamp 1698175906
transform 1 0 240464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1856
timestamp 1698175906
transform 1 0 248304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1857
timestamp 1698175906
transform 1 0 256144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1858
timestamp 1698175906
transform 1 0 263984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1859
timestamp 1698175906
transform 1 0 271824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1860
timestamp 1698175906
transform 1 0 279664 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1861
timestamp 1698175906
transform 1 0 287504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1862
timestamp 1698175906
transform 1 0 295344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1863
timestamp 1698175906
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1864
timestamp 1698175906
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1865
timestamp 1698175906
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1866
timestamp 1698175906
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1867
timestamp 1698175906
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1868
timestamp 1698175906
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1869
timestamp 1698175906
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1870
timestamp 1698175906
transform 1 0 64064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1871
timestamp 1698175906
transform 1 0 71904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1872
timestamp 1698175906
transform 1 0 79744 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1873
timestamp 1698175906
transform 1 0 87584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1874
timestamp 1698175906
transform 1 0 95424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1875
timestamp 1698175906
transform 1 0 103264 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1876
timestamp 1698175906
transform 1 0 111104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1877
timestamp 1698175906
transform 1 0 118944 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1878
timestamp 1698175906
transform 1 0 126784 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1879
timestamp 1698175906
transform 1 0 134624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1880
timestamp 1698175906
transform 1 0 142464 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1881
timestamp 1698175906
transform 1 0 150304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1882
timestamp 1698175906
transform 1 0 158144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1883
timestamp 1698175906
transform 1 0 165984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1884
timestamp 1698175906
transform 1 0 173824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1885
timestamp 1698175906
transform 1 0 181664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1886
timestamp 1698175906
transform 1 0 189504 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1887
timestamp 1698175906
transform 1 0 197344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1888
timestamp 1698175906
transform 1 0 205184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1889
timestamp 1698175906
transform 1 0 213024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1890
timestamp 1698175906
transform 1 0 220864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1891
timestamp 1698175906
transform 1 0 228704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1892
timestamp 1698175906
transform 1 0 236544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1893
timestamp 1698175906
transform 1 0 244384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1894
timestamp 1698175906
transform 1 0 252224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1895
timestamp 1698175906
transform 1 0 260064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1896
timestamp 1698175906
transform 1 0 267904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1897
timestamp 1698175906
transform 1 0 275744 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1898
timestamp 1698175906
transform 1 0 283584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1899
timestamp 1698175906
transform 1 0 291424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1900
timestamp 1698175906
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1901
timestamp 1698175906
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1902
timestamp 1698175906
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1903
timestamp 1698175906
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1904
timestamp 1698175906
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1905
timestamp 1698175906
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1906
timestamp 1698175906
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1907
timestamp 1698175906
transform 1 0 60144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1908
timestamp 1698175906
transform 1 0 67984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1909
timestamp 1698175906
transform 1 0 75824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1910
timestamp 1698175906
transform 1 0 83664 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1911
timestamp 1698175906
transform 1 0 91504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1912
timestamp 1698175906
transform 1 0 99344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1913
timestamp 1698175906
transform 1 0 107184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1914
timestamp 1698175906
transform 1 0 115024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1915
timestamp 1698175906
transform 1 0 122864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1916
timestamp 1698175906
transform 1 0 130704 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1917
timestamp 1698175906
transform 1 0 138544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1918
timestamp 1698175906
transform 1 0 146384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1919
timestamp 1698175906
transform 1 0 154224 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1920
timestamp 1698175906
transform 1 0 162064 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1921
timestamp 1698175906
transform 1 0 169904 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1922
timestamp 1698175906
transform 1 0 177744 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1923
timestamp 1698175906
transform 1 0 185584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1924
timestamp 1698175906
transform 1 0 193424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1925
timestamp 1698175906
transform 1 0 201264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1926
timestamp 1698175906
transform 1 0 209104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1927
timestamp 1698175906
transform 1 0 216944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1928
timestamp 1698175906
transform 1 0 224784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1929
timestamp 1698175906
transform 1 0 232624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1930
timestamp 1698175906
transform 1 0 240464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1931
timestamp 1698175906
transform 1 0 248304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1932
timestamp 1698175906
transform 1 0 256144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1933
timestamp 1698175906
transform 1 0 263984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1934
timestamp 1698175906
transform 1 0 271824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1935
timestamp 1698175906
transform 1 0 279664 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1936
timestamp 1698175906
transform 1 0 287504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1937
timestamp 1698175906
transform 1 0 295344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1938
timestamp 1698175906
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1939
timestamp 1698175906
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1940
timestamp 1698175906
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1941
timestamp 1698175906
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1942
timestamp 1698175906
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1943
timestamp 1698175906
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1944
timestamp 1698175906
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1945
timestamp 1698175906
transform 1 0 64064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1946
timestamp 1698175906
transform 1 0 71904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1947
timestamp 1698175906
transform 1 0 79744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1948
timestamp 1698175906
transform 1 0 87584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1949
timestamp 1698175906
transform 1 0 95424 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1950
timestamp 1698175906
transform 1 0 103264 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1951
timestamp 1698175906
transform 1 0 111104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1952
timestamp 1698175906
transform 1 0 118944 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1953
timestamp 1698175906
transform 1 0 126784 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1954
timestamp 1698175906
transform 1 0 134624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1955
timestamp 1698175906
transform 1 0 142464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1956
timestamp 1698175906
transform 1 0 150304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1957
timestamp 1698175906
transform 1 0 158144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1958
timestamp 1698175906
transform 1 0 165984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1959
timestamp 1698175906
transform 1 0 173824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1960
timestamp 1698175906
transform 1 0 181664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1961
timestamp 1698175906
transform 1 0 189504 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1962
timestamp 1698175906
transform 1 0 197344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1963
timestamp 1698175906
transform 1 0 205184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1964
timestamp 1698175906
transform 1 0 213024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1965
timestamp 1698175906
transform 1 0 220864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1966
timestamp 1698175906
transform 1 0 228704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1967
timestamp 1698175906
transform 1 0 236544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1968
timestamp 1698175906
transform 1 0 244384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1969
timestamp 1698175906
transform 1 0 252224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1970
timestamp 1698175906
transform 1 0 260064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1971
timestamp 1698175906
transform 1 0 267904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1972
timestamp 1698175906
transform 1 0 275744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1973
timestamp 1698175906
transform 1 0 283584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1974
timestamp 1698175906
transform 1 0 291424 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1975
timestamp 1698175906
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1976
timestamp 1698175906
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1977
timestamp 1698175906
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1978
timestamp 1698175906
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1979
timestamp 1698175906
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1980
timestamp 1698175906
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1981
timestamp 1698175906
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1982
timestamp 1698175906
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1983
timestamp 1698175906
transform 1 0 67984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1984
timestamp 1698175906
transform 1 0 75824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1985
timestamp 1698175906
transform 1 0 83664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1986
timestamp 1698175906
transform 1 0 91504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1987
timestamp 1698175906
transform 1 0 99344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1988
timestamp 1698175906
transform 1 0 107184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1989
timestamp 1698175906
transform 1 0 115024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1990
timestamp 1698175906
transform 1 0 122864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1991
timestamp 1698175906
transform 1 0 130704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1992
timestamp 1698175906
transform 1 0 138544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1993
timestamp 1698175906
transform 1 0 146384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1994
timestamp 1698175906
transform 1 0 154224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1995
timestamp 1698175906
transform 1 0 162064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1996
timestamp 1698175906
transform 1 0 169904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1997
timestamp 1698175906
transform 1 0 177744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1998
timestamp 1698175906
transform 1 0 185584 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1999
timestamp 1698175906
transform 1 0 193424 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2000
timestamp 1698175906
transform 1 0 201264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2001
timestamp 1698175906
transform 1 0 209104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2002
timestamp 1698175906
transform 1 0 216944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2003
timestamp 1698175906
transform 1 0 224784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2004
timestamp 1698175906
transform 1 0 232624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2005
timestamp 1698175906
transform 1 0 240464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2006
timestamp 1698175906
transform 1 0 248304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2007
timestamp 1698175906
transform 1 0 256144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2008
timestamp 1698175906
transform 1 0 263984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2009
timestamp 1698175906
transform 1 0 271824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2010
timestamp 1698175906
transform 1 0 279664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2011
timestamp 1698175906
transform 1 0 287504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2012
timestamp 1698175906
transform 1 0 295344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2013
timestamp 1698175906
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2014
timestamp 1698175906
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2015
timestamp 1698175906
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2016
timestamp 1698175906
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2017
timestamp 1698175906
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2018
timestamp 1698175906
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2019
timestamp 1698175906
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2020
timestamp 1698175906
transform 1 0 64064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2021
timestamp 1698175906
transform 1 0 71904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2022
timestamp 1698175906
transform 1 0 79744 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2023
timestamp 1698175906
transform 1 0 87584 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2024
timestamp 1698175906
transform 1 0 95424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2025
timestamp 1698175906
transform 1 0 103264 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2026
timestamp 1698175906
transform 1 0 111104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2027
timestamp 1698175906
transform 1 0 118944 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2028
timestamp 1698175906
transform 1 0 126784 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2029
timestamp 1698175906
transform 1 0 134624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2030
timestamp 1698175906
transform 1 0 142464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2031
timestamp 1698175906
transform 1 0 150304 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2032
timestamp 1698175906
transform 1 0 158144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2033
timestamp 1698175906
transform 1 0 165984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2034
timestamp 1698175906
transform 1 0 173824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2035
timestamp 1698175906
transform 1 0 181664 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2036
timestamp 1698175906
transform 1 0 189504 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2037
timestamp 1698175906
transform 1 0 197344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2038
timestamp 1698175906
transform 1 0 205184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2039
timestamp 1698175906
transform 1 0 213024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2040
timestamp 1698175906
transform 1 0 220864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2041
timestamp 1698175906
transform 1 0 228704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2042
timestamp 1698175906
transform 1 0 236544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2043
timestamp 1698175906
transform 1 0 244384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2044
timestamp 1698175906
transform 1 0 252224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2045
timestamp 1698175906
transform 1 0 260064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2046
timestamp 1698175906
transform 1 0 267904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2047
timestamp 1698175906
transform 1 0 275744 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2048
timestamp 1698175906
transform 1 0 283584 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2049
timestamp 1698175906
transform 1 0 291424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2050
timestamp 1698175906
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2051
timestamp 1698175906
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2052
timestamp 1698175906
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2053
timestamp 1698175906
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2054
timestamp 1698175906
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2055
timestamp 1698175906
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2056
timestamp 1698175906
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2057
timestamp 1698175906
transform 1 0 60144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2058
timestamp 1698175906
transform 1 0 67984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2059
timestamp 1698175906
transform 1 0 75824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2060
timestamp 1698175906
transform 1 0 83664 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2061
timestamp 1698175906
transform 1 0 91504 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2062
timestamp 1698175906
transform 1 0 99344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2063
timestamp 1698175906
transform 1 0 107184 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2064
timestamp 1698175906
transform 1 0 115024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2065
timestamp 1698175906
transform 1 0 122864 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2066
timestamp 1698175906
transform 1 0 130704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2067
timestamp 1698175906
transform 1 0 138544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2068
timestamp 1698175906
transform 1 0 146384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2069
timestamp 1698175906
transform 1 0 154224 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2070
timestamp 1698175906
transform 1 0 162064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2071
timestamp 1698175906
transform 1 0 169904 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2072
timestamp 1698175906
transform 1 0 177744 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2073
timestamp 1698175906
transform 1 0 185584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2074
timestamp 1698175906
transform 1 0 193424 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2075
timestamp 1698175906
transform 1 0 201264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2076
timestamp 1698175906
transform 1 0 209104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2077
timestamp 1698175906
transform 1 0 216944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2078
timestamp 1698175906
transform 1 0 224784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2079
timestamp 1698175906
transform 1 0 232624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2080
timestamp 1698175906
transform 1 0 240464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2081
timestamp 1698175906
transform 1 0 248304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2082
timestamp 1698175906
transform 1 0 256144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2083
timestamp 1698175906
transform 1 0 263984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2084
timestamp 1698175906
transform 1 0 271824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2085
timestamp 1698175906
transform 1 0 279664 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2086
timestamp 1698175906
transform 1 0 287504 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2087
timestamp 1698175906
transform 1 0 295344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2088
timestamp 1698175906
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2089
timestamp 1698175906
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2090
timestamp 1698175906
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2091
timestamp 1698175906
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2092
timestamp 1698175906
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2093
timestamp 1698175906
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2094
timestamp 1698175906
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2095
timestamp 1698175906
transform 1 0 64064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2096
timestamp 1698175906
transform 1 0 71904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2097
timestamp 1698175906
transform 1 0 79744 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2098
timestamp 1698175906
transform 1 0 87584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2099
timestamp 1698175906
transform 1 0 95424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2100
timestamp 1698175906
transform 1 0 103264 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2101
timestamp 1698175906
transform 1 0 111104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2102
timestamp 1698175906
transform 1 0 118944 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2103
timestamp 1698175906
transform 1 0 126784 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2104
timestamp 1698175906
transform 1 0 134624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2105
timestamp 1698175906
transform 1 0 142464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2106
timestamp 1698175906
transform 1 0 150304 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2107
timestamp 1698175906
transform 1 0 158144 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2108
timestamp 1698175906
transform 1 0 165984 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2109
timestamp 1698175906
transform 1 0 173824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2110
timestamp 1698175906
transform 1 0 181664 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2111
timestamp 1698175906
transform 1 0 189504 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2112
timestamp 1698175906
transform 1 0 197344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2113
timestamp 1698175906
transform 1 0 205184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2114
timestamp 1698175906
transform 1 0 213024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2115
timestamp 1698175906
transform 1 0 220864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2116
timestamp 1698175906
transform 1 0 228704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2117
timestamp 1698175906
transform 1 0 236544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2118
timestamp 1698175906
transform 1 0 244384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2119
timestamp 1698175906
transform 1 0 252224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2120
timestamp 1698175906
transform 1 0 260064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2121
timestamp 1698175906
transform 1 0 267904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2122
timestamp 1698175906
transform 1 0 275744 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2123
timestamp 1698175906
transform 1 0 283584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2124
timestamp 1698175906
transform 1 0 291424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2125
timestamp 1698175906
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2126
timestamp 1698175906
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2127
timestamp 1698175906
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2128
timestamp 1698175906
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2129
timestamp 1698175906
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2130
timestamp 1698175906
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2131
timestamp 1698175906
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2132
timestamp 1698175906
transform 1 0 60144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2133
timestamp 1698175906
transform 1 0 67984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2134
timestamp 1698175906
transform 1 0 75824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2135
timestamp 1698175906
transform 1 0 83664 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2136
timestamp 1698175906
transform 1 0 91504 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2137
timestamp 1698175906
transform 1 0 99344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2138
timestamp 1698175906
transform 1 0 107184 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2139
timestamp 1698175906
transform 1 0 115024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2140
timestamp 1698175906
transform 1 0 122864 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2141
timestamp 1698175906
transform 1 0 130704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2142
timestamp 1698175906
transform 1 0 138544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2143
timestamp 1698175906
transform 1 0 146384 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2144
timestamp 1698175906
transform 1 0 154224 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2145
timestamp 1698175906
transform 1 0 162064 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2146
timestamp 1698175906
transform 1 0 169904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2147
timestamp 1698175906
transform 1 0 177744 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2148
timestamp 1698175906
transform 1 0 185584 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2149
timestamp 1698175906
transform 1 0 193424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2150
timestamp 1698175906
transform 1 0 201264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2151
timestamp 1698175906
transform 1 0 209104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2152
timestamp 1698175906
transform 1 0 216944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2153
timestamp 1698175906
transform 1 0 224784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2154
timestamp 1698175906
transform 1 0 232624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2155
timestamp 1698175906
transform 1 0 240464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2156
timestamp 1698175906
transform 1 0 248304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2157
timestamp 1698175906
transform 1 0 256144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2158
timestamp 1698175906
transform 1 0 263984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2159
timestamp 1698175906
transform 1 0 271824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2160
timestamp 1698175906
transform 1 0 279664 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2161
timestamp 1698175906
transform 1 0 287504 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2162
timestamp 1698175906
transform 1 0 295344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2163
timestamp 1698175906
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2164
timestamp 1698175906
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2165
timestamp 1698175906
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2166
timestamp 1698175906
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2167
timestamp 1698175906
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2168
timestamp 1698175906
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2169
timestamp 1698175906
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2170
timestamp 1698175906
transform 1 0 64064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2171
timestamp 1698175906
transform 1 0 71904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2172
timestamp 1698175906
transform 1 0 79744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2173
timestamp 1698175906
transform 1 0 87584 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2174
timestamp 1698175906
transform 1 0 95424 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2175
timestamp 1698175906
transform 1 0 103264 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2176
timestamp 1698175906
transform 1 0 111104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2177
timestamp 1698175906
transform 1 0 118944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2178
timestamp 1698175906
transform 1 0 126784 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2179
timestamp 1698175906
transform 1 0 134624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2180
timestamp 1698175906
transform 1 0 142464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2181
timestamp 1698175906
transform 1 0 150304 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2182
timestamp 1698175906
transform 1 0 158144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2183
timestamp 1698175906
transform 1 0 165984 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2184
timestamp 1698175906
transform 1 0 173824 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2185
timestamp 1698175906
transform 1 0 181664 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2186
timestamp 1698175906
transform 1 0 189504 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2187
timestamp 1698175906
transform 1 0 197344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2188
timestamp 1698175906
transform 1 0 205184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2189
timestamp 1698175906
transform 1 0 213024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2190
timestamp 1698175906
transform 1 0 220864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2191
timestamp 1698175906
transform 1 0 228704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2192
timestamp 1698175906
transform 1 0 236544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2193
timestamp 1698175906
transform 1 0 244384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2194
timestamp 1698175906
transform 1 0 252224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2195
timestamp 1698175906
transform 1 0 260064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2196
timestamp 1698175906
transform 1 0 267904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2197
timestamp 1698175906
transform 1 0 275744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2198
timestamp 1698175906
transform 1 0 283584 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2199
timestamp 1698175906
transform 1 0 291424 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2200
timestamp 1698175906
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2201
timestamp 1698175906
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2202
timestamp 1698175906
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2203
timestamp 1698175906
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2204
timestamp 1698175906
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2205
timestamp 1698175906
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2206
timestamp 1698175906
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2207
timestamp 1698175906
transform 1 0 60144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2208
timestamp 1698175906
transform 1 0 67984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2209
timestamp 1698175906
transform 1 0 75824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2210
timestamp 1698175906
transform 1 0 83664 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2211
timestamp 1698175906
transform 1 0 91504 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2212
timestamp 1698175906
transform 1 0 99344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2213
timestamp 1698175906
transform 1 0 107184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2214
timestamp 1698175906
transform 1 0 115024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2215
timestamp 1698175906
transform 1 0 122864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2216
timestamp 1698175906
transform 1 0 130704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2217
timestamp 1698175906
transform 1 0 138544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2218
timestamp 1698175906
transform 1 0 146384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2219
timestamp 1698175906
transform 1 0 154224 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2220
timestamp 1698175906
transform 1 0 162064 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2221
timestamp 1698175906
transform 1 0 169904 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2222
timestamp 1698175906
transform 1 0 177744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2223
timestamp 1698175906
transform 1 0 185584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2224
timestamp 1698175906
transform 1 0 193424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2225
timestamp 1698175906
transform 1 0 201264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2226
timestamp 1698175906
transform 1 0 209104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2227
timestamp 1698175906
transform 1 0 216944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2228
timestamp 1698175906
transform 1 0 224784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2229
timestamp 1698175906
transform 1 0 232624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2230
timestamp 1698175906
transform 1 0 240464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2231
timestamp 1698175906
transform 1 0 248304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2232
timestamp 1698175906
transform 1 0 256144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2233
timestamp 1698175906
transform 1 0 263984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2234
timestamp 1698175906
transform 1 0 271824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2235
timestamp 1698175906
transform 1 0 279664 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2236
timestamp 1698175906
transform 1 0 287504 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2237
timestamp 1698175906
transform 1 0 295344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2238
timestamp 1698175906
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2239
timestamp 1698175906
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2240
timestamp 1698175906
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2241
timestamp 1698175906
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2242
timestamp 1698175906
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2243
timestamp 1698175906
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2244
timestamp 1698175906
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2245
timestamp 1698175906
transform 1 0 64064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2246
timestamp 1698175906
transform 1 0 71904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2247
timestamp 1698175906
transform 1 0 79744 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2248
timestamp 1698175906
transform 1 0 87584 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2249
timestamp 1698175906
transform 1 0 95424 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2250
timestamp 1698175906
transform 1 0 103264 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2251
timestamp 1698175906
transform 1 0 111104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2252
timestamp 1698175906
transform 1 0 118944 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2253
timestamp 1698175906
transform 1 0 126784 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2254
timestamp 1698175906
transform 1 0 134624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2255
timestamp 1698175906
transform 1 0 142464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2256
timestamp 1698175906
transform 1 0 150304 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2257
timestamp 1698175906
transform 1 0 158144 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2258
timestamp 1698175906
transform 1 0 165984 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2259
timestamp 1698175906
transform 1 0 173824 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2260
timestamp 1698175906
transform 1 0 181664 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2261
timestamp 1698175906
transform 1 0 189504 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2262
timestamp 1698175906
transform 1 0 197344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2263
timestamp 1698175906
transform 1 0 205184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2264
timestamp 1698175906
transform 1 0 213024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2265
timestamp 1698175906
transform 1 0 220864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2266
timestamp 1698175906
transform 1 0 228704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2267
timestamp 1698175906
transform 1 0 236544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2268
timestamp 1698175906
transform 1 0 244384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2269
timestamp 1698175906
transform 1 0 252224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2270
timestamp 1698175906
transform 1 0 260064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2271
timestamp 1698175906
transform 1 0 267904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2272
timestamp 1698175906
transform 1 0 275744 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2273
timestamp 1698175906
transform 1 0 283584 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2274
timestamp 1698175906
transform 1 0 291424 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2275
timestamp 1698175906
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2276
timestamp 1698175906
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2277
timestamp 1698175906
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2278
timestamp 1698175906
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2279
timestamp 1698175906
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2280
timestamp 1698175906
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2281
timestamp 1698175906
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2282
timestamp 1698175906
transform 1 0 60144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2283
timestamp 1698175906
transform 1 0 67984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2284
timestamp 1698175906
transform 1 0 75824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2285
timestamp 1698175906
transform 1 0 83664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2286
timestamp 1698175906
transform 1 0 91504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2287
timestamp 1698175906
transform 1 0 99344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2288
timestamp 1698175906
transform 1 0 107184 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2289
timestamp 1698175906
transform 1 0 115024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2290
timestamp 1698175906
transform 1 0 122864 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2291
timestamp 1698175906
transform 1 0 130704 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2292
timestamp 1698175906
transform 1 0 138544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2293
timestamp 1698175906
transform 1 0 146384 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2294
timestamp 1698175906
transform 1 0 154224 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2295
timestamp 1698175906
transform 1 0 162064 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2296
timestamp 1698175906
transform 1 0 169904 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2297
timestamp 1698175906
transform 1 0 177744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2298
timestamp 1698175906
transform 1 0 185584 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2299
timestamp 1698175906
transform 1 0 193424 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2300
timestamp 1698175906
transform 1 0 201264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2301
timestamp 1698175906
transform 1 0 209104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2302
timestamp 1698175906
transform 1 0 216944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2303
timestamp 1698175906
transform 1 0 224784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2304
timestamp 1698175906
transform 1 0 232624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2305
timestamp 1698175906
transform 1 0 240464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2306
timestamp 1698175906
transform 1 0 248304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2307
timestamp 1698175906
transform 1 0 256144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2308
timestamp 1698175906
transform 1 0 263984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2309
timestamp 1698175906
transform 1 0 271824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2310
timestamp 1698175906
transform 1 0 279664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2311
timestamp 1698175906
transform 1 0 287504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2312
timestamp 1698175906
transform 1 0 295344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2313
timestamp 1698175906
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2314
timestamp 1698175906
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2315
timestamp 1698175906
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2316
timestamp 1698175906
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2317
timestamp 1698175906
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2318
timestamp 1698175906
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2319
timestamp 1698175906
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2320
timestamp 1698175906
transform 1 0 64064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2321
timestamp 1698175906
transform 1 0 71904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2322
timestamp 1698175906
transform 1 0 79744 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2323
timestamp 1698175906
transform 1 0 87584 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2324
timestamp 1698175906
transform 1 0 95424 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2325
timestamp 1698175906
transform 1 0 103264 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2326
timestamp 1698175906
transform 1 0 111104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2327
timestamp 1698175906
transform 1 0 118944 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2328
timestamp 1698175906
transform 1 0 126784 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2329
timestamp 1698175906
transform 1 0 134624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2330
timestamp 1698175906
transform 1 0 142464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2331
timestamp 1698175906
transform 1 0 150304 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2332
timestamp 1698175906
transform 1 0 158144 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2333
timestamp 1698175906
transform 1 0 165984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2334
timestamp 1698175906
transform 1 0 173824 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2335
timestamp 1698175906
transform 1 0 181664 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2336
timestamp 1698175906
transform 1 0 189504 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2337
timestamp 1698175906
transform 1 0 197344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2338
timestamp 1698175906
transform 1 0 205184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2339
timestamp 1698175906
transform 1 0 213024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2340
timestamp 1698175906
transform 1 0 220864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2341
timestamp 1698175906
transform 1 0 228704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2342
timestamp 1698175906
transform 1 0 236544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2343
timestamp 1698175906
transform 1 0 244384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2344
timestamp 1698175906
transform 1 0 252224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2345
timestamp 1698175906
transform 1 0 260064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2346
timestamp 1698175906
transform 1 0 267904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2347
timestamp 1698175906
transform 1 0 275744 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2348
timestamp 1698175906
transform 1 0 283584 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2349
timestamp 1698175906
transform 1 0 291424 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2350
timestamp 1698175906
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2351
timestamp 1698175906
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2352
timestamp 1698175906
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2353
timestamp 1698175906
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2354
timestamp 1698175906
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2355
timestamp 1698175906
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2356
timestamp 1698175906
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2357
timestamp 1698175906
transform 1 0 60144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2358
timestamp 1698175906
transform 1 0 67984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2359
timestamp 1698175906
transform 1 0 75824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2360
timestamp 1698175906
transform 1 0 83664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2361
timestamp 1698175906
transform 1 0 91504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2362
timestamp 1698175906
transform 1 0 99344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2363
timestamp 1698175906
transform 1 0 107184 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2364
timestamp 1698175906
transform 1 0 115024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2365
timestamp 1698175906
transform 1 0 122864 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2366
timestamp 1698175906
transform 1 0 130704 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2367
timestamp 1698175906
transform 1 0 138544 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2368
timestamp 1698175906
transform 1 0 146384 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2369
timestamp 1698175906
transform 1 0 154224 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2370
timestamp 1698175906
transform 1 0 162064 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2371
timestamp 1698175906
transform 1 0 169904 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2372
timestamp 1698175906
transform 1 0 177744 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2373
timestamp 1698175906
transform 1 0 185584 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2374
timestamp 1698175906
transform 1 0 193424 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2375
timestamp 1698175906
transform 1 0 201264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2376
timestamp 1698175906
transform 1 0 209104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2377
timestamp 1698175906
transform 1 0 216944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2378
timestamp 1698175906
transform 1 0 224784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2379
timestamp 1698175906
transform 1 0 232624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2380
timestamp 1698175906
transform 1 0 240464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2381
timestamp 1698175906
transform 1 0 248304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2382
timestamp 1698175906
transform 1 0 256144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2383
timestamp 1698175906
transform 1 0 263984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2384
timestamp 1698175906
transform 1 0 271824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2385
timestamp 1698175906
transform 1 0 279664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2386
timestamp 1698175906
transform 1 0 287504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2387
timestamp 1698175906
transform 1 0 295344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2388
timestamp 1698175906
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2389
timestamp 1698175906
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2390
timestamp 1698175906
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2391
timestamp 1698175906
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2392
timestamp 1698175906
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2393
timestamp 1698175906
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2394
timestamp 1698175906
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2395
timestamp 1698175906
transform 1 0 64064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2396
timestamp 1698175906
transform 1 0 71904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2397
timestamp 1698175906
transform 1 0 79744 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2398
timestamp 1698175906
transform 1 0 87584 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2399
timestamp 1698175906
transform 1 0 95424 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2400
timestamp 1698175906
transform 1 0 103264 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2401
timestamp 1698175906
transform 1 0 111104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2402
timestamp 1698175906
transform 1 0 118944 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2403
timestamp 1698175906
transform 1 0 126784 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2404
timestamp 1698175906
transform 1 0 134624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2405
timestamp 1698175906
transform 1 0 142464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2406
timestamp 1698175906
transform 1 0 150304 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2407
timestamp 1698175906
transform 1 0 158144 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2408
timestamp 1698175906
transform 1 0 165984 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2409
timestamp 1698175906
transform 1 0 173824 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2410
timestamp 1698175906
transform 1 0 181664 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2411
timestamp 1698175906
transform 1 0 189504 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2412
timestamp 1698175906
transform 1 0 197344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2413
timestamp 1698175906
transform 1 0 205184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2414
timestamp 1698175906
transform 1 0 213024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2415
timestamp 1698175906
transform 1 0 220864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2416
timestamp 1698175906
transform 1 0 228704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2417
timestamp 1698175906
transform 1 0 236544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2418
timestamp 1698175906
transform 1 0 244384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2419
timestamp 1698175906
transform 1 0 252224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2420
timestamp 1698175906
transform 1 0 260064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2421
timestamp 1698175906
transform 1 0 267904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2422
timestamp 1698175906
transform 1 0 275744 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2423
timestamp 1698175906
transform 1 0 283584 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2424
timestamp 1698175906
transform 1 0 291424 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2425
timestamp 1698175906
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2426
timestamp 1698175906
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2427
timestamp 1698175906
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2428
timestamp 1698175906
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2429
timestamp 1698175906
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2430
timestamp 1698175906
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2431
timestamp 1698175906
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2432
timestamp 1698175906
transform 1 0 60144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2433
timestamp 1698175906
transform 1 0 67984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2434
timestamp 1698175906
transform 1 0 75824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2435
timestamp 1698175906
transform 1 0 83664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2436
timestamp 1698175906
transform 1 0 91504 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2437
timestamp 1698175906
transform 1 0 99344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2438
timestamp 1698175906
transform 1 0 107184 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2439
timestamp 1698175906
transform 1 0 115024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2440
timestamp 1698175906
transform 1 0 122864 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2441
timestamp 1698175906
transform 1 0 130704 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2442
timestamp 1698175906
transform 1 0 138544 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2443
timestamp 1698175906
transform 1 0 146384 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2444
timestamp 1698175906
transform 1 0 154224 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2445
timestamp 1698175906
transform 1 0 162064 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2446
timestamp 1698175906
transform 1 0 169904 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2447
timestamp 1698175906
transform 1 0 177744 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2448
timestamp 1698175906
transform 1 0 185584 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2449
timestamp 1698175906
transform 1 0 193424 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2450
timestamp 1698175906
transform 1 0 201264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2451
timestamp 1698175906
transform 1 0 209104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2452
timestamp 1698175906
transform 1 0 216944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2453
timestamp 1698175906
transform 1 0 224784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2454
timestamp 1698175906
transform 1 0 232624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2455
timestamp 1698175906
transform 1 0 240464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2456
timestamp 1698175906
transform 1 0 248304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2457
timestamp 1698175906
transform 1 0 256144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2458
timestamp 1698175906
transform 1 0 263984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2459
timestamp 1698175906
transform 1 0 271824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2460
timestamp 1698175906
transform 1 0 279664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2461
timestamp 1698175906
transform 1 0 287504 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2462
timestamp 1698175906
transform 1 0 295344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2463
timestamp 1698175906
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2464
timestamp 1698175906
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2465
timestamp 1698175906
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2466
timestamp 1698175906
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2467
timestamp 1698175906
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2468
timestamp 1698175906
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2469
timestamp 1698175906
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2470
timestamp 1698175906
transform 1 0 64064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2471
timestamp 1698175906
transform 1 0 71904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2472
timestamp 1698175906
transform 1 0 79744 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2473
timestamp 1698175906
transform 1 0 87584 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2474
timestamp 1698175906
transform 1 0 95424 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2475
timestamp 1698175906
transform 1 0 103264 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2476
timestamp 1698175906
transform 1 0 111104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2477
timestamp 1698175906
transform 1 0 118944 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2478
timestamp 1698175906
transform 1 0 126784 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2479
timestamp 1698175906
transform 1 0 134624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2480
timestamp 1698175906
transform 1 0 142464 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2481
timestamp 1698175906
transform 1 0 150304 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2482
timestamp 1698175906
transform 1 0 158144 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2483
timestamp 1698175906
transform 1 0 165984 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2484
timestamp 1698175906
transform 1 0 173824 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2485
timestamp 1698175906
transform 1 0 181664 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2486
timestamp 1698175906
transform 1 0 189504 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2487
timestamp 1698175906
transform 1 0 197344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2488
timestamp 1698175906
transform 1 0 205184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2489
timestamp 1698175906
transform 1 0 213024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2490
timestamp 1698175906
transform 1 0 220864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2491
timestamp 1698175906
transform 1 0 228704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2492
timestamp 1698175906
transform 1 0 236544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2493
timestamp 1698175906
transform 1 0 244384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2494
timestamp 1698175906
transform 1 0 252224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2495
timestamp 1698175906
transform 1 0 260064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2496
timestamp 1698175906
transform 1 0 267904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2497
timestamp 1698175906
transform 1 0 275744 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2498
timestamp 1698175906
transform 1 0 283584 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2499
timestamp 1698175906
transform 1 0 291424 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2500
timestamp 1698175906
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2501
timestamp 1698175906
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2502
timestamp 1698175906
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2503
timestamp 1698175906
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2504
timestamp 1698175906
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2505
timestamp 1698175906
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2506
timestamp 1698175906
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2507
timestamp 1698175906
transform 1 0 60144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2508
timestamp 1698175906
transform 1 0 67984 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2509
timestamp 1698175906
transform 1 0 75824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2510
timestamp 1698175906
transform 1 0 83664 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2511
timestamp 1698175906
transform 1 0 91504 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2512
timestamp 1698175906
transform 1 0 99344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2513
timestamp 1698175906
transform 1 0 107184 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2514
timestamp 1698175906
transform 1 0 115024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2515
timestamp 1698175906
transform 1 0 122864 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2516
timestamp 1698175906
transform 1 0 130704 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2517
timestamp 1698175906
transform 1 0 138544 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2518
timestamp 1698175906
transform 1 0 146384 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2519
timestamp 1698175906
transform 1 0 154224 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2520
timestamp 1698175906
transform 1 0 162064 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2521
timestamp 1698175906
transform 1 0 169904 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2522
timestamp 1698175906
transform 1 0 177744 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2523
timestamp 1698175906
transform 1 0 185584 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2524
timestamp 1698175906
transform 1 0 193424 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2525
timestamp 1698175906
transform 1 0 201264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2526
timestamp 1698175906
transform 1 0 209104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2527
timestamp 1698175906
transform 1 0 216944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2528
timestamp 1698175906
transform 1 0 224784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2529
timestamp 1698175906
transform 1 0 232624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2530
timestamp 1698175906
transform 1 0 240464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2531
timestamp 1698175906
transform 1 0 248304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2532
timestamp 1698175906
transform 1 0 256144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2533
timestamp 1698175906
transform 1 0 263984 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2534
timestamp 1698175906
transform 1 0 271824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2535
timestamp 1698175906
transform 1 0 279664 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2536
timestamp 1698175906
transform 1 0 287504 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2537
timestamp 1698175906
transform 1 0 295344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2538
timestamp 1698175906
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2539
timestamp 1698175906
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2540
timestamp 1698175906
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2541
timestamp 1698175906
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2542
timestamp 1698175906
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2543
timestamp 1698175906
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2544
timestamp 1698175906
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2545
timestamp 1698175906
transform 1 0 64064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2546
timestamp 1698175906
transform 1 0 71904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2547
timestamp 1698175906
transform 1 0 79744 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2548
timestamp 1698175906
transform 1 0 87584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2549
timestamp 1698175906
transform 1 0 95424 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2550
timestamp 1698175906
transform 1 0 103264 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2551
timestamp 1698175906
transform 1 0 111104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2552
timestamp 1698175906
transform 1 0 118944 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2553
timestamp 1698175906
transform 1 0 126784 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2554
timestamp 1698175906
transform 1 0 134624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2555
timestamp 1698175906
transform 1 0 142464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2556
timestamp 1698175906
transform 1 0 150304 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2557
timestamp 1698175906
transform 1 0 158144 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2558
timestamp 1698175906
transform 1 0 165984 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2559
timestamp 1698175906
transform 1 0 173824 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2560
timestamp 1698175906
transform 1 0 181664 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2561
timestamp 1698175906
transform 1 0 189504 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2562
timestamp 1698175906
transform 1 0 197344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2563
timestamp 1698175906
transform 1 0 205184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2564
timestamp 1698175906
transform 1 0 213024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2565
timestamp 1698175906
transform 1 0 220864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2566
timestamp 1698175906
transform 1 0 228704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2567
timestamp 1698175906
transform 1 0 236544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2568
timestamp 1698175906
transform 1 0 244384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2569
timestamp 1698175906
transform 1 0 252224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2570
timestamp 1698175906
transform 1 0 260064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2571
timestamp 1698175906
transform 1 0 267904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2572
timestamp 1698175906
transform 1 0 275744 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2573
timestamp 1698175906
transform 1 0 283584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2574
timestamp 1698175906
transform 1 0 291424 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2575
timestamp 1698175906
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2576
timestamp 1698175906
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2577
timestamp 1698175906
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2578
timestamp 1698175906
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2579
timestamp 1698175906
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2580
timestamp 1698175906
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2581
timestamp 1698175906
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2582
timestamp 1698175906
transform 1 0 60144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2583
timestamp 1698175906
transform 1 0 67984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2584
timestamp 1698175906
transform 1 0 75824 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2585
timestamp 1698175906
transform 1 0 83664 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2586
timestamp 1698175906
transform 1 0 91504 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2587
timestamp 1698175906
transform 1 0 99344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2588
timestamp 1698175906
transform 1 0 107184 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2589
timestamp 1698175906
transform 1 0 115024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2590
timestamp 1698175906
transform 1 0 122864 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2591
timestamp 1698175906
transform 1 0 130704 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2592
timestamp 1698175906
transform 1 0 138544 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2593
timestamp 1698175906
transform 1 0 146384 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2594
timestamp 1698175906
transform 1 0 154224 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2595
timestamp 1698175906
transform 1 0 162064 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2596
timestamp 1698175906
transform 1 0 169904 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2597
timestamp 1698175906
transform 1 0 177744 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2598
timestamp 1698175906
transform 1 0 185584 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2599
timestamp 1698175906
transform 1 0 193424 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2600
timestamp 1698175906
transform 1 0 201264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2601
timestamp 1698175906
transform 1 0 209104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2602
timestamp 1698175906
transform 1 0 216944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2603
timestamp 1698175906
transform 1 0 224784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2604
timestamp 1698175906
transform 1 0 232624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2605
timestamp 1698175906
transform 1 0 240464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2606
timestamp 1698175906
transform 1 0 248304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2607
timestamp 1698175906
transform 1 0 256144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2608
timestamp 1698175906
transform 1 0 263984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2609
timestamp 1698175906
transform 1 0 271824 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2610
timestamp 1698175906
transform 1 0 279664 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2611
timestamp 1698175906
transform 1 0 287504 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2612
timestamp 1698175906
transform 1 0 295344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2613
timestamp 1698175906
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2614
timestamp 1698175906
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2615
timestamp 1698175906
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2616
timestamp 1698175906
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2617
timestamp 1698175906
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2618
timestamp 1698175906
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2619
timestamp 1698175906
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2620
timestamp 1698175906
transform 1 0 64064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2621
timestamp 1698175906
transform 1 0 71904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2622
timestamp 1698175906
transform 1 0 79744 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2623
timestamp 1698175906
transform 1 0 87584 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2624
timestamp 1698175906
transform 1 0 95424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2625
timestamp 1698175906
transform 1 0 103264 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2626
timestamp 1698175906
transform 1 0 111104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2627
timestamp 1698175906
transform 1 0 118944 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2628
timestamp 1698175906
transform 1 0 126784 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2629
timestamp 1698175906
transform 1 0 134624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2630
timestamp 1698175906
transform 1 0 142464 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2631
timestamp 1698175906
transform 1 0 150304 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2632
timestamp 1698175906
transform 1 0 158144 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2633
timestamp 1698175906
transform 1 0 165984 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2634
timestamp 1698175906
transform 1 0 173824 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2635
timestamp 1698175906
transform 1 0 181664 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2636
timestamp 1698175906
transform 1 0 189504 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2637
timestamp 1698175906
transform 1 0 197344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2638
timestamp 1698175906
transform 1 0 205184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2639
timestamp 1698175906
transform 1 0 213024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2640
timestamp 1698175906
transform 1 0 220864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2641
timestamp 1698175906
transform 1 0 228704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2642
timestamp 1698175906
transform 1 0 236544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2643
timestamp 1698175906
transform 1 0 244384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2644
timestamp 1698175906
transform 1 0 252224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2645
timestamp 1698175906
transform 1 0 260064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2646
timestamp 1698175906
transform 1 0 267904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2647
timestamp 1698175906
transform 1 0 275744 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2648
timestamp 1698175906
transform 1 0 283584 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2649
timestamp 1698175906
transform 1 0 291424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2650
timestamp 1698175906
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2651
timestamp 1698175906
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2652
timestamp 1698175906
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2653
timestamp 1698175906
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2654
timestamp 1698175906
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2655
timestamp 1698175906
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2656
timestamp 1698175906
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2657
timestamp 1698175906
transform 1 0 60144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2658
timestamp 1698175906
transform 1 0 67984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2659
timestamp 1698175906
transform 1 0 75824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2660
timestamp 1698175906
transform 1 0 83664 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2661
timestamp 1698175906
transform 1 0 91504 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2662
timestamp 1698175906
transform 1 0 99344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2663
timestamp 1698175906
transform 1 0 107184 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2664
timestamp 1698175906
transform 1 0 115024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2665
timestamp 1698175906
transform 1 0 122864 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2666
timestamp 1698175906
transform 1 0 130704 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2667
timestamp 1698175906
transform 1 0 138544 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2668
timestamp 1698175906
transform 1 0 146384 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2669
timestamp 1698175906
transform 1 0 154224 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2670
timestamp 1698175906
transform 1 0 162064 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2671
timestamp 1698175906
transform 1 0 169904 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2672
timestamp 1698175906
transform 1 0 177744 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2673
timestamp 1698175906
transform 1 0 185584 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2674
timestamp 1698175906
transform 1 0 193424 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2675
timestamp 1698175906
transform 1 0 201264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2676
timestamp 1698175906
transform 1 0 209104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2677
timestamp 1698175906
transform 1 0 216944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2678
timestamp 1698175906
transform 1 0 224784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2679
timestamp 1698175906
transform 1 0 232624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2680
timestamp 1698175906
transform 1 0 240464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2681
timestamp 1698175906
transform 1 0 248304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2682
timestamp 1698175906
transform 1 0 256144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2683
timestamp 1698175906
transform 1 0 263984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2684
timestamp 1698175906
transform 1 0 271824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2685
timestamp 1698175906
transform 1 0 279664 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2686
timestamp 1698175906
transform 1 0 287504 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2687
timestamp 1698175906
transform 1 0 295344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2688
timestamp 1698175906
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2689
timestamp 1698175906
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2690
timestamp 1698175906
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2691
timestamp 1698175906
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2692
timestamp 1698175906
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2693
timestamp 1698175906
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2694
timestamp 1698175906
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2695
timestamp 1698175906
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2696
timestamp 1698175906
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2697
timestamp 1698175906
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2698
timestamp 1698175906
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2699
timestamp 1698175906
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2700
timestamp 1698175906
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2701
timestamp 1698175906
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2702
timestamp 1698175906
transform 1 0 58464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2703
timestamp 1698175906
transform 1 0 62272 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2704
timestamp 1698175906
transform 1 0 66080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2705
timestamp 1698175906
transform 1 0 69888 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2706
timestamp 1698175906
transform 1 0 73696 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2707
timestamp 1698175906
transform 1 0 77504 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2708
timestamp 1698175906
transform 1 0 81312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2709
timestamp 1698175906
transform 1 0 85120 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2710
timestamp 1698175906
transform 1 0 88928 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2711
timestamp 1698175906
transform 1 0 92736 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2712
timestamp 1698175906
transform 1 0 96544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2713
timestamp 1698175906
transform 1 0 100352 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2714
timestamp 1698175906
transform 1 0 104160 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2715
timestamp 1698175906
transform 1 0 107968 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2716
timestamp 1698175906
transform 1 0 111776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2717
timestamp 1698175906
transform 1 0 115584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2718
timestamp 1698175906
transform 1 0 119392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2719
timestamp 1698175906
transform 1 0 123200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2720
timestamp 1698175906
transform 1 0 127008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2721
timestamp 1698175906
transform 1 0 130816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2722
timestamp 1698175906
transform 1 0 134624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2723
timestamp 1698175906
transform 1 0 138432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2724
timestamp 1698175906
transform 1 0 142240 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2725
timestamp 1698175906
transform 1 0 146048 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2726
timestamp 1698175906
transform 1 0 149856 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2727
timestamp 1698175906
transform 1 0 153664 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2728
timestamp 1698175906
transform 1 0 157472 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2729
timestamp 1698175906
transform 1 0 161280 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2730
timestamp 1698175906
transform 1 0 165088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2731
timestamp 1698175906
transform 1 0 168896 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2732
timestamp 1698175906
transform 1 0 172704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2733
timestamp 1698175906
transform 1 0 176512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2734
timestamp 1698175906
transform 1 0 180320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2735
timestamp 1698175906
transform 1 0 184128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2736
timestamp 1698175906
transform 1 0 187936 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2737
timestamp 1698175906
transform 1 0 191744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2738
timestamp 1698175906
transform 1 0 195552 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2739
timestamp 1698175906
transform 1 0 199360 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2740
timestamp 1698175906
transform 1 0 203168 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2741
timestamp 1698175906
transform 1 0 206976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2742
timestamp 1698175906
transform 1 0 210784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2743
timestamp 1698175906
transform 1 0 214592 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2744
timestamp 1698175906
transform 1 0 218400 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2745
timestamp 1698175906
transform 1 0 222208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2746
timestamp 1698175906
transform 1 0 226016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2747
timestamp 1698175906
transform 1 0 229824 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2748
timestamp 1698175906
transform 1 0 233632 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2749
timestamp 1698175906
transform 1 0 237440 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2750
timestamp 1698175906
transform 1 0 241248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2751
timestamp 1698175906
transform 1 0 245056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2752
timestamp 1698175906
transform 1 0 248864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2753
timestamp 1698175906
transform 1 0 252672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2754
timestamp 1698175906
transform 1 0 256480 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2755
timestamp 1698175906
transform 1 0 260288 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2756
timestamp 1698175906
transform 1 0 264096 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2757
timestamp 1698175906
transform 1 0 267904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2758
timestamp 1698175906
transform 1 0 271712 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2759
timestamp 1698175906
transform 1 0 275520 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2760
timestamp 1698175906
transform 1 0 279328 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2761
timestamp 1698175906
transform 1 0 283136 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2762
timestamp 1698175906
transform 1 0 286944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2763
timestamp 1698175906
transform 1 0 290752 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2764
timestamp 1698175906
transform 1 0 294560 0 -1 56448
box -86 -86 310 870
<< labels >>
flabel metal2 s 40544 0 40656 800 0 FreeSans 448 90 0 0 A_all[0]
port 0 nsew signal tristate
flabel metal2 s 44128 0 44240 800 0 FreeSans 448 90 0 0 A_all[1]
port 1 nsew signal tristate
flabel metal2 s 47712 0 47824 800 0 FreeSans 448 90 0 0 A_all[2]
port 2 nsew signal tristate
flabel metal2 s 51296 0 51408 800 0 FreeSans 448 90 0 0 A_all[3]
port 3 nsew signal tristate
flabel metal2 s 54880 0 54992 800 0 FreeSans 448 90 0 0 A_all[4]
port 4 nsew signal tristate
flabel metal2 s 58464 0 58576 800 0 FreeSans 448 90 0 0 A_all[5]
port 5 nsew signal tristate
flabel metal2 s 62048 0 62160 800 0 FreeSans 448 90 0 0 A_all[6]
port 6 nsew signal tristate
flabel metal2 s 65632 0 65744 800 0 FreeSans 448 90 0 0 A_all[7]
port 7 nsew signal tristate
flabel metal2 s 69216 0 69328 800 0 FreeSans 448 90 0 0 A_all[8]
port 8 nsew signal tristate
flabel metal2 s 8288 0 8400 800 0 FreeSans 448 90 0 0 CEN_all
port 9 nsew signal tristate
flabel metal2 s 72800 0 72912 800 0 FreeSans 448 90 0 0 D_all[0]
port 10 nsew signal tristate
flabel metal2 s 76384 0 76496 800 0 FreeSans 448 90 0 0 D_all[1]
port 11 nsew signal tristate
flabel metal2 s 79968 0 80080 800 0 FreeSans 448 90 0 0 D_all[2]
port 12 nsew signal tristate
flabel metal2 s 83552 0 83664 800 0 FreeSans 448 90 0 0 D_all[3]
port 13 nsew signal tristate
flabel metal2 s 87136 0 87248 800 0 FreeSans 448 90 0 0 D_all[4]
port 14 nsew signal tristate
flabel metal2 s 90720 0 90832 800 0 FreeSans 448 90 0 0 D_all[5]
port 15 nsew signal tristate
flabel metal2 s 94304 0 94416 800 0 FreeSans 448 90 0 0 D_all[6]
port 16 nsew signal tristate
flabel metal2 s 97888 0 98000 800 0 FreeSans 448 90 0 0 D_all[7]
port 17 nsew signal tristate
flabel metal2 s 101472 0 101584 800 0 FreeSans 448 90 0 0 GWEN_0
port 18 nsew signal tristate
flabel metal2 s 105056 0 105168 800 0 FreeSans 448 90 0 0 GWEN_1
port 19 nsew signal tristate
flabel metal2 s 108640 0 108752 800 0 FreeSans 448 90 0 0 GWEN_2
port 20 nsew signal tristate
flabel metal2 s 112224 0 112336 800 0 FreeSans 448 90 0 0 GWEN_3
port 21 nsew signal tristate
flabel metal2 s 115808 0 115920 800 0 FreeSans 448 90 0 0 GWEN_4
port 22 nsew signal tristate
flabel metal2 s 119392 0 119504 800 0 FreeSans 448 90 0 0 GWEN_5
port 23 nsew signal tristate
flabel metal2 s 200928 59200 201040 60000 0 FreeSans 448 90 0 0 GWEN_6
port 24 nsew signal tristate
flabel metal2 s 206304 59200 206416 60000 0 FreeSans 448 90 0 0 GWEN_7
port 25 nsew signal tristate
flabel metal2 s 122976 0 123088 800 0 FreeSans 448 90 0 0 Q0[0]
port 26 nsew signal input
flabel metal2 s 126560 0 126672 800 0 FreeSans 448 90 0 0 Q0[1]
port 27 nsew signal input
flabel metal2 s 130144 0 130256 800 0 FreeSans 448 90 0 0 Q0[2]
port 28 nsew signal input
flabel metal2 s 133728 0 133840 800 0 FreeSans 448 90 0 0 Q0[3]
port 29 nsew signal input
flabel metal2 s 137312 0 137424 800 0 FreeSans 448 90 0 0 Q0[4]
port 30 nsew signal input
flabel metal2 s 140896 0 141008 800 0 FreeSans 448 90 0 0 Q0[5]
port 31 nsew signal input
flabel metal2 s 144480 0 144592 800 0 FreeSans 448 90 0 0 Q0[6]
port 32 nsew signal input
flabel metal2 s 148064 0 148176 800 0 FreeSans 448 90 0 0 Q0[7]
port 33 nsew signal input
flabel metal2 s 151648 0 151760 800 0 FreeSans 448 90 0 0 Q1[0]
port 34 nsew signal input
flabel metal2 s 155232 0 155344 800 0 FreeSans 448 90 0 0 Q1[1]
port 35 nsew signal input
flabel metal2 s 158816 0 158928 800 0 FreeSans 448 90 0 0 Q1[2]
port 36 nsew signal input
flabel metal2 s 162400 0 162512 800 0 FreeSans 448 90 0 0 Q1[3]
port 37 nsew signal input
flabel metal2 s 165984 0 166096 800 0 FreeSans 448 90 0 0 Q1[4]
port 38 nsew signal input
flabel metal2 s 169568 0 169680 800 0 FreeSans 448 90 0 0 Q1[5]
port 39 nsew signal input
flabel metal2 s 173152 0 173264 800 0 FreeSans 448 90 0 0 Q1[6]
port 40 nsew signal input
flabel metal2 s 176736 0 176848 800 0 FreeSans 448 90 0 0 Q1[7]
port 41 nsew signal input
flabel metal2 s 180320 0 180432 800 0 FreeSans 448 90 0 0 Q2[0]
port 42 nsew signal input
flabel metal2 s 183904 0 184016 800 0 FreeSans 448 90 0 0 Q2[1]
port 43 nsew signal input
flabel metal2 s 187488 0 187600 800 0 FreeSans 448 90 0 0 Q2[2]
port 44 nsew signal input
flabel metal2 s 191072 0 191184 800 0 FreeSans 448 90 0 0 Q2[3]
port 45 nsew signal input
flabel metal2 s 194656 0 194768 800 0 FreeSans 448 90 0 0 Q2[4]
port 46 nsew signal input
flabel metal2 s 198240 0 198352 800 0 FreeSans 448 90 0 0 Q2[5]
port 47 nsew signal input
flabel metal2 s 201824 0 201936 800 0 FreeSans 448 90 0 0 Q2[6]
port 48 nsew signal input
flabel metal2 s 205408 0 205520 800 0 FreeSans 448 90 0 0 Q2[7]
port 49 nsew signal input
flabel metal2 s 208992 0 209104 800 0 FreeSans 448 90 0 0 Q3[0]
port 50 nsew signal input
flabel metal2 s 212576 0 212688 800 0 FreeSans 448 90 0 0 Q3[1]
port 51 nsew signal input
flabel metal2 s 216160 0 216272 800 0 FreeSans 448 90 0 0 Q3[2]
port 52 nsew signal input
flabel metal2 s 219744 0 219856 800 0 FreeSans 448 90 0 0 Q3[3]
port 53 nsew signal input
flabel metal2 s 223328 0 223440 800 0 FreeSans 448 90 0 0 Q3[4]
port 54 nsew signal input
flabel metal2 s 226912 0 227024 800 0 FreeSans 448 90 0 0 Q3[5]
port 55 nsew signal input
flabel metal2 s 230496 0 230608 800 0 FreeSans 448 90 0 0 Q3[6]
port 56 nsew signal input
flabel metal2 s 234080 0 234192 800 0 FreeSans 448 90 0 0 Q3[7]
port 57 nsew signal input
flabel metal2 s 237664 0 237776 800 0 FreeSans 448 90 0 0 Q4[0]
port 58 nsew signal input
flabel metal2 s 241248 0 241360 800 0 FreeSans 448 90 0 0 Q4[1]
port 59 nsew signal input
flabel metal2 s 244832 0 244944 800 0 FreeSans 448 90 0 0 Q4[2]
port 60 nsew signal input
flabel metal2 s 248416 0 248528 800 0 FreeSans 448 90 0 0 Q4[3]
port 61 nsew signal input
flabel metal2 s 252000 0 252112 800 0 FreeSans 448 90 0 0 Q4[4]
port 62 nsew signal input
flabel metal2 s 255584 0 255696 800 0 FreeSans 448 90 0 0 Q4[5]
port 63 nsew signal input
flabel metal2 s 259168 0 259280 800 0 FreeSans 448 90 0 0 Q4[6]
port 64 nsew signal input
flabel metal2 s 262752 0 262864 800 0 FreeSans 448 90 0 0 Q4[7]
port 65 nsew signal input
flabel metal2 s 266336 0 266448 800 0 FreeSans 448 90 0 0 Q5[0]
port 66 nsew signal input
flabel metal2 s 269920 0 270032 800 0 FreeSans 448 90 0 0 Q5[1]
port 67 nsew signal input
flabel metal2 s 273504 0 273616 800 0 FreeSans 448 90 0 0 Q5[2]
port 68 nsew signal input
flabel metal2 s 277088 0 277200 800 0 FreeSans 448 90 0 0 Q5[3]
port 69 nsew signal input
flabel metal2 s 280672 0 280784 800 0 FreeSans 448 90 0 0 Q5[4]
port 70 nsew signal input
flabel metal2 s 284256 0 284368 800 0 FreeSans 448 90 0 0 Q5[5]
port 71 nsew signal input
flabel metal2 s 287840 0 287952 800 0 FreeSans 448 90 0 0 Q5[6]
port 72 nsew signal input
flabel metal2 s 291424 0 291536 800 0 FreeSans 448 90 0 0 Q5[7]
port 73 nsew signal input
flabel metal2 s 211680 59200 211792 60000 0 FreeSans 448 90 0 0 Q6[0]
port 74 nsew signal input
flabel metal2 s 217056 59200 217168 60000 0 FreeSans 448 90 0 0 Q6[1]
port 75 nsew signal input
flabel metal2 s 222432 59200 222544 60000 0 FreeSans 448 90 0 0 Q6[2]
port 76 nsew signal input
flabel metal2 s 227808 59200 227920 60000 0 FreeSans 448 90 0 0 Q6[3]
port 77 nsew signal input
flabel metal2 s 233184 59200 233296 60000 0 FreeSans 448 90 0 0 Q6[4]
port 78 nsew signal input
flabel metal2 s 238560 59200 238672 60000 0 FreeSans 448 90 0 0 Q6[5]
port 79 nsew signal input
flabel metal2 s 243936 59200 244048 60000 0 FreeSans 448 90 0 0 Q6[6]
port 80 nsew signal input
flabel metal2 s 249312 59200 249424 60000 0 FreeSans 448 90 0 0 Q6[7]
port 81 nsew signal input
flabel metal2 s 254688 59200 254800 60000 0 FreeSans 448 90 0 0 Q7[0]
port 82 nsew signal input
flabel metal2 s 260064 59200 260176 60000 0 FreeSans 448 90 0 0 Q7[1]
port 83 nsew signal input
flabel metal2 s 265440 59200 265552 60000 0 FreeSans 448 90 0 0 Q7[2]
port 84 nsew signal input
flabel metal2 s 270816 59200 270928 60000 0 FreeSans 448 90 0 0 Q7[3]
port 85 nsew signal input
flabel metal2 s 276192 59200 276304 60000 0 FreeSans 448 90 0 0 Q7[4]
port 86 nsew signal input
flabel metal2 s 281568 59200 281680 60000 0 FreeSans 448 90 0 0 Q7[5]
port 87 nsew signal input
flabel metal2 s 286944 59200 287056 60000 0 FreeSans 448 90 0 0 Q7[6]
port 88 nsew signal input
flabel metal2 s 292320 59200 292432 60000 0 FreeSans 448 90 0 0 Q7[7]
port 89 nsew signal input
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 WEN_all[0]
port 90 nsew signal tristate
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 WEN_all[1]
port 91 nsew signal tristate
flabel metal2 s 19040 0 19152 800 0 FreeSans 448 90 0 0 WEN_all[2]
port 92 nsew signal tristate
flabel metal2 s 22624 0 22736 800 0 FreeSans 448 90 0 0 WEN_all[3]
port 93 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 WEN_all[4]
port 94 nsew signal tristate
flabel metal2 s 29792 0 29904 800 0 FreeSans 448 90 0 0 WEN_all[5]
port 95 nsew signal tristate
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 WEN_all[6]
port 96 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 WEN_all[7]
port 97 nsew signal tristate
flabel metal2 s 18144 59200 18256 60000 0 FreeSans 448 90 0 0 WEb_raw
port 98 nsew signal input
flabel metal2 s 23520 59200 23632 60000 0 FreeSans 448 90 0 0 bus_in[0]
port 99 nsew signal input
flabel metal2 s 28896 59200 29008 60000 0 FreeSans 448 90 0 0 bus_in[1]
port 100 nsew signal input
flabel metal2 s 34272 59200 34384 60000 0 FreeSans 448 90 0 0 bus_in[2]
port 101 nsew signal input
flabel metal2 s 39648 59200 39760 60000 0 FreeSans 448 90 0 0 bus_in[3]
port 102 nsew signal input
flabel metal2 s 45024 59200 45136 60000 0 FreeSans 448 90 0 0 bus_in[4]
port 103 nsew signal input
flabel metal2 s 50400 59200 50512 60000 0 FreeSans 448 90 0 0 bus_in[5]
port 104 nsew signal input
flabel metal2 s 55776 59200 55888 60000 0 FreeSans 448 90 0 0 bus_in[6]
port 105 nsew signal input
flabel metal2 s 61152 59200 61264 60000 0 FreeSans 448 90 0 0 bus_in[7]
port 106 nsew signal input
flabel metal2 s 66528 59200 66640 60000 0 FreeSans 448 90 0 0 bus_out[0]
port 107 nsew signal tristate
flabel metal2 s 71904 59200 72016 60000 0 FreeSans 448 90 0 0 bus_out[1]
port 108 nsew signal tristate
flabel metal2 s 77280 59200 77392 60000 0 FreeSans 448 90 0 0 bus_out[2]
port 109 nsew signal tristate
flabel metal2 s 82656 59200 82768 60000 0 FreeSans 448 90 0 0 bus_out[3]
port 110 nsew signal tristate
flabel metal2 s 88032 59200 88144 60000 0 FreeSans 448 90 0 0 bus_out[4]
port 111 nsew signal tristate
flabel metal2 s 93408 59200 93520 60000 0 FreeSans 448 90 0 0 bus_out[5]
port 112 nsew signal tristate
flabel metal2 s 98784 59200 98896 60000 0 FreeSans 448 90 0 0 bus_out[6]
port 113 nsew signal tristate
flabel metal2 s 104160 59200 104272 60000 0 FreeSans 448 90 0 0 bus_out[7]
port 114 nsew signal tristate
flabel metal2 s 109536 59200 109648 60000 0 FreeSans 448 90 0 0 ram_enabled
port 115 nsew signal input
flabel metal2 s 114912 59200 115024 60000 0 FreeSans 448 90 0 0 requested_addr[0]
port 116 nsew signal input
flabel metal2 s 168672 59200 168784 60000 0 FreeSans 448 90 0 0 requested_addr[10]
port 117 nsew signal input
flabel metal2 s 174048 59200 174160 60000 0 FreeSans 448 90 0 0 requested_addr[11]
port 118 nsew signal input
flabel metal2 s 179424 59200 179536 60000 0 FreeSans 448 90 0 0 requested_addr[12]
port 119 nsew signal input
flabel metal2 s 184800 59200 184912 60000 0 FreeSans 448 90 0 0 requested_addr[13]
port 120 nsew signal input
flabel metal2 s 190176 59200 190288 60000 0 FreeSans 448 90 0 0 requested_addr[14]
port 121 nsew signal input
flabel metal2 s 195552 59200 195664 60000 0 FreeSans 448 90 0 0 requested_addr[15]
port 122 nsew signal input
flabel metal2 s 120288 59200 120400 60000 0 FreeSans 448 90 0 0 requested_addr[1]
port 123 nsew signal input
flabel metal2 s 125664 59200 125776 60000 0 FreeSans 448 90 0 0 requested_addr[2]
port 124 nsew signal input
flabel metal2 s 131040 59200 131152 60000 0 FreeSans 448 90 0 0 requested_addr[3]
port 125 nsew signal input
flabel metal2 s 136416 59200 136528 60000 0 FreeSans 448 90 0 0 requested_addr[4]
port 126 nsew signal input
flabel metal2 s 141792 59200 141904 60000 0 FreeSans 448 90 0 0 requested_addr[5]
port 127 nsew signal input
flabel metal2 s 147168 59200 147280 60000 0 FreeSans 448 90 0 0 requested_addr[6]
port 128 nsew signal input
flabel metal2 s 152544 59200 152656 60000 0 FreeSans 448 90 0 0 requested_addr[7]
port 129 nsew signal input
flabel metal2 s 157920 59200 158032 60000 0 FreeSans 448 90 0 0 requested_addr[8]
port 130 nsew signal input
flabel metal2 s 163296 59200 163408 60000 0 FreeSans 448 90 0 0 requested_addr[9]
port 131 nsew signal input
flabel metal2 s 12768 59200 12880 60000 0 FreeSans 448 90 0 0 rst
port 132 nsew signal input
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 65888 3076 66208 56508 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 96608 3076 96928 56508 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 127328 3076 127648 56508 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 158048 3076 158368 56508 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 188768 3076 189088 56508 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 219488 3076 219808 56508 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 250208 3076 250528 56508 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 280928 3076 281248 56508 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 81248 3076 81568 56508 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 111968 3076 112288 56508 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 142688 3076 143008 56508 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 173408 3076 173728 56508 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 204128 3076 204448 56508 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 234848 3076 235168 56508 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 265568 3076 265888 56508 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 296288 3076 296608 56508 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal2 s 7392 59200 7504 60000 0 FreeSans 448 90 0 0 wb_clk_i
port 135 nsew signal input
rlabel metal1 149968 55664 149968 55664 0 vdd
rlabel metal1 149968 56448 149968 56448 0 vss
rlabel metal2 40600 2198 40600 2198 0 A_all[0]
rlabel metal2 44184 2198 44184 2198 0 A_all[1]
rlabel metal2 47768 2198 47768 2198 0 A_all[2]
rlabel metal2 51352 2198 51352 2198 0 A_all[3]
rlabel metal2 54936 2198 54936 2198 0 A_all[4]
rlabel metal2 58520 2198 58520 2198 0 A_all[5]
rlabel metal2 62104 2198 62104 2198 0 A_all[6]
rlabel metal2 65688 2086 65688 2086 0 A_all[7]
rlabel metal2 69272 2198 69272 2198 0 A_all[8]
rlabel metal2 8344 2086 8344 2086 0 CEN_all
rlabel metal2 72856 1190 72856 1190 0 D_all[0]
rlabel metal2 76440 2422 76440 2422 0 D_all[1]
rlabel metal2 80024 2422 80024 2422 0 D_all[2]
rlabel metal2 83608 2422 83608 2422 0 D_all[3]
rlabel metal2 87192 2478 87192 2478 0 D_all[4]
rlabel metal2 90776 2422 90776 2422 0 D_all[5]
rlabel metal2 94360 2030 94360 2030 0 D_all[6]
rlabel metal2 97944 854 97944 854 0 D_all[7]
rlabel metal2 101528 2198 101528 2198 0 GWEN_0
rlabel metal2 105112 2198 105112 2198 0 GWEN_1
rlabel metal2 108696 854 108696 854 0 GWEN_2
rlabel metal2 112280 1190 112280 1190 0 GWEN_3
rlabel metal2 115864 2198 115864 2198 0 GWEN_4
rlabel metal2 119448 2198 119448 2198 0 GWEN_5
rlabel metal2 200984 57610 200984 57610 0 GWEN_6
rlabel metal2 206360 57778 206360 57778 0 GWEN_7
rlabel metal2 123088 3416 123088 3416 0 Q0[0]
rlabel metal2 126952 2800 126952 2800 0 Q0[1]
rlabel metal2 130760 2800 130760 2800 0 Q0[2]
rlabel metal2 133784 2086 133784 2086 0 Q0[3]
rlabel metal2 137368 2086 137368 2086 0 Q0[4]
rlabel metal2 140952 2086 140952 2086 0 Q0[5]
rlabel metal2 144536 2086 144536 2086 0 Q0[6]
rlabel metal2 148120 2086 148120 2086 0 Q0[7]
rlabel metal2 151704 2086 151704 2086 0 Q1[0]
rlabel metal2 155288 2086 155288 2086 0 Q1[1]
rlabel metal2 158872 2086 158872 2086 0 Q1[2]
rlabel metal2 162456 2086 162456 2086 0 Q1[3]
rlabel metal2 166040 2086 166040 2086 0 Q1[4]
rlabel metal2 169624 2086 169624 2086 0 Q1[5]
rlabel metal2 173208 2086 173208 2086 0 Q1[6]
rlabel metal2 176624 3416 176624 3416 0 Q1[7]
rlabel metal2 180320 3416 180320 3416 0 Q2[0]
rlabel metal2 183736 3024 183736 3024 0 Q2[1]
rlabel metal2 187880 2800 187880 2800 0 Q2[2]
rlabel metal2 191184 3416 191184 3416 0 Q2[3]
rlabel metal3 195328 3416 195328 3416 0 Q2[4]
rlabel metal2 198856 2800 198856 2800 0 Q2[5]
rlabel metal2 206136 3696 206136 3696 0 Q2[6]
rlabel metal2 208488 4592 208488 4592 0 Q2[7]
rlabel metal2 210056 3472 210056 3472 0 Q3[0]
rlabel metal2 212632 2086 212632 2086 0 Q3[1]
rlabel metal1 215824 3752 215824 3752 0 Q3[2]
rlabel metal2 219800 2058 219800 2058 0 Q3[3]
rlabel metal2 223608 3528 223608 3528 0 Q3[4]
rlabel metal2 226968 2086 226968 2086 0 Q3[5]
rlabel metal2 230552 2086 230552 2086 0 Q3[6]
rlabel metal2 233576 2800 233576 2800 0 Q3[7]
rlabel metal2 237384 2800 237384 2800 0 Q4[0]
rlabel metal2 241248 3416 241248 3416 0 Q4[1]
rlabel metal2 244944 3416 244944 3416 0 Q4[2]
rlabel metal2 248640 3416 248640 3416 0 Q4[3]
rlabel metal2 252616 2800 252616 2800 0 Q4[4]
rlabel metal2 255640 2086 255640 2086 0 Q4[5]
rlabel metal2 259224 2086 259224 2086 0 Q4[6]
rlabel metal2 262808 2086 262808 2086 0 Q4[7]
rlabel metal2 266392 2086 266392 2086 0 Q5[0]
rlabel metal2 269976 2086 269976 2086 0 Q5[1]
rlabel metal2 273560 2086 273560 2086 0 Q5[2]
rlabel metal2 277144 2086 277144 2086 0 Q5[3]
rlabel metal2 280728 2086 280728 2086 0 Q5[4]
rlabel metal2 284312 2086 284312 2086 0 Q5[5]
rlabel metal2 287896 2086 287896 2086 0 Q5[6]
rlabel metal2 291480 2086 291480 2086 0 Q5[7]
rlabel metal2 211736 57778 211736 57778 0 Q6[0]
rlabel metal2 217112 57778 217112 57778 0 Q6[1]
rlabel metal2 222152 56728 222152 56728 0 Q6[2]
rlabel metal2 227864 57778 227864 57778 0 Q6[3]
rlabel metal2 233408 56280 233408 56280 0 Q6[4]
rlabel metal2 238616 57778 238616 57778 0 Q6[5]
rlabel metal2 243992 57778 243992 57778 0 Q6[6]
rlabel metal2 249480 56280 249480 56280 0 Q6[7]
rlabel metal2 254744 57778 254744 57778 0 Q7[0]
rlabel metal2 260120 57778 260120 57778 0 Q7[1]
rlabel metal2 265496 57778 265496 57778 0 Q7[2]
rlabel metal2 271544 56672 271544 56672 0 Q7[3]
rlabel metal2 276248 57778 276248 57778 0 Q7[4]
rlabel metal3 282184 56056 282184 56056 0 Q7[5]
rlabel metal2 286944 56280 286944 56280 0 Q7[6]
rlabel metal2 292376 57778 292376 57778 0 Q7[7]
rlabel metal2 18200 57778 18200 57778 0 WEb_raw
rlabel metal3 188552 56168 188552 56168 0 _000_
rlabel metal3 189952 8232 189952 8232 0 _001_
rlabel metal2 186760 3920 186760 3920 0 _002_
rlabel metal2 203448 8120 203448 8120 0 _003_
rlabel metal3 207032 8904 207032 8904 0 _004_
rlabel metal2 204680 7896 204680 7896 0 _005_
rlabel metal2 205800 5712 205800 5712 0 _006_
rlabel metal2 207368 7784 207368 7784 0 _007_
rlabel metal2 209832 7896 209832 7896 0 _008_
rlabel metal2 195328 4536 195328 4536 0 _009_
rlabel metal2 184632 5096 184632 5096 0 _010_
rlabel metal2 205576 6664 205576 6664 0 _011_
rlabel metal2 206472 5432 206472 5432 0 _012_
rlabel metal3 205464 4312 205464 4312 0 _013_
rlabel metal2 200872 8176 200872 8176 0 _014_
rlabel metal2 208824 5320 208824 5320 0 _015_
rlabel metal3 210616 4312 210616 4312 0 _016_
rlabel metal2 208712 3696 208712 3696 0 _017_
rlabel metal2 202888 7112 202888 7112 0 _018_
rlabel metal2 188888 4704 188888 4704 0 _019_
rlabel metal2 209496 6608 209496 6608 0 _020_
rlabel metal3 210336 4424 210336 4424 0 _021_
rlabel metal2 210392 7784 210392 7784 0 _022_
rlabel metal2 214536 7392 214536 7392 0 _023_
rlabel metal2 214088 7504 214088 7504 0 _024_
rlabel metal2 212520 9688 212520 9688 0 _025_
rlabel metal2 189392 4536 189392 4536 0 _026_
rlabel metal2 190680 5152 190680 5152 0 _027_
rlabel metal3 212352 9128 212352 9128 0 _028_
rlabel metal2 211120 8008 211120 8008 0 _029_
rlabel metal3 193592 5880 193592 5880 0 _030_
rlabel metal2 192360 5152 192360 5152 0 _031_
rlabel metal2 182392 5208 182392 5208 0 _032_
rlabel metal2 189896 4816 189896 4816 0 _033_
rlabel metal2 213864 6776 213864 6776 0 _034_
rlabel metal2 213640 5712 213640 5712 0 _035_
rlabel metal3 208908 5096 208908 5096 0 _036_
rlabel metal2 209160 4088 209160 4088 0 _037_
rlabel metal2 215208 5544 215208 5544 0 _038_
rlabel metal2 209944 5040 209944 5040 0 _039_
rlabel metal2 210280 5600 210280 5600 0 _040_
rlabel metal2 186760 6776 186760 6776 0 _041_
rlabel metal3 183288 4312 183288 4312 0 _042_
rlabel metal2 186200 4592 186200 4592 0 _043_
rlabel metal2 211624 5600 211624 5600 0 _044_
rlabel metal2 211400 4760 211400 4760 0 _045_
rlabel metal2 215320 5544 215320 5544 0 _046_
rlabel metal2 210840 7140 210840 7140 0 _047_
rlabel metal2 186760 2744 186760 2744 0 _048_
rlabel metal2 182448 3752 182448 3752 0 _049_
rlabel metal2 187432 5880 187432 5880 0 _050_
rlabel metal3 202384 4424 202384 4424 0 _051_
rlabel metal2 212856 4368 212856 4368 0 _052_
rlabel metal2 212520 4648 212520 4648 0 _053_
rlabel metal2 212632 4760 212632 4760 0 _054_
rlabel metal2 214536 4760 214536 4760 0 _055_
rlabel metal2 212408 4760 212408 4760 0 _056_
rlabel metal2 212184 7952 212184 7952 0 _057_
rlabel metal2 212296 6776 212296 6776 0 _058_
rlabel metal2 187096 3696 187096 3696 0 _059_
rlabel metal2 190904 5096 190904 5096 0 _060_
rlabel metal2 193816 4200 193816 4200 0 _061_
rlabel metal2 199192 6272 199192 6272 0 _062_
rlabel metal2 197960 4760 197960 4760 0 _063_
rlabel metal2 201096 5152 201096 5152 0 _064_
rlabel metal2 195160 6272 195160 6272 0 _065_
rlabel metal2 201712 5096 201712 5096 0 _066_
rlabel metal3 203000 3528 203000 3528 0 _067_
rlabel metal2 219184 2744 219184 2744 0 _068_
rlabel metal3 217168 4424 217168 4424 0 _069_
rlabel metal2 220024 4592 220024 4592 0 _070_
rlabel metal2 218568 5768 218568 5768 0 _071_
rlabel metal3 221760 4200 221760 4200 0 _072_
rlabel metal3 218456 9240 218456 9240 0 _073_
rlabel metal2 218064 9016 218064 9016 0 _074_
rlabel metal2 220584 6384 220584 6384 0 _075_
rlabel metal2 196112 7672 196112 7672 0 _076_
rlabel metal2 193144 4200 193144 4200 0 _077_
rlabel metal2 194824 4200 194824 4200 0 _078_
rlabel metal2 203224 3248 203224 3248 0 _079_
rlabel metal2 220808 4032 220808 4032 0 _080_
rlabel metal2 221816 4480 221816 4480 0 _081_
rlabel metal2 221368 6384 221368 6384 0 _082_
rlabel metal2 197624 2744 197624 2744 0 _083_
rlabel metal3 192360 5992 192360 5992 0 _084_
rlabel metal2 195384 5992 195384 5992 0 _085_
rlabel metal3 220248 4424 220248 4424 0 _086_
rlabel metal2 221704 4368 221704 4368 0 _087_
rlabel metal3 222824 5096 222824 5096 0 _088_
rlabel metal2 221144 6664 221144 6664 0 _089_
rlabel metal2 196112 6664 196112 6664 0 _090_
rlabel metal2 192920 5320 192920 5320 0 _091_
rlabel metal2 195384 8344 195384 8344 0 _092_
rlabel metal2 204120 5712 204120 5712 0 _093_
rlabel metal2 217448 4592 217448 4592 0 _094_
rlabel metal2 217784 5040 217784 5040 0 _095_
rlabel metal2 218008 6944 218008 6944 0 _096_
rlabel metal2 196056 9520 196056 9520 0 _097_
rlabel metal2 184520 7056 184520 7056 0 _098_
rlabel metal2 187880 7728 187880 7728 0 _099_
rlabel metal2 206136 6328 206136 6328 0 _100_
rlabel metal2 216552 6608 216552 6608 0 _101_
rlabel metal2 217784 7112 217784 7112 0 _102_
rlabel metal2 216216 8176 216216 8176 0 _103_
rlabel metal3 189616 7560 189616 7560 0 _104_
rlabel metal2 186704 55160 186704 55160 0 _105_
rlabel metal2 189336 52472 189336 52472 0 aaaa\[0\]
rlabel metal3 184296 55384 184296 55384 0 aaaa\[12\]
rlabel metal2 186144 54376 186144 54376 0 aaaa\[13\]
rlabel metal3 187376 55384 187376 55384 0 aaaa\[14\]
rlabel metal3 191352 56056 191352 56056 0 aaaa\[15\]
rlabel metal3 194544 53816 194544 53816 0 aaaa\[1\]
rlabel metal2 185416 36064 185416 36064 0 aaaa\[2\]
rlabel metal2 24136 56448 24136 56448 0 bus_in[0]
rlabel metal2 28952 57778 28952 57778 0 bus_in[1]
rlabel metal2 34328 57778 34328 57778 0 bus_in[2]
rlabel metal2 39816 56280 39816 56280 0 bus_in[3]
rlabel metal2 45080 57778 45080 57778 0 bus_in[4]
rlabel metal2 50624 56280 50624 56280 0 bus_in[5]
rlabel metal2 55832 57778 55832 57778 0 bus_in[6]
rlabel metal2 61208 57778 61208 57778 0 bus_in[7]
rlabel metal2 67032 56728 67032 56728 0 bus_out[0]
rlabel metal2 72408 55412 72408 55412 0 bus_out[1]
rlabel metal2 77336 58170 77336 58170 0 bus_out[2]
rlabel metal2 82712 57610 82712 57610 0 bus_out[3]
rlabel metal2 88088 57610 88088 57610 0 bus_out[4]
rlabel metal2 93464 57610 93464 57610 0 bus_out[5]
rlabel metal3 99456 55384 99456 55384 0 bus_out[6]
rlabel metal2 104216 57610 104216 57610 0 bus_out[7]
rlabel metal2 166264 54320 166264 54320 0 clknet_0_wb_clk_i
rlabel metal3 139440 55272 139440 55272 0 clknet_1_0__leaf_wb_clk_i
rlabel metal3 170072 55272 170072 55272 0 clknet_1_1__leaf_wb_clk_i
rlabel metal2 123928 3752 123928 3752 0 net1
rlabel metal2 156296 2912 156296 2912 0 net10
rlabel metal2 72856 3584 72856 3584 0 net100
rlabel metal2 11592 3976 11592 3976 0 net101
rlabel metal2 71736 3976 71736 3976 0 net102
rlabel metal2 75432 4368 75432 4368 0 net103
rlabel metal2 79016 3864 79016 3864 0 net104
rlabel metal2 83496 4368 83496 4368 0 net105
rlabel metal2 87080 4368 87080 4368 0 net106
rlabel metal2 89656 3864 89656 3864 0 net107
rlabel metal2 94248 3976 94248 3976 0 net108
rlabel metal3 97216 4424 97216 4424 0 net109
rlabel metal2 159656 2688 159656 2688 0 net11
rlabel metal3 106120 3416 106120 3416 0 net110
rlabel metal3 108976 3416 108976 3416 0 net111
rlabel metal2 186872 3192 186872 3192 0 net112
rlabel metal3 119728 3528 119728 3528 0 net113
rlabel metal2 118664 3584 118664 3584 0 net114
rlabel metal2 122584 4816 122584 4816 0 net115
rlabel metal2 210056 19600 210056 19600 0 net116
rlabel metal2 189336 7616 189336 7616 0 net117
rlabel metal3 71792 55944 71792 55944 0 net118
rlabel metal2 74760 55160 74760 55160 0 net119
rlabel metal2 163016 3080 163016 3080 0 net12
rlabel metal3 82096 55944 82096 55944 0 net120
rlabel metal2 192696 7980 192696 7980 0 net121
rlabel metal2 193368 2912 193368 2912 0 net122
rlabel metal3 98560 55944 98560 55944 0 net123
rlabel metal2 102312 55160 102312 55160 0 net124
rlabel metal3 183848 7560 183848 7560 0 net125
rlabel metal2 11928 2030 11928 2030 0 net126
rlabel metal2 15512 2030 15512 2030 0 net127
rlabel metal2 19096 2030 19096 2030 0 net128
rlabel metal2 22680 2030 22680 2030 0 net129
rlabel metal2 169960 3080 169960 3080 0 net13
rlabel metal2 26264 2030 26264 2030 0 net130
rlabel metal2 29848 2030 29848 2030 0 net131
rlabel metal2 33432 2030 33432 2030 0 net132
rlabel metal2 37016 2030 37016 2030 0 net133
rlabel metal2 170184 3640 170184 3640 0 net14
rlabel metal2 173768 3976 173768 3976 0 net15
rlabel metal2 177352 2240 177352 2240 0 net16
rlabel metal2 189896 3976 189896 3976 0 net17
rlabel metal2 187544 4424 187544 4424 0 net18
rlabel metal2 187768 6496 187768 6496 0 net19
rlabel metal2 127736 3472 127736 3472 0 net2
rlabel metal2 191632 3416 191632 3416 0 net20
rlabel metal2 196280 4256 196280 4256 0 net21
rlabel metal2 198184 5880 198184 5880 0 net22
rlabel metal2 201152 6664 201152 6664 0 net23
rlabel metal2 206360 5880 206360 5880 0 net24
rlabel metal2 209832 3360 209832 3360 0 net25
rlabel metal3 212128 3416 212128 3416 0 net26
rlabel metal2 212296 3920 212296 3920 0 net27
rlabel metal2 219912 3864 219912 3864 0 net28
rlabel metal2 223776 3304 223776 3304 0 net29
rlabel metal2 131544 3584 131544 3584 0 net3
rlabel metal3 227192 3360 227192 3360 0 net30
rlabel metal2 230776 3920 230776 3920 0 net31
rlabel metal2 234360 4536 234360 4536 0 net32
rlabel metal2 237944 3528 237944 3528 0 net33
rlabel metal2 241640 4144 241640 4144 0 net34
rlabel metal3 231840 5264 231840 5264 0 net35
rlabel metal2 249256 3864 249256 3864 0 net36
rlabel metal2 253064 3696 253064 3696 0 net37
rlabel metal2 255864 3528 255864 3528 0 net38
rlabel metal2 259448 3024 259448 3024 0 net39
rlabel metal2 190456 3416 190456 3416 0 net4
rlabel metal2 263032 4704 263032 4704 0 net40
rlabel metal2 195832 2912 195832 2912 0 net41
rlabel metal2 195496 5264 195496 5264 0 net42
rlabel metal3 192976 6440 192976 6440 0 net43
rlabel metal2 208040 4816 208040 4816 0 net44
rlabel metal2 281400 3696 281400 3696 0 net45
rlabel metal2 204904 5208 204904 5208 0 net46
rlabel metal2 288568 4032 288568 4032 0 net47
rlabel metal3 206080 6664 206080 6664 0 net48
rlabel metal3 212128 8120 212128 8120 0 net49
rlabel metal2 137928 5544 137928 5544 0 net5
rlabel metal2 211960 11256 211960 11256 0 net50
rlabel metal3 212912 8232 212912 8232 0 net51
rlabel metal3 226184 53816 226184 53816 0 net52
rlabel metal2 234024 55048 234024 55048 0 net53
rlabel metal2 239288 55272 239288 55272 0 net54
rlabel metal2 244776 33600 244776 33600 0 net55
rlabel metal2 250152 34440 250152 34440 0 net56
rlabel metal3 193480 4368 193480 4368 0 net57
rlabel metal2 194376 5768 194376 5768 0 net58
rlabel metal3 192136 6664 192136 6664 0 net59
rlabel metal2 141512 4760 141512 4760 0 net6
rlabel metal2 208208 3528 208208 3528 0 net60
rlabel metal2 209160 32368 209160 32368 0 net61
rlabel metal3 280784 55944 280784 55944 0 net62
rlabel metal2 288120 41776 288120 41776 0 net63
rlabel metal3 205520 6440 205520 6440 0 net64
rlabel metal3 188496 55944 188496 55944 0 net65
rlabel metal2 71176 6048 71176 6048 0 net66
rlabel metal2 75096 4480 75096 4480 0 net67
rlabel metal2 78512 3640 78512 3640 0 net68
rlabel metal2 82936 4032 82936 4032 0 net69
rlabel metal2 145096 5152 145096 5152 0 net7
rlabel metal2 45864 38472 45864 38472 0 net70
rlabel metal3 52360 55944 52360 55944 0 net71
rlabel metal2 93576 5544 93576 5544 0 net72
rlabel metal3 93968 4536 93968 4536 0 net73
rlabel metal3 187264 55160 187264 55160 0 net74
rlabel metal2 186200 52528 186200 52528 0 net75
rlabel metal2 168952 54936 168952 54936 0 net76
rlabel metal3 173544 54712 173544 54712 0 net77
rlabel metal2 180264 55412 180264 55412 0 net78
rlabel metal2 184072 55384 184072 55384 0 net79
rlabel metal2 148680 4928 148680 4928 0 net8
rlabel metal2 190456 55412 190456 55412 0 net80
rlabel metal3 194936 56168 194936 56168 0 net81
rlabel metal2 191128 53536 191128 53536 0 net82
rlabel metal3 182392 52808 182392 52808 0 net83
rlabel metal3 131040 54376 131040 54376 0 net84
rlabel metal3 136248 56168 136248 56168 0 net85
rlabel metal3 141960 55384 141960 55384 0 net86
rlabel metal3 146720 54376 146720 54376 0 net87
rlabel metal3 152376 54376 152376 54376 0 net88
rlabel metal2 157416 54936 157416 54936 0 net89
rlabel metal2 186312 3416 186312 3416 0 net9
rlabel metal2 163240 54936 163240 54936 0 net90
rlabel metal2 12208 4536 12208 4536 0 net91
rlabel metal2 43848 14056 43848 14056 0 net92
rlabel metal2 46872 3584 46872 3584 0 net93
rlabel metal2 50792 3864 50792 3864 0 net94
rlabel metal2 54152 4032 54152 4032 0 net95
rlabel metal2 57792 3640 57792 3640 0 net96
rlabel metal2 61488 3640 61488 3640 0 net97
rlabel metal2 68264 19936 68264 19936 0 net98
rlabel metal3 69272 3528 69272 3528 0 net99
rlabel metal2 109592 57778 109592 57778 0 ram_enabled
rlabel metal2 115528 56448 115528 56448 0 requested_addr[0]
rlabel metal2 168784 56280 168784 56280 0 requested_addr[10]
rlabel metal2 174104 57778 174104 57778 0 requested_addr[11]
rlabel metal2 179480 57778 179480 57778 0 requested_addr[12]
rlabel metal2 184856 57778 184856 57778 0 requested_addr[13]
rlabel metal2 191464 56336 191464 56336 0 requested_addr[14]
rlabel metal2 195552 56280 195552 56280 0 requested_addr[15]
rlabel metal2 120344 57778 120344 57778 0 requested_addr[1]
rlabel metal2 125720 57778 125720 57778 0 requested_addr[2]
rlabel metal2 130760 56672 130760 56672 0 requested_addr[3]
rlabel metal2 136472 57778 136472 57778 0 requested_addr[4]
rlabel metal2 142184 56728 142184 56728 0 requested_addr[5]
rlabel metal2 147224 57778 147224 57778 0 requested_addr[6]
rlabel metal2 152600 57778 152600 57778 0 requested_addr[7]
rlabel metal2 157416 56672 157416 56672 0 requested_addr[8]
rlabel metal2 163352 57778 163352 57778 0 requested_addr[9]
rlabel metal2 12768 56280 12768 56280 0 rst
rlabel metal2 162232 53704 162232 53704 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 300000 60000
<< end >>
