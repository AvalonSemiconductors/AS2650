magic
tech gf180mcuD
magscale 1 10
timestamp 1700229967
<< metal1 >>
rect 8530 41694 8542 41746
rect 8594 41743 8606 41746
rect 9426 41743 9438 41746
rect 8594 41697 9438 41743
rect 8594 41694 8606 41697
rect 9426 41694 9438 41697
rect 9490 41694 9502 41746
rect 1344 41578 43568 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 43568 41578
rect 1344 41492 43568 41526
rect 22430 41410 22482 41422
rect 22430 41346 22482 41358
rect 25566 41410 25618 41422
rect 25566 41346 25618 41358
rect 29374 41410 29426 41422
rect 29374 41346 29426 41358
rect 33182 41410 33234 41422
rect 33182 41346 33234 41358
rect 36990 41410 37042 41422
rect 36990 41346 37042 41358
rect 40798 41410 40850 41422
rect 40798 41346 40850 41358
rect 1934 41298 1986 41310
rect 1934 41234 1986 41246
rect 5630 41298 5682 41310
rect 5630 41234 5682 41246
rect 9438 41298 9490 41310
rect 9438 41234 9490 41246
rect 11230 41298 11282 41310
rect 11230 41234 11282 41246
rect 15038 41298 15090 41310
rect 15038 41234 15090 41246
rect 17278 41298 17330 41310
rect 17278 41234 17330 41246
rect 18398 41298 18450 41310
rect 18398 41234 18450 41246
rect 19518 41298 19570 41310
rect 19518 41234 19570 41246
rect 12126 41186 12178 41198
rect 4274 41134 4286 41186
rect 4338 41134 4350 41186
rect 4722 41134 4734 41186
rect 4786 41134 4798 41186
rect 7858 41134 7870 41186
rect 7922 41134 7934 41186
rect 8530 41134 8542 41186
rect 8594 41134 8606 41186
rect 11666 41134 11678 41186
rect 11730 41134 11742 41186
rect 12126 41122 12178 41134
rect 13134 41186 13186 41198
rect 15262 41186 15314 41198
rect 14354 41134 14366 41186
rect 14418 41134 14430 41186
rect 16146 41134 16158 41186
rect 16210 41134 16222 41186
rect 17714 41134 17726 41186
rect 17778 41134 17790 41186
rect 18834 41134 18846 41186
rect 18898 41134 18910 41186
rect 19954 41134 19966 41186
rect 20018 41134 20030 41186
rect 20962 41134 20974 41186
rect 21026 41134 21038 41186
rect 21410 41134 21422 41186
rect 21474 41134 21486 41186
rect 24546 41134 24558 41186
rect 24610 41134 24622 41186
rect 28354 41134 28366 41186
rect 28418 41134 28430 41186
rect 32162 41134 32174 41186
rect 32226 41134 32238 41186
rect 35970 41134 35982 41186
rect 36034 41134 36046 41186
rect 39778 41134 39790 41186
rect 39842 41134 39854 41186
rect 13134 41122 13186 41134
rect 15262 41122 15314 41134
rect 11454 41074 11506 41086
rect 11454 41010 11506 41022
rect 43150 41074 43202 41086
rect 43150 41010 43202 41022
rect 4958 40962 5010 40974
rect 4958 40898 5010 40910
rect 7646 40962 7698 40974
rect 7646 40898 7698 40910
rect 8766 40962 8818 40974
rect 13470 40962 13522 40974
rect 12450 40910 12462 40962
rect 12514 40910 12526 40962
rect 8766 40898 8818 40910
rect 13470 40898 13522 40910
rect 14142 40962 14194 40974
rect 14142 40898 14194 40910
rect 15598 40962 15650 40974
rect 15598 40898 15650 40910
rect 16382 40962 16434 40974
rect 16382 40898 16434 40910
rect 17502 40962 17554 40974
rect 17502 40898 17554 40910
rect 18622 40962 18674 40974
rect 18622 40898 18674 40910
rect 19742 40962 19794 40974
rect 19742 40898 19794 40910
rect 20750 40962 20802 40974
rect 20750 40898 20802 40910
rect 42814 40962 42866 40974
rect 42814 40898 42866 40910
rect 1344 40794 43568 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 43568 40794
rect 1344 40708 43568 40742
rect 9662 40626 9714 40638
rect 9662 40562 9714 40574
rect 13134 40626 13186 40638
rect 13134 40562 13186 40574
rect 13918 40626 13970 40638
rect 13918 40562 13970 40574
rect 16606 40626 16658 40638
rect 16606 40562 16658 40574
rect 21310 40626 21362 40638
rect 21310 40562 21362 40574
rect 26350 40626 26402 40638
rect 26350 40562 26402 40574
rect 29262 40626 29314 40638
rect 29262 40562 29314 40574
rect 34078 40626 34130 40638
rect 34078 40562 34130 40574
rect 36990 40626 37042 40638
rect 36990 40562 37042 40574
rect 7534 40514 7586 40526
rect 5394 40462 5406 40514
rect 5458 40462 5470 40514
rect 7534 40450 7586 40462
rect 7870 40514 7922 40526
rect 7870 40450 7922 40462
rect 8430 40514 8482 40526
rect 8430 40450 8482 40462
rect 8766 40514 8818 40526
rect 8766 40450 8818 40462
rect 11678 40514 11730 40526
rect 11678 40450 11730 40462
rect 12686 40514 12738 40526
rect 12686 40450 12738 40462
rect 24670 40514 24722 40526
rect 24670 40450 24722 40462
rect 31502 40514 31554 40526
rect 31502 40450 31554 40462
rect 11454 40402 11506 40414
rect 12350 40402 12402 40414
rect 31166 40402 31218 40414
rect 43150 40402 43202 40414
rect 4274 40350 4286 40402
rect 4338 40350 4350 40402
rect 7186 40350 7198 40402
rect 7250 40350 7262 40402
rect 11890 40350 11902 40402
rect 11954 40350 11966 40402
rect 24434 40350 24446 40402
rect 24498 40350 24510 40402
rect 25330 40350 25342 40402
rect 25394 40350 25406 40402
rect 28242 40350 28254 40402
rect 28306 40350 28318 40402
rect 33058 40350 33070 40402
rect 33122 40350 33134 40402
rect 35970 40350 35982 40402
rect 36034 40350 36046 40402
rect 11454 40338 11506 40350
rect 12350 40338 12402 40350
rect 31166 40338 31218 40350
rect 43150 40338 43202 40350
rect 15374 40290 15426 40302
rect 15374 40226 15426 40238
rect 1934 40178 1986 40190
rect 1934 40114 1986 40126
rect 1344 40010 43568 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 43568 40010
rect 1344 39924 43568 39958
rect 24110 39842 24162 39854
rect 6850 39790 6862 39842
rect 6914 39839 6926 39842
rect 7522 39839 7534 39842
rect 6914 39793 7534 39839
rect 6914 39790 6926 39793
rect 7522 39790 7534 39793
rect 7586 39790 7598 39842
rect 24110 39778 24162 39790
rect 29374 39842 29426 39854
rect 29374 39778 29426 39790
rect 33070 39842 33122 39854
rect 33070 39778 33122 39790
rect 37998 39842 38050 39854
rect 37998 39778 38050 39790
rect 40910 39842 40962 39854
rect 40910 39778 40962 39790
rect 6862 39730 6914 39742
rect 4610 39678 4622 39730
rect 4674 39678 4686 39730
rect 6862 39666 6914 39678
rect 7198 39730 7250 39742
rect 26238 39730 26290 39742
rect 11554 39678 11566 39730
rect 11618 39678 11630 39730
rect 13458 39678 13470 39730
rect 13522 39678 13534 39730
rect 20626 39678 20638 39730
rect 20690 39678 20702 39730
rect 7198 39666 7250 39678
rect 26238 39666 26290 39678
rect 26014 39618 26066 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 8642 39566 8654 39618
rect 8706 39566 8718 39618
rect 16258 39566 16270 39618
rect 16322 39566 16334 39618
rect 17714 39566 17726 39618
rect 17778 39566 17790 39618
rect 23090 39566 23102 39618
rect 23154 39566 23166 39618
rect 27234 39566 27246 39618
rect 27298 39566 27310 39618
rect 31266 39566 31278 39618
rect 31330 39566 31342 39618
rect 32050 39566 32062 39618
rect 32114 39566 32126 39618
rect 36978 39566 36990 39618
rect 37042 39566 37054 39618
rect 39890 39566 39902 39618
rect 39954 39566 39966 39618
rect 26014 39554 26066 39566
rect 8318 39506 8370 39518
rect 21310 39506 21362 39518
rect 2482 39454 2494 39506
rect 2546 39454 2558 39506
rect 9426 39454 9438 39506
rect 9490 39454 9502 39506
rect 15586 39454 15598 39506
rect 15650 39454 15662 39506
rect 18498 39454 18510 39506
rect 18562 39454 18574 39506
rect 8318 39442 8370 39454
rect 21310 39442 21362 39454
rect 21646 39506 21698 39518
rect 21646 39442 21698 39454
rect 22430 39506 22482 39518
rect 22430 39442 22482 39454
rect 22766 39506 22818 39518
rect 22766 39442 22818 39454
rect 27470 39506 27522 39518
rect 27470 39442 27522 39454
rect 27806 39506 27858 39518
rect 27806 39442 27858 39454
rect 28142 39506 28194 39518
rect 28142 39442 28194 39454
rect 34974 39506 35026 39518
rect 34974 39442 35026 39454
rect 35310 39506 35362 39518
rect 35310 39442 35362 39454
rect 35982 39506 36034 39518
rect 35982 39442 36034 39454
rect 36318 39506 36370 39518
rect 36318 39442 36370 39454
rect 5070 39394 5122 39406
rect 5070 39330 5122 39342
rect 5742 39394 5794 39406
rect 5742 39330 5794 39342
rect 7646 39394 7698 39406
rect 7646 39330 7698 39342
rect 7982 39394 8034 39406
rect 7982 39330 8034 39342
rect 12014 39394 12066 39406
rect 12014 39330 12066 39342
rect 12910 39394 12962 39406
rect 12910 39330 12962 39342
rect 17390 39394 17442 39406
rect 28702 39394 28754 39406
rect 26562 39342 26574 39394
rect 26626 39342 26638 39394
rect 17390 39330 17442 39342
rect 28702 39330 28754 39342
rect 1344 39226 43568 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 43568 39226
rect 1344 39140 43568 39174
rect 8318 39058 8370 39070
rect 8318 38994 8370 39006
rect 9662 39058 9714 39070
rect 9662 38994 9714 39006
rect 15710 39058 15762 39070
rect 18286 39058 18338 39070
rect 16818 39006 16830 39058
rect 16882 39006 16894 39058
rect 15710 38994 15762 39006
rect 18286 38994 18338 39006
rect 20414 39058 20466 39070
rect 20414 38994 20466 39006
rect 23886 39058 23938 39070
rect 26686 39058 26738 39070
rect 24658 39006 24670 39058
rect 24722 39006 24734 39058
rect 25778 39006 25790 39058
rect 25842 39006 25854 39058
rect 23886 38994 23938 39006
rect 26686 38994 26738 39006
rect 27918 39058 27970 39070
rect 27918 38994 27970 39006
rect 30830 39058 30882 39070
rect 30830 38994 30882 39006
rect 31502 39058 31554 39070
rect 31502 38994 31554 39006
rect 32174 39058 32226 39070
rect 32174 38994 32226 39006
rect 33406 39058 33458 39070
rect 33406 38994 33458 39006
rect 36430 39058 36482 39070
rect 36430 38994 36482 39006
rect 19630 38946 19682 38958
rect 38334 38946 38386 38958
rect 29138 38894 29150 38946
rect 29202 38894 29214 38946
rect 19630 38882 19682 38894
rect 38334 38882 38386 38894
rect 38670 38946 38722 38958
rect 38670 38882 38722 38894
rect 39118 38946 39170 38958
rect 39118 38882 39170 38894
rect 39454 38946 39506 38958
rect 39454 38882 39506 38894
rect 9438 38834 9490 38846
rect 1922 38782 1934 38834
rect 1986 38782 1998 38834
rect 5170 38782 5182 38834
rect 5234 38782 5246 38834
rect 9438 38770 9490 38782
rect 9886 38834 9938 38846
rect 9886 38770 9938 38782
rect 10110 38834 10162 38846
rect 15486 38834 15538 38846
rect 14914 38782 14926 38834
rect 14978 38782 14990 38834
rect 10110 38770 10162 38782
rect 15486 38770 15538 38782
rect 15598 38834 15650 38846
rect 15598 38770 15650 38782
rect 16046 38834 16098 38846
rect 16046 38770 16098 38782
rect 16494 38834 16546 38846
rect 16494 38770 16546 38782
rect 18062 38834 18114 38846
rect 18062 38770 18114 38782
rect 18286 38834 18338 38846
rect 18286 38770 18338 38782
rect 18622 38834 18674 38846
rect 24334 38834 24386 38846
rect 20178 38782 20190 38834
rect 20242 38782 20254 38834
rect 18622 38770 18674 38782
rect 24334 38770 24386 38782
rect 25230 38834 25282 38846
rect 25230 38770 25282 38782
rect 27582 38834 27634 38846
rect 29710 38834 29762 38846
rect 28914 38782 28926 38834
rect 28978 38782 28990 38834
rect 27582 38770 27634 38782
rect 29710 38770 29762 38782
rect 30046 38834 30098 38846
rect 31166 38834 31218 38846
rect 33070 38834 33122 38846
rect 30594 38782 30606 38834
rect 30658 38782 30670 38834
rect 31938 38782 31950 38834
rect 32002 38782 32014 38834
rect 35634 38782 35646 38834
rect 35698 38782 35710 38834
rect 30046 38770 30098 38782
rect 31166 38770 31218 38782
rect 33070 38770 33122 38782
rect 16270 38722 16322 38734
rect 2594 38670 2606 38722
rect 2658 38670 2670 38722
rect 4722 38670 4734 38722
rect 4786 38670 4798 38722
rect 5842 38670 5854 38722
rect 5906 38670 5918 38722
rect 7970 38670 7982 38722
rect 8034 38670 8046 38722
rect 8754 38670 8766 38722
rect 8818 38670 8830 38722
rect 12114 38670 12126 38722
rect 12178 38670 12190 38722
rect 14242 38670 14254 38722
rect 14306 38670 14318 38722
rect 16270 38658 16322 38670
rect 17614 38722 17666 38734
rect 17614 38658 17666 38670
rect 19518 38722 19570 38734
rect 19518 38658 19570 38670
rect 24110 38722 24162 38734
rect 24110 38658 24162 38670
rect 26238 38722 26290 38734
rect 26238 38658 26290 38670
rect 28366 38722 28418 38734
rect 28366 38658 28418 38670
rect 25454 38610 25506 38622
rect 25454 38546 25506 38558
rect 1344 38442 43568 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 43568 38442
rect 1344 38356 43568 38390
rect 13918 38274 13970 38286
rect 40910 38274 40962 38286
rect 15810 38222 15822 38274
rect 15874 38222 15886 38274
rect 13918 38210 13970 38222
rect 40910 38210 40962 38222
rect 1934 38162 1986 38174
rect 11790 38162 11842 38174
rect 8418 38110 8430 38162
rect 8482 38110 8494 38162
rect 1934 38098 1986 38110
rect 11790 38098 11842 38110
rect 14478 38162 14530 38174
rect 14478 38098 14530 38110
rect 16942 38162 16994 38174
rect 20738 38110 20750 38162
rect 20802 38110 20814 38162
rect 25778 38110 25790 38162
rect 25842 38110 25854 38162
rect 16942 38098 16994 38110
rect 5742 38050 5794 38062
rect 14030 38050 14082 38062
rect 4274 37998 4286 38050
rect 4338 37998 4350 38050
rect 4834 37998 4846 38050
rect 4898 37998 4910 38050
rect 11330 37998 11342 38050
rect 11394 37998 11406 38050
rect 5742 37986 5794 37998
rect 14030 37986 14082 37998
rect 14254 38050 14306 38062
rect 14254 37986 14306 37998
rect 14814 38050 14866 38062
rect 14814 37986 14866 37998
rect 15262 38050 15314 38062
rect 15262 37986 15314 37998
rect 15486 38050 15538 38062
rect 15486 37986 15538 37998
rect 16046 38050 16098 38062
rect 16046 37986 16098 37998
rect 16382 38050 16434 38062
rect 16382 37986 16434 37998
rect 17278 38050 17330 38062
rect 17826 37998 17838 38050
rect 17890 37998 17902 38050
rect 22978 37998 22990 38050
rect 23042 37998 23054 38050
rect 29250 37998 29262 38050
rect 29314 37998 29326 38050
rect 39890 37998 39902 38050
rect 39954 37998 39966 38050
rect 17278 37986 17330 37998
rect 8094 37938 8146 37950
rect 14702 37938 14754 37950
rect 10546 37886 10558 37938
rect 10610 37886 10622 37938
rect 8094 37874 8146 37886
rect 14702 37874 14754 37886
rect 16270 37938 16322 37950
rect 16270 37874 16322 37886
rect 17614 37938 17666 37950
rect 28702 37938 28754 37950
rect 18610 37886 18622 37938
rect 18674 37886 18686 37938
rect 23650 37886 23662 37938
rect 23714 37886 23726 37938
rect 17614 37874 17666 37886
rect 28702 37874 28754 37886
rect 29486 37938 29538 37950
rect 29486 37874 29538 37886
rect 5070 37826 5122 37838
rect 5070 37762 5122 37774
rect 7534 37826 7586 37838
rect 7534 37762 7586 37774
rect 7758 37826 7810 37838
rect 7758 37762 7810 37774
rect 12910 37826 12962 37838
rect 12910 37762 12962 37774
rect 13918 37826 13970 37838
rect 13918 37762 13970 37774
rect 17390 37826 17442 37838
rect 17390 37762 17442 37774
rect 26238 37826 26290 37838
rect 26238 37762 26290 37774
rect 31502 37826 31554 37838
rect 31502 37762 31554 37774
rect 1344 37658 43568 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 43568 37658
rect 1344 37572 43568 37606
rect 7534 37490 7586 37502
rect 7534 37426 7586 37438
rect 9774 37490 9826 37502
rect 9774 37426 9826 37438
rect 15262 37490 15314 37502
rect 15262 37426 15314 37438
rect 15486 37490 15538 37502
rect 15486 37426 15538 37438
rect 15934 37490 15986 37502
rect 15934 37426 15986 37438
rect 16270 37490 16322 37502
rect 16270 37426 16322 37438
rect 17502 37490 17554 37502
rect 17502 37426 17554 37438
rect 18286 37490 18338 37502
rect 18286 37426 18338 37438
rect 18622 37490 18674 37502
rect 18622 37426 18674 37438
rect 6750 37378 6802 37390
rect 6750 37314 6802 37326
rect 8430 37378 8482 37390
rect 8430 37314 8482 37326
rect 8654 37378 8706 37390
rect 8654 37314 8706 37326
rect 10110 37378 10162 37390
rect 10110 37314 10162 37326
rect 10558 37378 10610 37390
rect 17390 37378 17442 37390
rect 12562 37326 12574 37378
rect 12626 37326 12638 37378
rect 14578 37326 14590 37378
rect 14642 37326 14654 37378
rect 10558 37314 10610 37326
rect 17390 37314 17442 37326
rect 18062 37378 18114 37390
rect 18062 37314 18114 37326
rect 19518 37378 19570 37390
rect 19518 37314 19570 37326
rect 7422 37266 7474 37278
rect 4274 37214 4286 37266
rect 4338 37214 4350 37266
rect 6962 37214 6974 37266
rect 7026 37214 7038 37266
rect 7422 37202 7474 37214
rect 7758 37266 7810 37278
rect 7758 37202 7810 37214
rect 7982 37266 8034 37278
rect 7982 37202 8034 37214
rect 8318 37266 8370 37278
rect 8318 37202 8370 37214
rect 9438 37266 9490 37278
rect 9438 37202 9490 37214
rect 9774 37266 9826 37278
rect 9774 37202 9826 37214
rect 10446 37266 10498 37278
rect 10446 37202 10498 37214
rect 12350 37266 12402 37278
rect 15150 37266 15202 37278
rect 13346 37214 13358 37266
rect 13410 37214 13422 37266
rect 13906 37214 13918 37266
rect 13970 37214 13982 37266
rect 14354 37214 14366 37266
rect 14418 37214 14430 37266
rect 12350 37202 12402 37214
rect 15150 37202 15202 37214
rect 17726 37266 17778 37278
rect 17726 37202 17778 37214
rect 17950 37266 18002 37278
rect 17950 37202 18002 37214
rect 18398 37266 18450 37278
rect 18398 37202 18450 37214
rect 18734 37266 18786 37278
rect 18734 37202 18786 37214
rect 19070 37266 19122 37278
rect 19070 37202 19122 37214
rect 6526 37154 6578 37166
rect 6526 37090 6578 37102
rect 8990 37154 9042 37166
rect 8990 37090 9042 37102
rect 11118 37154 11170 37166
rect 13010 37102 13022 37154
rect 13074 37102 13086 37154
rect 11118 37090 11170 37102
rect 1934 37042 1986 37054
rect 1934 36978 1986 36990
rect 10558 37042 10610 37054
rect 10558 36978 10610 36990
rect 1344 36874 43568 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 43568 36874
rect 1344 36788 43568 36822
rect 15374 36706 15426 36718
rect 15374 36642 15426 36654
rect 18286 36706 18338 36718
rect 18286 36642 18338 36654
rect 41582 36706 41634 36718
rect 41582 36642 41634 36654
rect 5854 36594 5906 36606
rect 2034 36542 2046 36594
rect 2098 36542 2110 36594
rect 5854 36530 5906 36542
rect 14926 36594 14978 36606
rect 14926 36530 14978 36542
rect 23214 36594 23266 36606
rect 28578 36542 28590 36594
rect 28642 36542 28654 36594
rect 23214 36530 23266 36542
rect 5630 36482 5682 36494
rect 4050 36430 4062 36482
rect 4114 36430 4126 36482
rect 4834 36430 4846 36482
rect 4898 36430 4910 36482
rect 5630 36418 5682 36430
rect 5966 36482 6018 36494
rect 5966 36418 6018 36430
rect 6526 36482 6578 36494
rect 6526 36418 6578 36430
rect 7310 36482 7362 36494
rect 7310 36418 7362 36430
rect 7646 36482 7698 36494
rect 7646 36418 7698 36430
rect 7758 36482 7810 36494
rect 7758 36418 7810 36430
rect 8094 36482 8146 36494
rect 8094 36418 8146 36430
rect 8430 36482 8482 36494
rect 8430 36418 8482 36430
rect 9438 36482 9490 36494
rect 9438 36418 9490 36430
rect 9774 36482 9826 36494
rect 9774 36418 9826 36430
rect 15486 36482 15538 36494
rect 15486 36418 15538 36430
rect 16830 36482 16882 36494
rect 23326 36482 23378 36494
rect 20514 36430 20526 36482
rect 20578 36430 20590 36482
rect 16830 36418 16882 36430
rect 23326 36418 23378 36430
rect 23662 36482 23714 36494
rect 23662 36418 23714 36430
rect 23886 36482 23938 36494
rect 23886 36418 23938 36430
rect 24446 36482 24498 36494
rect 25666 36430 25678 36482
rect 25730 36430 25742 36482
rect 40562 36430 40574 36482
rect 40626 36430 40638 36482
rect 24446 36418 24498 36430
rect 6302 36370 6354 36382
rect 5058 36318 5070 36370
rect 5122 36318 5134 36370
rect 6302 36306 6354 36318
rect 6750 36370 6802 36382
rect 6750 36306 6802 36318
rect 6862 36370 6914 36382
rect 6862 36306 6914 36318
rect 8766 36370 8818 36382
rect 8766 36306 8818 36318
rect 16494 36370 16546 36382
rect 16494 36306 16546 36318
rect 18174 36370 18226 36382
rect 22542 36370 22594 36382
rect 20290 36318 20302 36370
rect 20354 36318 20366 36370
rect 18174 36306 18226 36318
rect 22542 36306 22594 36318
rect 22654 36370 22706 36382
rect 22654 36306 22706 36318
rect 22878 36370 22930 36382
rect 22878 36306 22930 36318
rect 23102 36370 23154 36382
rect 23102 36306 23154 36318
rect 24334 36370 24386 36382
rect 26450 36318 26462 36370
rect 26514 36318 26526 36370
rect 24334 36306 24386 36318
rect 7422 36258 7474 36270
rect 7422 36194 7474 36206
rect 7982 36258 8034 36270
rect 7982 36194 8034 36206
rect 9550 36258 9602 36270
rect 9550 36194 9602 36206
rect 10222 36258 10274 36270
rect 10222 36194 10274 36206
rect 15374 36258 15426 36270
rect 15374 36194 15426 36206
rect 16046 36258 16098 36270
rect 16046 36194 16098 36206
rect 18286 36258 18338 36270
rect 18286 36194 18338 36206
rect 18958 36258 19010 36270
rect 18958 36194 19010 36206
rect 24222 36258 24274 36270
rect 24222 36194 24274 36206
rect 25006 36258 25058 36270
rect 25006 36194 25058 36206
rect 1344 36090 43568 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 43568 36090
rect 1344 36004 43568 36038
rect 5070 35922 5122 35934
rect 5070 35858 5122 35870
rect 5294 35922 5346 35934
rect 5294 35858 5346 35870
rect 6750 35922 6802 35934
rect 6750 35858 6802 35870
rect 7086 35922 7138 35934
rect 7086 35858 7138 35870
rect 7422 35922 7474 35934
rect 7422 35858 7474 35870
rect 12350 35922 12402 35934
rect 21198 35922 21250 35934
rect 22542 35922 22594 35934
rect 17714 35870 17726 35922
rect 17778 35870 17790 35922
rect 21522 35870 21534 35922
rect 21586 35870 21598 35922
rect 12350 35858 12402 35870
rect 21198 35858 21250 35870
rect 22542 35858 22594 35870
rect 23326 35922 23378 35934
rect 23326 35858 23378 35870
rect 4958 35810 5010 35822
rect 4958 35746 5010 35758
rect 7198 35810 7250 35822
rect 7198 35746 7250 35758
rect 7646 35810 7698 35822
rect 7646 35746 7698 35758
rect 7758 35810 7810 35822
rect 21982 35810 22034 35822
rect 12786 35758 12798 35810
rect 12850 35758 12862 35810
rect 14578 35758 14590 35810
rect 14642 35758 14654 35810
rect 7758 35746 7810 35758
rect 21982 35746 22034 35758
rect 22990 35810 23042 35822
rect 22990 35746 23042 35758
rect 23102 35810 23154 35822
rect 23102 35746 23154 35758
rect 23662 35810 23714 35822
rect 23662 35746 23714 35758
rect 25230 35810 25282 35822
rect 25230 35746 25282 35758
rect 8990 35698 9042 35710
rect 1810 35646 1822 35698
rect 1874 35646 1886 35698
rect 8990 35634 9042 35646
rect 11902 35698 11954 35710
rect 15262 35698 15314 35710
rect 21870 35698 21922 35710
rect 13346 35646 13358 35698
rect 13410 35646 13422 35698
rect 13906 35646 13918 35698
rect 13970 35646 13982 35698
rect 14354 35646 14366 35698
rect 14418 35646 14430 35698
rect 17938 35646 17950 35698
rect 18002 35646 18014 35698
rect 11902 35634 11954 35646
rect 15262 35634 15314 35646
rect 21870 35634 21922 35646
rect 22430 35698 22482 35710
rect 22430 35634 22482 35646
rect 22766 35698 22818 35710
rect 22766 35634 22818 35646
rect 23550 35698 23602 35710
rect 23550 35634 23602 35646
rect 23998 35698 24050 35710
rect 23998 35634 24050 35646
rect 24334 35698 24386 35710
rect 24334 35634 24386 35646
rect 24558 35698 24610 35710
rect 24558 35634 24610 35646
rect 25454 35698 25506 35710
rect 25454 35634 25506 35646
rect 25790 35698 25842 35710
rect 28802 35646 28814 35698
rect 28866 35646 28878 35698
rect 25790 35634 25842 35646
rect 5630 35586 5682 35598
rect 2482 35534 2494 35586
rect 2546 35534 2558 35586
rect 4610 35534 4622 35586
rect 4674 35534 4686 35586
rect 5630 35522 5682 35534
rect 8542 35586 8594 35598
rect 8542 35522 8594 35534
rect 10894 35586 10946 35598
rect 16270 35586 16322 35598
rect 13010 35534 13022 35586
rect 13074 35534 13086 35586
rect 10894 35522 10946 35534
rect 16270 35522 16322 35534
rect 20862 35586 20914 35598
rect 20862 35522 20914 35534
rect 24222 35586 24274 35598
rect 24222 35522 24274 35534
rect 25678 35586 25730 35598
rect 29586 35534 29598 35586
rect 29650 35534 29662 35586
rect 31714 35534 31726 35586
rect 31778 35534 31790 35586
rect 25678 35522 25730 35534
rect 7086 35474 7138 35486
rect 7086 35410 7138 35422
rect 21982 35474 22034 35486
rect 21982 35410 22034 35422
rect 23662 35474 23714 35486
rect 23662 35410 23714 35422
rect 1344 35306 43568 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 43568 35306
rect 1344 35220 43568 35254
rect 15822 35138 15874 35150
rect 15822 35074 15874 35086
rect 1934 35026 1986 35038
rect 1934 34962 1986 34974
rect 4734 35026 4786 35038
rect 4734 34962 4786 34974
rect 11006 35026 11058 35038
rect 11006 34962 11058 34974
rect 11342 35026 11394 35038
rect 11342 34962 11394 34974
rect 13582 35026 13634 35038
rect 13582 34962 13634 34974
rect 21982 35026 22034 35038
rect 21982 34962 22034 34974
rect 22990 35026 23042 35038
rect 22990 34962 23042 34974
rect 23438 35026 23490 35038
rect 26338 34974 26350 35026
rect 26402 34974 26414 35026
rect 28466 34974 28478 35026
rect 28530 34974 28542 35026
rect 23438 34962 23490 34974
rect 5518 34914 5570 34926
rect 4274 34862 4286 34914
rect 4338 34862 4350 34914
rect 5518 34850 5570 34862
rect 5966 34914 6018 34926
rect 5966 34850 6018 34862
rect 6190 34914 6242 34926
rect 6190 34850 6242 34862
rect 7422 34914 7474 34926
rect 7422 34850 7474 34862
rect 10558 34914 10610 34926
rect 10558 34850 10610 34862
rect 11566 34914 11618 34926
rect 15374 34914 15426 34926
rect 11778 34862 11790 34914
rect 11842 34862 11854 34914
rect 14914 34862 14926 34914
rect 14978 34862 14990 34914
rect 11566 34850 11618 34862
rect 15374 34850 15426 34862
rect 16942 34914 16994 34926
rect 16942 34850 16994 34862
rect 22654 34914 22706 34926
rect 22654 34850 22706 34862
rect 23774 34914 23826 34926
rect 23774 34850 23826 34862
rect 24110 34914 24162 34926
rect 24546 34862 24558 34914
rect 24610 34862 24622 34914
rect 25554 34862 25566 34914
rect 25618 34862 25630 34914
rect 24110 34850 24162 34862
rect 6862 34802 6914 34814
rect 6862 34738 6914 34750
rect 7086 34802 7138 34814
rect 14590 34802 14642 34814
rect 10210 34750 10222 34802
rect 10274 34750 10286 34802
rect 7086 34738 7138 34750
rect 14590 34738 14642 34750
rect 15710 34802 15762 34814
rect 15710 34738 15762 34750
rect 20190 34802 20242 34814
rect 22318 34802 22370 34814
rect 20514 34750 20526 34802
rect 20578 34750 20590 34802
rect 20190 34738 20242 34750
rect 22318 34738 22370 34750
rect 22430 34802 22482 34814
rect 22430 34738 22482 34750
rect 24334 34802 24386 34814
rect 24334 34738 24386 34750
rect 4622 34690 4674 34702
rect 4622 34626 4674 34638
rect 5742 34690 5794 34702
rect 5742 34626 5794 34638
rect 7310 34690 7362 34702
rect 7310 34626 7362 34638
rect 11454 34690 11506 34702
rect 11454 34626 11506 34638
rect 12014 34690 12066 34702
rect 12014 34626 12066 34638
rect 12126 34690 12178 34702
rect 12126 34626 12178 34638
rect 12798 34690 12850 34702
rect 12798 34626 12850 34638
rect 15822 34690 15874 34702
rect 15822 34626 15874 34638
rect 16494 34690 16546 34702
rect 16494 34626 16546 34638
rect 17390 34690 17442 34702
rect 17390 34626 17442 34638
rect 17726 34690 17778 34702
rect 17726 34626 17778 34638
rect 23886 34690 23938 34702
rect 23886 34626 23938 34638
rect 1344 34522 43568 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 43568 34522
rect 1344 34436 43568 34470
rect 18734 34354 18786 34366
rect 2818 34302 2830 34354
rect 2882 34302 2894 34354
rect 17938 34302 17950 34354
rect 18002 34302 18014 34354
rect 18734 34290 18786 34302
rect 20638 34354 20690 34366
rect 20638 34290 20690 34302
rect 24110 34354 24162 34366
rect 24110 34290 24162 34302
rect 26910 34354 26962 34366
rect 26910 34290 26962 34302
rect 28254 34354 28306 34366
rect 28254 34290 28306 34302
rect 29934 34354 29986 34366
rect 29934 34290 29986 34302
rect 30830 34354 30882 34366
rect 30830 34290 30882 34302
rect 32510 34354 32562 34366
rect 32510 34290 32562 34302
rect 2046 34242 2098 34254
rect 23774 34242 23826 34254
rect 2706 34190 2718 34242
rect 2770 34190 2782 34242
rect 5730 34190 5742 34242
rect 5794 34190 5806 34242
rect 7634 34190 7646 34242
rect 7698 34190 7710 34242
rect 19618 34190 19630 34242
rect 19682 34190 19694 34242
rect 2046 34178 2098 34190
rect 23774 34178 23826 34190
rect 23886 34242 23938 34254
rect 28914 34190 28926 34242
rect 28978 34190 28990 34242
rect 29138 34190 29150 34242
rect 29202 34190 29214 34242
rect 31714 34190 31726 34242
rect 31778 34190 31790 34242
rect 23886 34178 23938 34190
rect 2158 34130 2210 34142
rect 2158 34066 2210 34078
rect 2494 34130 2546 34142
rect 6974 34130 7026 34142
rect 3266 34078 3278 34130
rect 3330 34078 3342 34130
rect 6514 34078 6526 34130
rect 6578 34078 6590 34130
rect 2494 34066 2546 34078
rect 6974 34066 7026 34078
rect 7422 34130 7474 34142
rect 17390 34130 17442 34142
rect 12786 34078 12798 34130
rect 12850 34078 12862 34130
rect 7422 34066 7474 34078
rect 17390 34066 17442 34078
rect 17614 34130 17666 34142
rect 20302 34130 20354 34142
rect 19506 34078 19518 34130
rect 19570 34078 19582 34130
rect 31938 34078 31950 34130
rect 32002 34078 32014 34130
rect 17614 34066 17666 34078
rect 20302 34066 20354 34078
rect 7758 34018 7810 34030
rect 3602 33966 3614 34018
rect 3666 33966 3678 34018
rect 7758 33954 7810 33966
rect 8318 34018 8370 34030
rect 8318 33954 8370 33966
rect 10558 34018 10610 34030
rect 19070 34018 19122 34030
rect 13346 33966 13358 34018
rect 13410 33966 13422 34018
rect 10558 33954 10610 33966
rect 19070 33954 19122 33966
rect 24446 34018 24498 34030
rect 24446 33954 24498 33966
rect 30382 34018 30434 34030
rect 30382 33954 30434 33966
rect 33182 34018 33234 34030
rect 33182 33954 33234 33966
rect 6750 33906 6802 33918
rect 3042 33854 3054 33906
rect 3106 33854 3118 33906
rect 6750 33842 6802 33854
rect 28590 33906 28642 33918
rect 28590 33842 28642 33854
rect 31166 33906 31218 33918
rect 31166 33842 31218 33854
rect 1344 33738 43568 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 43568 33738
rect 1344 33652 43568 33686
rect 25566 33570 25618 33582
rect 25566 33506 25618 33518
rect 27358 33570 27410 33582
rect 27358 33506 27410 33518
rect 1934 33458 1986 33470
rect 1934 33394 1986 33406
rect 6750 33458 6802 33470
rect 6750 33394 6802 33406
rect 7310 33458 7362 33470
rect 7310 33394 7362 33406
rect 11902 33458 11954 33470
rect 11902 33394 11954 33406
rect 12350 33458 12402 33470
rect 30158 33458 30210 33470
rect 16930 33406 16942 33458
rect 16994 33406 17006 33458
rect 12350 33394 12402 33406
rect 30158 33394 30210 33406
rect 4622 33346 4674 33358
rect 4274 33294 4286 33346
rect 4338 33294 4350 33346
rect 4622 33282 4674 33294
rect 4958 33346 5010 33358
rect 4958 33282 5010 33294
rect 9774 33346 9826 33358
rect 9774 33282 9826 33294
rect 10894 33346 10946 33358
rect 10894 33282 10946 33294
rect 11230 33346 11282 33358
rect 11230 33282 11282 33294
rect 11566 33346 11618 33358
rect 15710 33346 15762 33358
rect 14690 33294 14702 33346
rect 14754 33294 14766 33346
rect 15250 33294 15262 33346
rect 15314 33294 15326 33346
rect 11566 33282 11618 33294
rect 15710 33282 15762 33294
rect 16494 33346 16546 33358
rect 25230 33346 25282 33358
rect 19730 33294 19742 33346
rect 19794 33294 19806 33346
rect 24434 33294 24446 33346
rect 24498 33294 24510 33346
rect 16494 33282 16546 33294
rect 25230 33282 25282 33294
rect 26574 33346 26626 33358
rect 26574 33282 26626 33294
rect 27694 33346 27746 33358
rect 27694 33282 27746 33294
rect 7758 33234 7810 33246
rect 7758 33170 7810 33182
rect 8094 33234 8146 33246
rect 8094 33170 8146 33182
rect 10222 33234 10274 33246
rect 10222 33170 10274 33182
rect 10782 33234 10834 33246
rect 14242 33182 14254 33234
rect 14306 33182 14318 33234
rect 16258 33182 16270 33234
rect 16322 33182 16334 33234
rect 19058 33182 19070 33234
rect 19122 33182 19134 33234
rect 24658 33182 24670 33234
rect 24722 33182 24734 33234
rect 27906 33182 27918 33234
rect 27970 33182 27982 33234
rect 28466 33182 28478 33234
rect 28530 33182 28542 33234
rect 10782 33170 10834 33182
rect 4734 33122 4786 33134
rect 4734 33058 4786 33070
rect 9662 33122 9714 33134
rect 9662 33058 9714 33070
rect 9886 33122 9938 33134
rect 9886 33058 9938 33070
rect 9998 33122 10050 33134
rect 9998 33058 10050 33070
rect 10670 33122 10722 33134
rect 10670 33058 10722 33070
rect 11342 33122 11394 33134
rect 11342 33058 11394 33070
rect 12910 33122 12962 33134
rect 12910 33058 12962 33070
rect 13806 33122 13858 33134
rect 13806 33058 13858 33070
rect 14030 33122 14082 33134
rect 14030 33058 14082 33070
rect 26126 33122 26178 33134
rect 26126 33058 26178 33070
rect 29262 33122 29314 33134
rect 29262 33058 29314 33070
rect 1344 32954 43568 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 43568 32954
rect 1344 32868 43568 32902
rect 5294 32786 5346 32798
rect 2370 32734 2382 32786
rect 2434 32734 2446 32786
rect 5294 32722 5346 32734
rect 6414 32786 6466 32798
rect 6414 32722 6466 32734
rect 8654 32786 8706 32798
rect 8654 32722 8706 32734
rect 10334 32786 10386 32798
rect 16718 32786 16770 32798
rect 14578 32734 14590 32786
rect 14642 32734 14654 32786
rect 10334 32722 10386 32734
rect 16718 32722 16770 32734
rect 18174 32786 18226 32798
rect 18174 32722 18226 32734
rect 2046 32674 2098 32686
rect 6190 32674 6242 32686
rect 2258 32622 2270 32674
rect 2322 32622 2334 32674
rect 2046 32610 2098 32622
rect 6190 32610 6242 32622
rect 8318 32674 8370 32686
rect 10546 32622 10558 32674
rect 10610 32622 10622 32674
rect 12562 32622 12574 32674
rect 12626 32622 12638 32674
rect 14354 32622 14366 32674
rect 14418 32622 14430 32674
rect 16258 32622 16270 32674
rect 16322 32622 16334 32674
rect 8318 32610 8370 32622
rect 6078 32562 6130 32574
rect 2818 32510 2830 32562
rect 2882 32510 2894 32562
rect 5506 32510 5518 32562
rect 5570 32510 5582 32562
rect 6078 32498 6130 32510
rect 6638 32562 6690 32574
rect 6638 32498 6690 32510
rect 7198 32562 7250 32574
rect 7198 32498 7250 32510
rect 7646 32562 7698 32574
rect 7646 32498 7698 32510
rect 7758 32562 7810 32574
rect 7758 32498 7810 32510
rect 8542 32562 8594 32574
rect 8542 32498 8594 32510
rect 8766 32562 8818 32574
rect 8766 32498 8818 32510
rect 8878 32562 8930 32574
rect 18062 32562 18114 32574
rect 11218 32510 11230 32562
rect 11282 32510 11294 32562
rect 11666 32510 11678 32562
rect 11730 32510 11742 32562
rect 12338 32510 12350 32562
rect 12402 32510 12414 32562
rect 13906 32510 13918 32562
rect 13970 32510 13982 32562
rect 14914 32510 14926 32562
rect 14978 32510 14990 32562
rect 15138 32510 15150 32562
rect 15202 32510 15214 32562
rect 15810 32510 15822 32562
rect 15874 32510 15886 32562
rect 17490 32510 17502 32562
rect 17554 32510 17566 32562
rect 8878 32498 8930 32510
rect 18062 32498 18114 32510
rect 18622 32562 18674 32574
rect 26674 32510 26686 32562
rect 26738 32510 26750 32562
rect 18622 32498 18674 32510
rect 3278 32450 3330 32462
rect 3278 32386 3330 32398
rect 3726 32450 3778 32462
rect 3726 32386 3778 32398
rect 7982 32450 8034 32462
rect 13134 32450 13186 32462
rect 24670 32450 24722 32462
rect 10994 32398 11006 32450
rect 11058 32398 11070 32450
rect 13570 32398 13582 32450
rect 13634 32398 13646 32450
rect 17714 32398 17726 32450
rect 17778 32398 17790 32450
rect 27234 32398 27246 32450
rect 27298 32398 27310 32450
rect 7982 32386 8034 32398
rect 13134 32386 13186 32398
rect 24670 32386 24722 32398
rect 2494 32338 2546 32350
rect 2494 32274 2546 32286
rect 6974 32338 7026 32350
rect 6974 32274 7026 32286
rect 1344 32170 43568 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 43568 32170
rect 1344 32084 43568 32118
rect 13794 31950 13806 32002
rect 13858 31999 13870 32002
rect 14466 31999 14478 32002
rect 13858 31953 14478 31999
rect 13858 31950 13870 31953
rect 14466 31950 14478 31953
rect 14530 31950 14542 32002
rect 1934 31890 1986 31902
rect 1934 31826 1986 31838
rect 7086 31890 7138 31902
rect 7086 31826 7138 31838
rect 8094 31890 8146 31902
rect 8094 31826 8146 31838
rect 9886 31890 9938 31902
rect 24210 31838 24222 31890
rect 24274 31838 24286 31890
rect 32050 31838 32062 31890
rect 32114 31838 32126 31890
rect 9886 31826 9938 31838
rect 6526 31778 6578 31790
rect 4050 31726 4062 31778
rect 4114 31726 4126 31778
rect 5954 31726 5966 31778
rect 6018 31726 6030 31778
rect 6526 31714 6578 31726
rect 7310 31778 7362 31790
rect 7310 31714 7362 31726
rect 7870 31778 7922 31790
rect 15822 31778 15874 31790
rect 24558 31778 24610 31790
rect 9538 31726 9550 31778
rect 9602 31726 9614 31778
rect 10210 31726 10222 31778
rect 10274 31726 10286 31778
rect 15362 31726 15374 31778
rect 15426 31726 15438 31778
rect 21298 31726 21310 31778
rect 21362 31726 21374 31778
rect 7870 31714 7922 31726
rect 15822 31714 15874 31726
rect 24558 31714 24610 31726
rect 24782 31778 24834 31790
rect 25106 31726 25118 31778
rect 25170 31726 25182 31778
rect 29250 31726 29262 31778
rect 29314 31726 29326 31778
rect 24782 31714 24834 31726
rect 8318 31666 8370 31678
rect 7634 31614 7646 31666
rect 7698 31614 7710 31666
rect 8318 31602 8370 31614
rect 9998 31666 10050 31678
rect 11342 31666 11394 31678
rect 10546 31614 10558 31666
rect 10610 31614 10622 31666
rect 9998 31602 10050 31614
rect 11342 31602 11394 31614
rect 17054 31666 17106 31678
rect 42814 31666 42866 31678
rect 22082 31614 22094 31666
rect 22146 31614 22158 31666
rect 29922 31614 29934 31666
rect 29986 31614 29998 31666
rect 37314 31614 37326 31666
rect 37378 31614 37390 31666
rect 17054 31602 17106 31614
rect 42814 31602 42866 31614
rect 43150 31666 43202 31678
rect 43150 31602 43202 31614
rect 8206 31554 8258 31566
rect 6178 31502 6190 31554
rect 6242 31502 6254 31554
rect 8206 31490 8258 31502
rect 9214 31554 9266 31566
rect 9214 31490 9266 31502
rect 9774 31554 9826 31566
rect 9774 31490 9826 31502
rect 10894 31554 10946 31566
rect 10894 31490 10946 31502
rect 14030 31554 14082 31566
rect 14030 31490 14082 31502
rect 14478 31554 14530 31566
rect 14478 31490 14530 31502
rect 14926 31554 14978 31566
rect 14926 31490 14978 31502
rect 16158 31554 16210 31566
rect 36990 31554 37042 31566
rect 16482 31502 16494 31554
rect 16546 31502 16558 31554
rect 16158 31490 16210 31502
rect 36990 31490 37042 31502
rect 42590 31554 42642 31566
rect 42590 31490 42642 31502
rect 1344 31386 43568 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 43568 31386
rect 1344 31300 43568 31334
rect 4062 31218 4114 31230
rect 4062 31154 4114 31166
rect 5406 31218 5458 31230
rect 5406 31154 5458 31166
rect 20302 31218 20354 31230
rect 20302 31154 20354 31166
rect 20974 31218 21026 31230
rect 20974 31154 21026 31166
rect 23662 31218 23714 31230
rect 23662 31154 23714 31166
rect 27694 31218 27746 31230
rect 27694 31154 27746 31166
rect 28142 31218 28194 31230
rect 28142 31154 28194 31166
rect 28702 31218 28754 31230
rect 31826 31166 31838 31218
rect 31890 31166 31902 31218
rect 28702 31154 28754 31166
rect 2606 31106 2658 31118
rect 10110 31106 10162 31118
rect 3042 31054 3054 31106
rect 3106 31054 3118 31106
rect 9426 31054 9438 31106
rect 9490 31103 9502 31106
rect 9762 31103 9774 31106
rect 9490 31057 9774 31103
rect 9490 31054 9502 31057
rect 9762 31054 9774 31057
rect 9826 31054 9838 31106
rect 2606 31042 2658 31054
rect 10110 31042 10162 31054
rect 20414 31106 20466 31118
rect 20414 31042 20466 31054
rect 23102 31106 23154 31118
rect 23102 31042 23154 31054
rect 28366 31106 28418 31118
rect 28366 31042 28418 31054
rect 32286 31106 32338 31118
rect 32286 31042 32338 31054
rect 3726 30994 3778 31006
rect 10222 30994 10274 31006
rect 3266 30942 3278 30994
rect 3330 30942 3342 30994
rect 9874 30942 9886 30994
rect 9938 30942 9950 30994
rect 3726 30930 3778 30942
rect 10222 30930 10274 30942
rect 12238 30994 12290 31006
rect 20638 30994 20690 31006
rect 14130 30942 14142 30994
rect 14194 30942 14206 30994
rect 12238 30930 12290 30942
rect 20638 30930 20690 30942
rect 20974 30994 21026 31006
rect 20974 30930 21026 30942
rect 21310 30994 21362 31006
rect 21310 30930 21362 30942
rect 21982 30994 22034 31006
rect 21982 30930 22034 30942
rect 22206 30994 22258 31006
rect 22206 30930 22258 30942
rect 22654 30994 22706 31006
rect 22654 30930 22706 30942
rect 28030 30994 28082 31006
rect 28030 30930 28082 30942
rect 28478 30994 28530 31006
rect 28478 30930 28530 30942
rect 28814 30994 28866 31006
rect 28814 30930 28866 30942
rect 29150 30994 29202 31006
rect 29150 30930 29202 30942
rect 31502 30994 31554 31006
rect 31502 30930 31554 30942
rect 1822 30882 1874 30894
rect 1822 30818 1874 30830
rect 2382 30882 2434 30894
rect 2382 30818 2434 30830
rect 4622 30882 4674 30894
rect 16158 30882 16210 30894
rect 14354 30830 14366 30882
rect 14418 30830 14430 30882
rect 4622 30818 4674 30830
rect 16158 30818 16210 30830
rect 22430 30882 22482 30894
rect 22430 30818 22482 30830
rect 24222 30882 24274 30894
rect 24222 30818 24274 30830
rect 31054 30882 31106 30894
rect 31054 30818 31106 30830
rect 31278 30882 31330 30894
rect 31278 30818 31330 30830
rect 2718 30770 2770 30782
rect 12014 30770 12066 30782
rect 10658 30718 10670 30770
rect 10722 30718 10734 30770
rect 11666 30718 11678 30770
rect 11730 30718 11742 30770
rect 2718 30706 2770 30718
rect 12014 30706 12066 30718
rect 20302 30770 20354 30782
rect 20302 30706 20354 30718
rect 23214 30770 23266 30782
rect 23426 30718 23438 30770
rect 23490 30767 23502 30770
rect 24210 30767 24222 30770
rect 23490 30721 24222 30767
rect 23490 30718 23502 30721
rect 24210 30718 24222 30721
rect 24274 30718 24286 30770
rect 23214 30706 23266 30718
rect 1344 30602 43568 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 43568 30602
rect 1344 30516 43568 30550
rect 6078 30434 6130 30446
rect 6078 30370 6130 30382
rect 11790 30434 11842 30446
rect 11790 30370 11842 30382
rect 20078 30434 20130 30446
rect 30482 30382 30494 30434
rect 30546 30431 30558 30434
rect 30930 30431 30942 30434
rect 30546 30385 30942 30431
rect 30546 30382 30558 30385
rect 30930 30382 30942 30385
rect 30994 30382 31006 30434
rect 20078 30370 20130 30382
rect 16270 30322 16322 30334
rect 1922 30270 1934 30322
rect 1986 30270 1998 30322
rect 16270 30258 16322 30270
rect 17614 30322 17666 30334
rect 17614 30258 17666 30270
rect 18062 30322 18114 30334
rect 34638 30322 34690 30334
rect 26450 30270 26462 30322
rect 26514 30270 26526 30322
rect 34066 30270 34078 30322
rect 34130 30270 34142 30322
rect 18062 30258 18114 30270
rect 34638 30258 34690 30270
rect 12014 30210 12066 30222
rect 4834 30158 4846 30210
rect 4898 30158 4910 30210
rect 12014 30146 12066 30158
rect 12238 30210 12290 30222
rect 15934 30210 15986 30222
rect 15474 30158 15486 30210
rect 15538 30158 15550 30210
rect 15698 30158 15710 30210
rect 15762 30158 15774 30210
rect 12238 30146 12290 30158
rect 15934 30146 15986 30158
rect 16158 30210 16210 30222
rect 16942 30210 16994 30222
rect 16706 30158 16718 30210
rect 16770 30158 16782 30210
rect 16158 30146 16210 30158
rect 16942 30146 16994 30158
rect 17054 30210 17106 30222
rect 17054 30146 17106 30158
rect 20862 30210 20914 30222
rect 22654 30210 22706 30222
rect 27918 30210 27970 30222
rect 21746 30158 21758 30210
rect 21810 30158 21822 30210
rect 23538 30158 23550 30210
rect 23602 30158 23614 30210
rect 24322 30158 24334 30210
rect 24386 30158 24398 30210
rect 20862 30146 20914 30158
rect 22654 30146 22706 30158
rect 27918 30146 27970 30158
rect 29486 30210 29538 30222
rect 29486 30146 29538 30158
rect 29710 30210 29762 30222
rect 29710 30146 29762 30158
rect 30046 30210 30098 30222
rect 30046 30146 30098 30158
rect 30270 30210 30322 30222
rect 30270 30146 30322 30158
rect 30830 30210 30882 30222
rect 34414 30210 34466 30222
rect 31154 30158 31166 30210
rect 31218 30158 31230 30210
rect 34962 30158 34974 30210
rect 35026 30158 35038 30210
rect 30830 30146 30882 30158
rect 34414 30146 34466 30158
rect 6302 30098 6354 30110
rect 4050 30046 4062 30098
rect 4114 30046 4126 30098
rect 6302 30034 6354 30046
rect 11118 30098 11170 30110
rect 11118 30034 11170 30046
rect 11342 30098 11394 30110
rect 16382 30098 16434 30110
rect 11554 30046 11566 30098
rect 11618 30046 11630 30098
rect 11342 30034 11394 30046
rect 16382 30034 16434 30046
rect 17390 30098 17442 30110
rect 17390 30034 17442 30046
rect 20190 30098 20242 30110
rect 20190 30034 20242 30046
rect 20526 30098 20578 30110
rect 20526 30034 20578 30046
rect 20638 30098 20690 30110
rect 20638 30034 20690 30046
rect 22318 30098 22370 30110
rect 22318 30034 22370 30046
rect 22990 30098 23042 30110
rect 22990 30034 23042 30046
rect 27582 30098 27634 30110
rect 27582 30034 27634 30046
rect 29150 30098 29202 30110
rect 29150 30034 29202 30046
rect 29934 30098 29986 30110
rect 31938 30046 31950 30098
rect 32002 30046 32014 30098
rect 29934 30034 29986 30046
rect 6750 29986 6802 29998
rect 15150 29986 15202 29998
rect 5730 29934 5742 29986
rect 5794 29934 5806 29986
rect 11666 29934 11678 29986
rect 11730 29934 11742 29986
rect 6750 29922 6802 29934
rect 15150 29922 15202 29934
rect 17502 29986 17554 29998
rect 17502 29922 17554 29934
rect 18398 29986 18450 29998
rect 18398 29922 18450 29934
rect 19630 29986 19682 29998
rect 19630 29922 19682 29934
rect 20078 29986 20130 29998
rect 20078 29922 20130 29934
rect 21982 29986 22034 29998
rect 21982 29922 22034 29934
rect 22430 29986 22482 29998
rect 22430 29922 22482 29934
rect 26798 29986 26850 29998
rect 27694 29986 27746 29998
rect 27122 29934 27134 29986
rect 27186 29934 27198 29986
rect 26798 29922 26850 29934
rect 27694 29922 27746 29934
rect 28254 29986 28306 29998
rect 28254 29922 28306 29934
rect 29262 29986 29314 29998
rect 29262 29922 29314 29934
rect 1344 29818 43568 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 43568 29818
rect 1344 29732 43568 29766
rect 2046 29650 2098 29662
rect 2046 29586 2098 29598
rect 2606 29650 2658 29662
rect 2606 29586 2658 29598
rect 3838 29650 3890 29662
rect 3838 29586 3890 29598
rect 4174 29650 4226 29662
rect 4174 29586 4226 29598
rect 17726 29650 17778 29662
rect 21198 29650 21250 29662
rect 20738 29598 20750 29650
rect 20802 29598 20814 29650
rect 26562 29598 26574 29650
rect 26626 29598 26638 29650
rect 17726 29586 17778 29598
rect 21198 29586 21250 29598
rect 2494 29538 2546 29550
rect 2494 29474 2546 29486
rect 2718 29538 2770 29550
rect 2718 29474 2770 29486
rect 3054 29538 3106 29550
rect 3054 29474 3106 29486
rect 4846 29538 4898 29550
rect 6078 29538 6130 29550
rect 5282 29486 5294 29538
rect 5346 29535 5358 29538
rect 5506 29535 5518 29538
rect 5346 29489 5518 29535
rect 5346 29486 5358 29489
rect 5506 29486 5518 29489
rect 5570 29486 5582 29538
rect 4846 29474 4898 29486
rect 6078 29474 6130 29486
rect 16718 29538 16770 29550
rect 16718 29474 16770 29486
rect 17838 29538 17890 29550
rect 17838 29474 17890 29486
rect 18062 29538 18114 29550
rect 18062 29474 18114 29486
rect 19070 29538 19122 29550
rect 19070 29474 19122 29486
rect 6190 29426 6242 29438
rect 1810 29374 1822 29426
rect 1874 29374 1886 29426
rect 3266 29374 3278 29426
rect 3330 29374 3342 29426
rect 3826 29374 3838 29426
rect 3890 29374 3902 29426
rect 4386 29374 4398 29426
rect 4450 29374 4462 29426
rect 5170 29374 5182 29426
rect 5234 29374 5246 29426
rect 6190 29362 6242 29374
rect 10110 29426 10162 29438
rect 10110 29362 10162 29374
rect 10334 29426 10386 29438
rect 16606 29426 16658 29438
rect 15362 29374 15374 29426
rect 15426 29374 15438 29426
rect 10334 29362 10386 29374
rect 16606 29362 16658 29374
rect 16942 29426 16994 29438
rect 17614 29426 17666 29438
rect 17378 29374 17390 29426
rect 17442 29374 17454 29426
rect 16942 29362 16994 29374
rect 17614 29362 17666 29374
rect 20414 29426 20466 29438
rect 20414 29362 20466 29374
rect 26238 29426 26290 29438
rect 26238 29362 26290 29374
rect 5630 29314 5682 29326
rect 5630 29250 5682 29262
rect 6638 29314 6690 29326
rect 18510 29314 18562 29326
rect 11778 29262 11790 29314
rect 11842 29262 11854 29314
rect 6638 29250 6690 29262
rect 18510 29250 18562 29262
rect 27134 29314 27186 29326
rect 27134 29250 27186 29262
rect 28926 29314 28978 29326
rect 28926 29250 28978 29262
rect 34078 29314 34130 29326
rect 34078 29250 34130 29262
rect 5182 29202 5234 29214
rect 3602 29150 3614 29202
rect 3666 29150 3678 29202
rect 5182 29138 5234 29150
rect 6078 29202 6130 29214
rect 9762 29150 9774 29202
rect 9826 29150 9838 29202
rect 6078 29138 6130 29150
rect 1344 29034 43568 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 43568 29034
rect 1344 28948 43568 28982
rect 4622 28866 4674 28878
rect 4622 28802 4674 28814
rect 11342 28866 11394 28878
rect 11342 28802 11394 28814
rect 17950 28866 18002 28878
rect 17950 28802 18002 28814
rect 30830 28866 30882 28878
rect 30830 28802 30882 28814
rect 1934 28754 1986 28766
rect 26910 28754 26962 28766
rect 6290 28702 6302 28754
rect 6354 28702 6366 28754
rect 1934 28690 1986 28702
rect 26910 28690 26962 28702
rect 33742 28754 33794 28766
rect 33742 28690 33794 28702
rect 10334 28642 10386 28654
rect 4274 28590 4286 28642
rect 4338 28590 4350 28642
rect 8418 28590 8430 28642
rect 8482 28590 8494 28642
rect 9090 28590 9102 28642
rect 9154 28590 9166 28642
rect 10334 28578 10386 28590
rect 10446 28642 10498 28654
rect 10446 28578 10498 28590
rect 10894 28642 10946 28654
rect 10894 28578 10946 28590
rect 11118 28642 11170 28654
rect 11118 28578 11170 28590
rect 11454 28642 11506 28654
rect 11454 28578 11506 28590
rect 11902 28642 11954 28654
rect 13918 28642 13970 28654
rect 13458 28590 13470 28642
rect 13522 28590 13534 28642
rect 11902 28578 11954 28590
rect 13918 28578 13970 28590
rect 14142 28642 14194 28654
rect 14142 28578 14194 28590
rect 17390 28642 17442 28654
rect 17390 28578 17442 28590
rect 17726 28642 17778 28654
rect 20638 28642 20690 28654
rect 26014 28642 26066 28654
rect 18274 28590 18286 28642
rect 18338 28590 18350 28642
rect 25554 28590 25566 28642
rect 25618 28590 25630 28642
rect 17726 28578 17778 28590
rect 20638 28578 20690 28590
rect 26014 28578 26066 28590
rect 27246 28642 27298 28654
rect 27246 28578 27298 28590
rect 29486 28642 29538 28654
rect 29486 28578 29538 28590
rect 29822 28642 29874 28654
rect 29822 28578 29874 28590
rect 30158 28642 30210 28654
rect 30158 28578 30210 28590
rect 30494 28642 30546 28654
rect 30494 28578 30546 28590
rect 32734 28642 32786 28654
rect 32734 28578 32786 28590
rect 32846 28642 32898 28654
rect 32846 28578 32898 28590
rect 4958 28530 5010 28542
rect 4958 28466 5010 28478
rect 12238 28530 12290 28542
rect 12238 28466 12290 28478
rect 14030 28530 14082 28542
rect 27806 28530 27858 28542
rect 16258 28478 16270 28530
rect 16322 28478 16334 28530
rect 16930 28478 16942 28530
rect 16994 28478 17006 28530
rect 25330 28478 25342 28530
rect 25394 28478 25406 28530
rect 26338 28478 26350 28530
rect 26402 28478 26414 28530
rect 14030 28466 14082 28478
rect 27806 28466 27858 28478
rect 29150 28530 29202 28542
rect 29150 28466 29202 28478
rect 30718 28530 30770 28542
rect 30718 28466 30770 28478
rect 4734 28418 4786 28430
rect 4734 28354 4786 28366
rect 10782 28418 10834 28430
rect 10782 28354 10834 28366
rect 15150 28418 15202 28430
rect 15150 28354 15202 28366
rect 15598 28418 15650 28430
rect 15598 28354 15650 28366
rect 15934 28418 15986 28430
rect 15934 28354 15986 28366
rect 16606 28418 16658 28430
rect 27358 28418 27410 28430
rect 20290 28366 20302 28418
rect 20354 28366 20366 28418
rect 16606 28354 16658 28366
rect 27358 28354 27410 28366
rect 27582 28418 27634 28430
rect 27582 28354 27634 28366
rect 27918 28418 27970 28430
rect 27918 28354 27970 28366
rect 28142 28418 28194 28430
rect 28142 28354 28194 28366
rect 28590 28418 28642 28430
rect 28590 28354 28642 28366
rect 29262 28418 29314 28430
rect 29262 28354 29314 28366
rect 30270 28418 30322 28430
rect 30270 28354 30322 28366
rect 30830 28418 30882 28430
rect 30830 28354 30882 28366
rect 31502 28418 31554 28430
rect 31502 28354 31554 28366
rect 33294 28418 33346 28430
rect 33294 28354 33346 28366
rect 1344 28250 43568 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 43568 28250
rect 1344 28164 43568 28198
rect 12910 28082 12962 28094
rect 11666 28030 11678 28082
rect 11730 28030 11742 28082
rect 12910 28018 12962 28030
rect 16270 28082 16322 28094
rect 16270 28018 16322 28030
rect 17502 28082 17554 28094
rect 17502 28018 17554 28030
rect 12462 27970 12514 27982
rect 10770 27918 10782 27970
rect 10834 27918 10846 27970
rect 12462 27906 12514 27918
rect 22206 27970 22258 27982
rect 30930 27918 30942 27970
rect 30994 27918 31006 27970
rect 33842 27918 33854 27970
rect 33906 27918 33918 27970
rect 22206 27906 22258 27918
rect 11118 27858 11170 27870
rect 12126 27858 12178 27870
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 10546 27806 10558 27858
rect 10610 27806 10622 27858
rect 11778 27806 11790 27858
rect 11842 27806 11854 27858
rect 11118 27794 11170 27806
rect 12126 27794 12178 27806
rect 21646 27858 21698 27870
rect 21646 27794 21698 27806
rect 21870 27858 21922 27870
rect 27234 27806 27246 27858
rect 27298 27806 27310 27858
rect 33058 27806 33070 27858
rect 33122 27806 33134 27858
rect 21870 27794 21922 27806
rect 4734 27746 4786 27758
rect 4734 27682 4786 27694
rect 11342 27746 11394 27758
rect 11342 27682 11394 27694
rect 12350 27746 12402 27758
rect 12350 27682 12402 27694
rect 21758 27746 21810 27758
rect 21758 27682 21810 27694
rect 26910 27746 26962 27758
rect 35970 27694 35982 27746
rect 36034 27694 36046 27746
rect 26910 27682 26962 27694
rect 1934 27634 1986 27646
rect 1934 27570 1986 27582
rect 11566 27634 11618 27646
rect 11566 27570 11618 27582
rect 1344 27466 43568 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 43568 27466
rect 1344 27380 43568 27414
rect 29374 27298 29426 27310
rect 30158 27298 30210 27310
rect 15138 27246 15150 27298
rect 15202 27246 15214 27298
rect 29698 27246 29710 27298
rect 29762 27246 29774 27298
rect 29374 27234 29426 27246
rect 30158 27234 30210 27246
rect 34414 27298 34466 27310
rect 34738 27246 34750 27298
rect 34802 27246 34814 27298
rect 34414 27234 34466 27246
rect 16718 27186 16770 27198
rect 35198 27186 35250 27198
rect 2034 27134 2046 27186
rect 2098 27134 2110 27186
rect 9986 27134 9998 27186
rect 10050 27134 10062 27186
rect 12114 27134 12126 27186
rect 12178 27134 12190 27186
rect 22642 27134 22654 27186
rect 22706 27134 22718 27186
rect 24770 27134 24782 27186
rect 24834 27134 24846 27186
rect 25666 27134 25678 27186
rect 25730 27134 25742 27186
rect 33618 27134 33630 27186
rect 33682 27134 33694 27186
rect 16718 27122 16770 27134
rect 35198 27122 35250 27134
rect 6750 27074 6802 27086
rect 4162 27022 4174 27074
rect 4226 27022 4238 27074
rect 6750 27010 6802 27022
rect 7870 27074 7922 27086
rect 14814 27074 14866 27086
rect 12786 27022 12798 27074
rect 12850 27022 12862 27074
rect 7870 27010 7922 27022
rect 14814 27010 14866 27022
rect 15710 27074 15762 27086
rect 16494 27074 16546 27086
rect 20526 27074 20578 27086
rect 15922 27022 15934 27074
rect 15986 27022 15998 27074
rect 17154 27022 17166 27074
rect 17218 27022 17230 27074
rect 15710 27010 15762 27022
rect 16494 27010 16546 27022
rect 20526 27010 20578 27022
rect 21310 27074 21362 27086
rect 21310 27010 21362 27022
rect 21646 27074 21698 27086
rect 25230 27074 25282 27086
rect 29150 27074 29202 27086
rect 21970 27022 21982 27074
rect 22034 27022 22046 27074
rect 28578 27022 28590 27074
rect 28642 27022 28654 27074
rect 21646 27010 21698 27022
rect 25230 27010 25282 27022
rect 29150 27010 29202 27022
rect 30046 27074 30098 27086
rect 34190 27074 34242 27086
rect 30818 27022 30830 27074
rect 30882 27022 30894 27074
rect 30046 27010 30098 27022
rect 34190 27010 34242 27022
rect 14478 26962 14530 26974
rect 7522 26910 7534 26962
rect 7586 26910 7598 26962
rect 14478 26898 14530 26910
rect 15598 26962 15650 26974
rect 15598 26898 15650 26910
rect 16270 26962 16322 26974
rect 20638 26962 20690 26974
rect 16930 26910 16942 26962
rect 16994 26910 17006 26962
rect 27794 26910 27806 26962
rect 27858 26910 27870 26962
rect 31490 26910 31502 26962
rect 31554 26910 31566 26962
rect 16270 26898 16322 26910
rect 20638 26898 20690 26910
rect 6862 26850 6914 26862
rect 6862 26786 6914 26798
rect 16158 26850 16210 26862
rect 16158 26786 16210 26798
rect 17726 26850 17778 26862
rect 17726 26786 17778 26798
rect 20862 26850 20914 26862
rect 20862 26786 20914 26798
rect 21422 26850 21474 26862
rect 21422 26786 21474 26798
rect 30158 26850 30210 26862
rect 30158 26786 30210 26798
rect 1344 26682 43568 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 43568 26682
rect 1344 26596 43568 26630
rect 6974 26514 7026 26526
rect 6974 26450 7026 26462
rect 15486 26514 15538 26526
rect 15486 26450 15538 26462
rect 16270 26514 16322 26526
rect 27806 26514 27858 26526
rect 25778 26462 25790 26514
rect 25842 26462 25854 26514
rect 16270 26450 16322 26462
rect 27806 26450 27858 26462
rect 28814 26514 28866 26526
rect 28814 26450 28866 26462
rect 29262 26514 29314 26526
rect 29262 26450 29314 26462
rect 34302 26514 34354 26526
rect 34302 26450 34354 26462
rect 7086 26402 7138 26414
rect 5842 26350 5854 26402
rect 5906 26350 5918 26402
rect 7086 26338 7138 26350
rect 7982 26402 8034 26414
rect 16382 26402 16434 26414
rect 15810 26350 15822 26402
rect 15874 26350 15886 26402
rect 7982 26338 8034 26350
rect 16382 26338 16434 26350
rect 18062 26402 18114 26414
rect 18062 26338 18114 26350
rect 27358 26402 27410 26414
rect 27358 26338 27410 26350
rect 27582 26402 27634 26414
rect 27582 26338 27634 26350
rect 7310 26290 7362 26302
rect 11566 26290 11618 26302
rect 12126 26290 12178 26302
rect 6514 26238 6526 26290
rect 6578 26238 6590 26290
rect 7746 26238 7758 26290
rect 7810 26238 7822 26290
rect 11890 26238 11902 26290
rect 11954 26238 11966 26290
rect 7310 26226 7362 26238
rect 11566 26226 11618 26238
rect 12126 26226 12178 26238
rect 12350 26290 12402 26302
rect 12350 26226 12402 26238
rect 12574 26290 12626 26302
rect 12574 26226 12626 26238
rect 16606 26290 16658 26302
rect 22766 26290 22818 26302
rect 16818 26238 16830 26290
rect 16882 26238 16894 26290
rect 22530 26238 22542 26290
rect 22594 26238 22606 26290
rect 16606 26226 16658 26238
rect 22766 26226 22818 26238
rect 23214 26290 23266 26302
rect 23214 26226 23266 26238
rect 23326 26290 23378 26302
rect 23326 26226 23378 26238
rect 25454 26290 25506 26302
rect 25454 26226 25506 26238
rect 28030 26290 28082 26302
rect 28030 26226 28082 26238
rect 11342 26178 11394 26190
rect 3714 26126 3726 26178
rect 3778 26126 3790 26178
rect 11342 26114 11394 26126
rect 12462 26178 12514 26190
rect 12462 26114 12514 26126
rect 13022 26178 13074 26190
rect 17502 26178 17554 26190
rect 22990 26178 23042 26190
rect 16258 26126 16270 26178
rect 16322 26126 16334 26178
rect 19618 26126 19630 26178
rect 19682 26126 19694 26178
rect 21746 26126 21758 26178
rect 21810 26126 21822 26178
rect 13022 26114 13074 26126
rect 17502 26114 17554 26126
rect 22990 26114 23042 26126
rect 25230 26178 25282 26190
rect 25230 26114 25282 26126
rect 33854 26178 33906 26190
rect 33854 26114 33906 26126
rect 7534 26066 7586 26078
rect 7534 26002 7586 26014
rect 1344 25898 43568 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 43568 25898
rect 1344 25812 43568 25846
rect 22318 25730 22370 25742
rect 22318 25666 22370 25678
rect 27134 25730 27186 25742
rect 27134 25666 27186 25678
rect 5854 25618 5906 25630
rect 1698 25566 1710 25618
rect 1762 25566 1774 25618
rect 5854 25554 5906 25566
rect 7310 25618 7362 25630
rect 7310 25554 7362 25566
rect 23102 25618 23154 25630
rect 23102 25554 23154 25566
rect 32174 25618 32226 25630
rect 32174 25554 32226 25566
rect 7086 25506 7138 25518
rect 4610 25454 4622 25506
rect 4674 25454 4686 25506
rect 7086 25442 7138 25454
rect 7534 25506 7586 25518
rect 7534 25442 7586 25454
rect 8094 25506 8146 25518
rect 8094 25442 8146 25454
rect 12350 25506 12402 25518
rect 12350 25442 12402 25454
rect 12462 25506 12514 25518
rect 12462 25442 12514 25454
rect 15598 25506 15650 25518
rect 15598 25442 15650 25454
rect 20526 25506 20578 25518
rect 20526 25442 20578 25454
rect 21646 25506 21698 25518
rect 21646 25442 21698 25454
rect 22094 25506 22146 25518
rect 31614 25506 31666 25518
rect 22642 25454 22654 25506
rect 22706 25454 22718 25506
rect 22094 25442 22146 25454
rect 31614 25442 31666 25454
rect 5742 25394 5794 25406
rect 12574 25394 12626 25406
rect 3826 25342 3838 25394
rect 3890 25342 3902 25394
rect 7746 25342 7758 25394
rect 7810 25342 7822 25394
rect 5742 25330 5794 25342
rect 12574 25330 12626 25342
rect 15710 25394 15762 25406
rect 21310 25394 21362 25406
rect 16706 25342 16718 25394
rect 16770 25342 16782 25394
rect 15710 25330 15762 25342
rect 21310 25330 21362 25342
rect 21422 25394 21474 25406
rect 21422 25330 21474 25342
rect 27022 25394 27074 25406
rect 27022 25330 27074 25342
rect 6974 25282 7026 25294
rect 6974 25218 7026 25230
rect 10558 25282 10610 25294
rect 15262 25282 15314 25294
rect 11890 25230 11902 25282
rect 11954 25230 11966 25282
rect 10558 25218 10610 25230
rect 15262 25218 15314 25230
rect 16494 25282 16546 25294
rect 16494 25218 16546 25230
rect 17054 25282 17106 25294
rect 17054 25218 17106 25230
rect 17502 25282 17554 25294
rect 17502 25218 17554 25230
rect 19854 25282 19906 25294
rect 19854 25218 19906 25230
rect 20302 25282 20354 25294
rect 20302 25218 20354 25230
rect 20638 25282 20690 25294
rect 20638 25218 20690 25230
rect 20862 25282 20914 25294
rect 20862 25218 20914 25230
rect 31726 25282 31778 25294
rect 31726 25218 31778 25230
rect 33854 25282 33906 25294
rect 33854 25218 33906 25230
rect 1344 25114 43568 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 43568 25114
rect 1344 25028 43568 25062
rect 12686 24946 12738 24958
rect 10546 24894 10558 24946
rect 10610 24894 10622 24946
rect 12686 24882 12738 24894
rect 12798 24946 12850 24958
rect 12798 24882 12850 24894
rect 13470 24946 13522 24958
rect 13470 24882 13522 24894
rect 15150 24946 15202 24958
rect 15150 24882 15202 24894
rect 15262 24946 15314 24958
rect 15262 24882 15314 24894
rect 16606 24946 16658 24958
rect 20078 24946 20130 24958
rect 17602 24894 17614 24946
rect 17666 24894 17678 24946
rect 16606 24882 16658 24894
rect 20078 24882 20130 24894
rect 23438 24946 23490 24958
rect 23438 24882 23490 24894
rect 23886 24946 23938 24958
rect 23886 24882 23938 24894
rect 28926 24946 28978 24958
rect 28926 24882 28978 24894
rect 33182 24946 33234 24958
rect 33182 24882 33234 24894
rect 6750 24834 6802 24846
rect 6750 24770 6802 24782
rect 7646 24834 7698 24846
rect 7646 24770 7698 24782
rect 9550 24834 9602 24846
rect 9550 24770 9602 24782
rect 9998 24834 10050 24846
rect 9998 24770 10050 24782
rect 15486 24834 15538 24846
rect 15486 24770 15538 24782
rect 16830 24834 16882 24846
rect 16830 24770 16882 24782
rect 19294 24834 19346 24846
rect 19294 24770 19346 24782
rect 19630 24834 19682 24846
rect 19630 24770 19682 24782
rect 34302 24834 34354 24846
rect 34302 24770 34354 24782
rect 7310 24722 7362 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 7310 24658 7362 24670
rect 9774 24722 9826 24734
rect 9774 24658 9826 24670
rect 10110 24722 10162 24734
rect 10110 24658 10162 24670
rect 10894 24722 10946 24734
rect 12462 24722 12514 24734
rect 12226 24670 12238 24722
rect 12290 24670 12302 24722
rect 10894 24658 10946 24670
rect 12462 24658 12514 24670
rect 12574 24722 12626 24734
rect 15038 24722 15090 24734
rect 16382 24722 16434 24734
rect 14802 24670 14814 24722
rect 14866 24670 14878 24722
rect 16146 24670 16158 24722
rect 16210 24670 16222 24722
rect 12574 24658 12626 24670
rect 15038 24658 15090 24670
rect 16382 24658 16434 24670
rect 17950 24722 18002 24734
rect 17950 24658 18002 24670
rect 18286 24722 18338 24734
rect 18286 24658 18338 24670
rect 23326 24722 23378 24734
rect 28466 24670 28478 24722
rect 28530 24670 28542 24722
rect 29362 24670 29374 24722
rect 29426 24670 29438 24722
rect 33954 24719 33966 24722
rect 33745 24673 33966 24719
rect 23326 24658 23378 24670
rect 6862 24610 6914 24622
rect 6862 24546 6914 24558
rect 6974 24610 7026 24622
rect 6974 24546 7026 24558
rect 9886 24610 9938 24622
rect 9886 24546 9938 24558
rect 11118 24610 11170 24622
rect 11118 24546 11170 24558
rect 11902 24610 11954 24622
rect 11902 24546 11954 24558
rect 14590 24610 14642 24622
rect 14590 24546 14642 24558
rect 16494 24610 16546 24622
rect 16494 24546 16546 24558
rect 18846 24610 18898 24622
rect 33630 24610 33682 24622
rect 25554 24558 25566 24610
rect 25618 24558 25630 24610
rect 27682 24558 27694 24610
rect 27746 24558 27758 24610
rect 30146 24558 30158 24610
rect 30210 24558 30222 24610
rect 32274 24558 32286 24610
rect 32338 24558 32350 24610
rect 18846 24546 18898 24558
rect 33630 24546 33682 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 7198 24498 7250 24510
rect 33618 24446 33630 24498
rect 33682 24495 33694 24498
rect 33745 24495 33791 24673
rect 33954 24670 33966 24673
rect 34018 24670 34030 24722
rect 33682 24449 33791 24495
rect 34078 24498 34130 24510
rect 33682 24446 33694 24449
rect 7198 24434 7250 24446
rect 34078 24434 34130 24446
rect 34414 24498 34466 24510
rect 34414 24434 34466 24446
rect 1344 24330 43568 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 43568 24330
rect 1344 24244 43568 24278
rect 5742 24162 5794 24174
rect 5742 24098 5794 24110
rect 11678 24050 11730 24062
rect 1698 23998 1710 24050
rect 1762 23998 1774 24050
rect 3826 23998 3838 24050
rect 3890 23998 3902 24050
rect 11106 23998 11118 24050
rect 11170 23998 11182 24050
rect 11678 23986 11730 23998
rect 16494 24050 16546 24062
rect 16494 23986 16546 23998
rect 29374 24050 29426 24062
rect 29374 23986 29426 23998
rect 32958 24050 33010 24062
rect 32958 23986 33010 23998
rect 36206 24050 36258 24062
rect 36206 23986 36258 23998
rect 9886 23938 9938 23950
rect 4610 23886 4622 23938
rect 4674 23886 4686 23938
rect 9886 23874 9938 23886
rect 10110 23938 10162 23950
rect 10110 23874 10162 23886
rect 10334 23938 10386 23950
rect 11454 23938 11506 23950
rect 10546 23886 10558 23938
rect 10610 23886 10622 23938
rect 10334 23874 10386 23886
rect 11454 23874 11506 23886
rect 16046 23938 16098 23950
rect 16046 23874 16098 23886
rect 17166 23938 17218 23950
rect 17166 23874 17218 23886
rect 17502 23938 17554 23950
rect 17502 23874 17554 23886
rect 18622 23938 18674 23950
rect 18622 23874 18674 23886
rect 29710 23938 29762 23950
rect 33282 23886 33294 23938
rect 33346 23886 33358 23938
rect 29710 23874 29762 23886
rect 5630 23826 5682 23838
rect 5630 23762 5682 23774
rect 10782 23826 10834 23838
rect 10782 23762 10834 23774
rect 15486 23826 15538 23838
rect 16818 23774 16830 23826
rect 16882 23774 16894 23826
rect 34066 23774 34078 23826
rect 34130 23774 34142 23826
rect 15486 23762 15538 23774
rect 9774 23714 9826 23726
rect 9774 23650 9826 23662
rect 15150 23714 15202 23726
rect 15150 23650 15202 23662
rect 17614 23714 17666 23726
rect 17614 23650 17666 23662
rect 17838 23714 17890 23726
rect 18274 23662 18286 23714
rect 18338 23662 18350 23714
rect 30034 23662 30046 23714
rect 30098 23662 30110 23714
rect 17838 23650 17890 23662
rect 1344 23546 43568 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 43568 23546
rect 1344 23460 43568 23494
rect 8430 23378 8482 23390
rect 8430 23314 8482 23326
rect 20190 23378 20242 23390
rect 30942 23378 30994 23390
rect 29474 23326 29486 23378
rect 29538 23326 29550 23378
rect 20190 23314 20242 23326
rect 30942 23314 30994 23326
rect 32510 23378 32562 23390
rect 32510 23314 32562 23326
rect 33294 23378 33346 23390
rect 33294 23314 33346 23326
rect 42814 23378 42866 23390
rect 42814 23314 42866 23326
rect 20078 23266 20130 23278
rect 5730 23214 5742 23266
rect 5794 23214 5806 23266
rect 34514 23214 34526 23266
rect 34578 23214 34590 23266
rect 20078 23202 20130 23214
rect 29822 23154 29874 23166
rect 6514 23102 6526 23154
rect 6578 23102 6590 23154
rect 28690 23102 28702 23154
rect 28754 23102 28766 23154
rect 29026 23102 29038 23154
rect 29090 23102 29102 23154
rect 29586 23102 29598 23154
rect 29650 23102 29662 23154
rect 29822 23090 29874 23102
rect 30158 23154 30210 23166
rect 30158 23090 30210 23102
rect 30494 23154 30546 23166
rect 43150 23154 43202 23166
rect 30706 23102 30718 23154
rect 30770 23102 30782 23154
rect 33058 23102 33070 23154
rect 33122 23102 33134 23154
rect 33730 23102 33742 23154
rect 33794 23102 33806 23154
rect 30494 23090 30546 23102
rect 43150 23090 43202 23102
rect 8318 23042 8370 23054
rect 3602 22990 3614 23042
rect 3666 22990 3678 23042
rect 8318 22978 8370 22990
rect 10670 23042 10722 23054
rect 10670 22978 10722 22990
rect 27358 23042 27410 23054
rect 27358 22978 27410 22990
rect 28030 23042 28082 23054
rect 28030 22978 28082 22990
rect 31390 23042 31442 23054
rect 42590 23042 42642 23054
rect 36642 22990 36654 23042
rect 36706 22990 36718 23042
rect 31390 22978 31442 22990
rect 42590 22978 42642 22990
rect 28366 22930 28418 22942
rect 28366 22866 28418 22878
rect 28702 22930 28754 22942
rect 30606 22930 30658 22942
rect 29250 22878 29262 22930
rect 29314 22878 29326 22930
rect 28702 22866 28754 22878
rect 30606 22866 30658 22878
rect 33406 22930 33458 22942
rect 33406 22866 33458 22878
rect 1344 22762 43568 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 43568 22762
rect 1344 22676 43568 22710
rect 1934 22594 1986 22606
rect 1934 22530 1986 22542
rect 29486 22594 29538 22606
rect 29486 22530 29538 22542
rect 9326 22482 9378 22494
rect 11118 22482 11170 22494
rect 10210 22430 10222 22482
rect 10274 22430 10286 22482
rect 9326 22418 9378 22430
rect 11118 22418 11170 22430
rect 12014 22482 12066 22494
rect 12014 22418 12066 22430
rect 20750 22482 20802 22494
rect 29934 22482 29986 22494
rect 25554 22430 25566 22482
rect 25618 22430 25630 22482
rect 27682 22430 27694 22482
rect 27746 22430 27758 22482
rect 20750 22418 20802 22430
rect 29934 22418 29986 22430
rect 33742 22482 33794 22494
rect 33742 22418 33794 22430
rect 34750 22482 34802 22494
rect 34750 22418 34802 22430
rect 10110 22370 10162 22382
rect 10670 22370 10722 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 9650 22318 9662 22370
rect 9714 22318 9726 22370
rect 10322 22318 10334 22370
rect 10386 22318 10398 22370
rect 10110 22306 10162 22318
rect 10670 22306 10722 22318
rect 10894 22370 10946 22382
rect 10894 22306 10946 22318
rect 11678 22370 11730 22382
rect 26910 22370 26962 22382
rect 27358 22370 27410 22382
rect 21410 22318 21422 22370
rect 21474 22318 21486 22370
rect 22754 22318 22766 22370
rect 22818 22318 22830 22370
rect 26786 22318 26798 22370
rect 26850 22318 26862 22370
rect 27122 22318 27134 22370
rect 27186 22318 27198 22370
rect 11678 22306 11730 22318
rect 26910 22306 26962 22318
rect 27358 22306 27410 22318
rect 33854 22370 33906 22382
rect 33854 22306 33906 22318
rect 34190 22370 34242 22382
rect 35422 22370 35474 22382
rect 34962 22318 34974 22370
rect 35026 22318 35038 22370
rect 34190 22306 34242 22318
rect 35422 22306 35474 22318
rect 14926 22258 14978 22270
rect 28030 22258 28082 22270
rect 11330 22206 11342 22258
rect 11394 22206 11406 22258
rect 21298 22206 21310 22258
rect 21362 22206 21374 22258
rect 21746 22206 21758 22258
rect 21810 22206 21822 22258
rect 23426 22206 23438 22258
rect 23490 22206 23502 22258
rect 14926 22194 14978 22206
rect 28030 22194 28082 22206
rect 28590 22258 28642 22270
rect 28590 22194 28642 22206
rect 29150 22258 29202 22270
rect 29150 22194 29202 22206
rect 33630 22258 33682 22270
rect 33630 22194 33682 22206
rect 34638 22258 34690 22270
rect 34638 22194 34690 22206
rect 9886 22146 9938 22158
rect 9886 22082 9938 22094
rect 10558 22146 10610 22158
rect 10558 22082 10610 22094
rect 14590 22146 14642 22158
rect 14590 22082 14642 22094
rect 15038 22146 15090 22158
rect 15038 22082 15090 22094
rect 15262 22146 15314 22158
rect 15262 22082 15314 22094
rect 26014 22146 26066 22158
rect 27806 22146 27858 22158
rect 27010 22094 27022 22146
rect 27074 22094 27086 22146
rect 26014 22082 26066 22094
rect 27806 22082 27858 22094
rect 29374 22146 29426 22158
rect 29374 22082 29426 22094
rect 30382 22146 30434 22158
rect 30382 22082 30434 22094
rect 1344 21978 43568 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 43568 21978
rect 1344 21892 43568 21926
rect 10110 21810 10162 21822
rect 10110 21746 10162 21758
rect 11342 21810 11394 21822
rect 11342 21746 11394 21758
rect 11790 21810 11842 21822
rect 11790 21746 11842 21758
rect 17614 21810 17666 21822
rect 17614 21746 17666 21758
rect 18174 21810 18226 21822
rect 18174 21746 18226 21758
rect 27022 21810 27074 21822
rect 27022 21746 27074 21758
rect 27694 21810 27746 21822
rect 27694 21746 27746 21758
rect 34414 21810 34466 21822
rect 34414 21746 34466 21758
rect 9998 21698 10050 21710
rect 9998 21634 10050 21646
rect 10894 21698 10946 21710
rect 27358 21698 27410 21710
rect 16258 21646 16270 21698
rect 16322 21646 16334 21698
rect 19282 21646 19294 21698
rect 19346 21646 19358 21698
rect 25890 21646 25902 21698
rect 25954 21646 25966 21698
rect 10894 21634 10946 21646
rect 27358 21634 27410 21646
rect 28142 21698 28194 21710
rect 28142 21634 28194 21646
rect 28366 21698 28418 21710
rect 28366 21634 28418 21646
rect 15934 21586 15986 21598
rect 4162 21534 4174 21586
rect 4226 21534 4238 21586
rect 8978 21534 8990 21586
rect 9042 21534 9054 21586
rect 10658 21534 10670 21586
rect 10722 21534 10734 21586
rect 12786 21534 12798 21586
rect 12850 21534 12862 21586
rect 15934 21522 15986 21534
rect 17502 21586 17554 21598
rect 26686 21586 26738 21598
rect 24322 21534 24334 21586
rect 24386 21534 24398 21586
rect 25330 21534 25342 21586
rect 25394 21534 25406 21586
rect 17502 21522 17554 21534
rect 26686 21522 26738 21534
rect 28814 21586 28866 21598
rect 28814 21522 28866 21534
rect 1934 21474 1986 21486
rect 1934 21410 1986 21422
rect 5070 21474 5122 21486
rect 5070 21410 5122 21422
rect 5182 21474 5234 21486
rect 10222 21474 10274 21486
rect 6066 21422 6078 21474
rect 6130 21422 6142 21474
rect 8194 21422 8206 21474
rect 8258 21422 8270 21474
rect 5182 21410 5234 21422
rect 10222 21410 10274 21422
rect 11230 21474 11282 21486
rect 16830 21474 16882 21486
rect 13458 21422 13470 21474
rect 13522 21422 13534 21474
rect 15586 21422 15598 21474
rect 15650 21422 15662 21474
rect 11230 21410 11282 21422
rect 16830 21410 16882 21422
rect 29374 21474 29426 21486
rect 29374 21410 29426 21422
rect 31838 21474 31890 21486
rect 31838 21410 31890 21422
rect 10446 21362 10498 21374
rect 10446 21298 10498 21310
rect 17614 21362 17666 21374
rect 17614 21298 17666 21310
rect 25790 21362 25842 21374
rect 25790 21298 25842 21310
rect 28030 21362 28082 21374
rect 28030 21298 28082 21310
rect 1344 21194 43568 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 43568 21194
rect 1344 21108 43568 21142
rect 27470 21026 27522 21038
rect 27470 20962 27522 20974
rect 29934 21026 29986 21038
rect 29934 20962 29986 20974
rect 31838 21026 31890 21038
rect 31838 20962 31890 20974
rect 32174 21026 32226 21038
rect 32174 20962 32226 20974
rect 12910 20914 12962 20926
rect 1698 20862 1710 20914
rect 1762 20862 1774 20914
rect 3826 20862 3838 20914
rect 3890 20862 3902 20914
rect 12910 20850 12962 20862
rect 14254 20914 14306 20926
rect 25230 20914 25282 20926
rect 18274 20862 18286 20914
rect 18338 20862 18350 20914
rect 14254 20850 14306 20862
rect 25230 20850 25282 20862
rect 25678 20914 25730 20926
rect 25678 20850 25730 20862
rect 28366 20914 28418 20926
rect 28366 20850 28418 20862
rect 30942 20914 30994 20926
rect 35086 20914 35138 20926
rect 31490 20862 31502 20914
rect 31554 20862 31566 20914
rect 30942 20850 30994 20862
rect 35086 20850 35138 20862
rect 12574 20802 12626 20814
rect 16942 20802 16994 20814
rect 18846 20802 18898 20814
rect 21646 20802 21698 20814
rect 22990 20802 23042 20814
rect 4610 20750 4622 20802
rect 4674 20750 4686 20802
rect 14914 20750 14926 20802
rect 14978 20750 14990 20802
rect 15698 20750 15710 20802
rect 15762 20750 15774 20802
rect 15922 20750 15934 20802
rect 15986 20750 15998 20802
rect 17826 20750 17838 20802
rect 17890 20750 17902 20802
rect 21522 20750 21534 20802
rect 21586 20750 21598 20802
rect 21858 20750 21870 20802
rect 21922 20750 21934 20802
rect 12574 20738 12626 20750
rect 16942 20738 16994 20750
rect 18846 20738 18898 20750
rect 21646 20738 21698 20750
rect 22990 20738 23042 20750
rect 23102 20802 23154 20814
rect 24110 20802 24162 20814
rect 23314 20750 23326 20802
rect 23378 20750 23390 20802
rect 23102 20738 23154 20750
rect 24110 20738 24162 20750
rect 24558 20802 24610 20814
rect 27918 20802 27970 20814
rect 27122 20750 27134 20802
rect 27186 20750 27198 20802
rect 27682 20750 27694 20802
rect 27746 20750 27758 20802
rect 24558 20738 24610 20750
rect 27918 20738 27970 20750
rect 29262 20802 29314 20814
rect 29262 20738 29314 20750
rect 30270 20802 30322 20814
rect 30270 20738 30322 20750
rect 33854 20802 33906 20814
rect 33854 20738 33906 20750
rect 34190 20802 34242 20814
rect 34190 20738 34242 20750
rect 10110 20690 10162 20702
rect 7746 20638 7758 20690
rect 7810 20638 7822 20690
rect 10110 20626 10162 20638
rect 13470 20690 13522 20702
rect 13470 20626 13522 20638
rect 13582 20690 13634 20702
rect 22094 20690 22146 20702
rect 14578 20638 14590 20690
rect 14642 20638 14654 20690
rect 16482 20638 16494 20690
rect 16546 20638 16558 20690
rect 18386 20638 18398 20690
rect 18450 20638 18462 20690
rect 13582 20626 13634 20638
rect 22094 20626 22146 20638
rect 22654 20690 22706 20702
rect 22654 20626 22706 20638
rect 23774 20690 23826 20702
rect 23774 20626 23826 20638
rect 24446 20690 24498 20702
rect 24446 20626 24498 20638
rect 29598 20690 29650 20702
rect 29598 20626 29650 20638
rect 29822 20690 29874 20702
rect 29822 20626 29874 20638
rect 31614 20690 31666 20702
rect 31614 20626 31666 20638
rect 34526 20690 34578 20702
rect 34526 20626 34578 20638
rect 5070 20578 5122 20590
rect 5070 20514 5122 20526
rect 8094 20578 8146 20590
rect 8094 20514 8146 20526
rect 13806 20578 13858 20590
rect 13806 20514 13858 20526
rect 14478 20578 14530 20590
rect 14478 20514 14530 20526
rect 21310 20578 21362 20590
rect 21310 20514 21362 20526
rect 23438 20578 23490 20590
rect 23438 20514 23490 20526
rect 24670 20578 24722 20590
rect 24670 20514 24722 20526
rect 27806 20578 27858 20590
rect 27806 20514 27858 20526
rect 32286 20578 32338 20590
rect 32286 20514 32338 20526
rect 32398 20578 32450 20590
rect 32398 20514 32450 20526
rect 32958 20578 33010 20590
rect 32958 20514 33010 20526
rect 34190 20578 34242 20590
rect 34190 20514 34242 20526
rect 1344 20410 43568 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 43568 20410
rect 1344 20324 43568 20358
rect 12014 20242 12066 20254
rect 10434 20190 10446 20242
rect 10498 20190 10510 20242
rect 12014 20178 12066 20190
rect 14814 20242 14866 20254
rect 14814 20178 14866 20190
rect 15598 20242 15650 20254
rect 15598 20178 15650 20190
rect 29262 20242 29314 20254
rect 29262 20178 29314 20190
rect 30046 20242 30098 20254
rect 30046 20178 30098 20190
rect 30382 20242 30434 20254
rect 30382 20178 30434 20190
rect 31278 20242 31330 20254
rect 31278 20178 31330 20190
rect 23886 20130 23938 20142
rect 13234 20078 13246 20130
rect 13298 20078 13310 20130
rect 13906 20078 13918 20130
rect 13970 20078 13982 20130
rect 21410 20078 21422 20130
rect 21474 20078 21486 20130
rect 23886 20066 23938 20078
rect 24110 20130 24162 20142
rect 24110 20066 24162 20078
rect 28030 20130 28082 20142
rect 28030 20066 28082 20078
rect 29038 20130 29090 20142
rect 29038 20066 29090 20078
rect 30270 20130 30322 20142
rect 30270 20066 30322 20078
rect 30718 20130 30770 20142
rect 30718 20066 30770 20078
rect 32062 20130 32114 20142
rect 32062 20066 32114 20078
rect 9550 20018 9602 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 5954 19966 5966 20018
rect 6018 19966 6030 20018
rect 9550 19954 9602 19966
rect 10110 20018 10162 20030
rect 10110 19954 10162 19966
rect 11006 20018 11058 20030
rect 15262 20018 15314 20030
rect 16046 20018 16098 20030
rect 12562 19966 12574 20018
rect 12626 19966 12638 20018
rect 13122 19966 13134 20018
rect 13186 19966 13198 20018
rect 14242 19966 14254 20018
rect 14306 19966 14318 20018
rect 15698 19966 15710 20018
rect 15762 19966 15774 20018
rect 11006 19954 11058 19966
rect 15262 19954 15314 19966
rect 16046 19954 16098 19966
rect 16382 20018 16434 20030
rect 29710 20018 29762 20030
rect 22194 19966 22206 20018
rect 22258 19966 22270 20018
rect 23090 19966 23102 20018
rect 23154 19966 23166 20018
rect 29474 19966 29486 20018
rect 29538 19966 29550 20018
rect 16382 19954 16434 19966
rect 29710 19954 29762 19966
rect 31502 20018 31554 20030
rect 31502 19954 31554 19966
rect 31726 20018 31778 20030
rect 31726 19954 31778 19966
rect 32510 20018 32562 20030
rect 33170 19966 33182 20018
rect 33234 19966 33246 20018
rect 32510 19954 32562 19966
rect 1934 19906 1986 19918
rect 1934 19842 1986 19854
rect 6414 19906 6466 19918
rect 6414 19842 6466 19854
rect 16830 19906 16882 19918
rect 16830 19842 16882 19854
rect 17502 19906 17554 19918
rect 22766 19906 22818 19918
rect 19282 19854 19294 19906
rect 19346 19854 19358 19906
rect 17502 19842 17554 19854
rect 22766 19842 22818 19854
rect 24558 19906 24610 19918
rect 24558 19842 24610 19854
rect 25342 19906 25394 19918
rect 25342 19842 25394 19854
rect 28478 19906 28530 19918
rect 28478 19842 28530 19854
rect 29374 19906 29426 19918
rect 29374 19842 29426 19854
rect 31614 19906 31666 19918
rect 36542 19906 36594 19918
rect 33954 19854 33966 19906
rect 34018 19854 34030 19906
rect 36082 19854 36094 19906
rect 36146 19854 36158 19906
rect 31614 19842 31666 19854
rect 36542 19842 36594 19854
rect 10782 19794 10834 19806
rect 10782 19730 10834 19742
rect 15934 19794 15986 19806
rect 15934 19730 15986 19742
rect 23102 19794 23154 19806
rect 23102 19730 23154 19742
rect 23438 19794 23490 19806
rect 23438 19730 23490 19742
rect 23774 19794 23826 19806
rect 27906 19742 27918 19794
rect 27970 19791 27982 19794
rect 28354 19791 28366 19794
rect 27970 19745 28366 19791
rect 27970 19742 27982 19745
rect 28354 19742 28366 19745
rect 28418 19742 28430 19794
rect 23774 19730 23826 19742
rect 1344 19626 43568 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 43568 19626
rect 1344 19540 43568 19574
rect 16046 19458 16098 19470
rect 23102 19458 23154 19470
rect 21746 19406 21758 19458
rect 21810 19406 21822 19458
rect 16046 19394 16098 19406
rect 23102 19394 23154 19406
rect 34750 19458 34802 19470
rect 34750 19394 34802 19406
rect 35086 19458 35138 19470
rect 35086 19394 35138 19406
rect 35422 19458 35474 19470
rect 35422 19394 35474 19406
rect 1934 19346 1986 19358
rect 15038 19346 15090 19358
rect 20750 19346 20802 19358
rect 12226 19294 12238 19346
rect 12290 19294 12302 19346
rect 14018 19294 14030 19346
rect 14082 19294 14094 19346
rect 17042 19294 17054 19346
rect 17106 19294 17118 19346
rect 17378 19294 17390 19346
rect 17442 19294 17454 19346
rect 1934 19282 1986 19294
rect 15038 19282 15090 19294
rect 20750 19282 20802 19294
rect 24334 19346 24386 19358
rect 24334 19282 24386 19294
rect 28590 19346 28642 19358
rect 36430 19346 36482 19358
rect 35746 19294 35758 19346
rect 35810 19294 35822 19346
rect 36194 19294 36206 19346
rect 36258 19294 36270 19346
rect 28590 19282 28642 19294
rect 36430 19282 36482 19294
rect 7310 19234 7362 19246
rect 10558 19234 10610 19246
rect 3938 19182 3950 19234
rect 4002 19182 4014 19234
rect 5730 19182 5742 19234
rect 5794 19182 5806 19234
rect 6626 19182 6638 19234
rect 6690 19182 6702 19234
rect 6962 19182 6974 19234
rect 7026 19182 7038 19234
rect 10098 19182 10110 19234
rect 10162 19182 10174 19234
rect 7310 19170 7362 19182
rect 10558 19170 10610 19182
rect 11230 19234 11282 19246
rect 13582 19234 13634 19246
rect 11554 19182 11566 19234
rect 11618 19182 11630 19234
rect 12338 19182 12350 19234
rect 12402 19182 12414 19234
rect 11230 19170 11282 19182
rect 13582 19170 13634 19182
rect 13918 19234 13970 19246
rect 22318 19234 22370 19246
rect 16034 19182 16046 19234
rect 16098 19182 16110 19234
rect 20290 19182 20302 19234
rect 20354 19182 20366 19234
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 13918 19170 13970 19182
rect 22318 19170 22370 19182
rect 22654 19234 22706 19246
rect 23886 19234 23938 19246
rect 22866 19182 22878 19234
rect 22930 19182 22942 19234
rect 23314 19182 23326 19234
rect 23378 19182 23390 19234
rect 22654 19170 22706 19182
rect 23886 19170 23938 19182
rect 24782 19234 24834 19246
rect 37102 19234 37154 19246
rect 29138 19182 29150 19234
rect 29202 19182 29214 19234
rect 36082 19182 36094 19234
rect 36146 19182 36158 19234
rect 24782 19170 24834 19182
rect 37102 19170 37154 19182
rect 16382 19122 16434 19134
rect 5842 19070 5854 19122
rect 5906 19070 5918 19122
rect 12674 19070 12686 19122
rect 12738 19070 12750 19122
rect 14242 19070 14254 19122
rect 14306 19119 14318 19122
rect 14306 19073 14527 19119
rect 14306 19070 14318 19073
rect 4734 19010 4786 19022
rect 4734 18946 4786 18958
rect 13694 19010 13746 19022
rect 13694 18946 13746 18958
rect 14030 19010 14082 19022
rect 14481 19010 14527 19073
rect 16382 19058 16434 19070
rect 16718 19122 16770 19134
rect 23774 19122 23826 19134
rect 34862 19122 34914 19134
rect 19506 19070 19518 19122
rect 19570 19070 19582 19122
rect 22082 19070 22094 19122
rect 22146 19070 22158 19122
rect 32050 19070 32062 19122
rect 32114 19070 32126 19122
rect 16718 19058 16770 19070
rect 23774 19058 23826 19070
rect 34862 19058 34914 19070
rect 35646 19122 35698 19134
rect 35646 19058 35698 19070
rect 14590 19010 14642 19022
rect 14466 18958 14478 19010
rect 14530 18958 14542 19010
rect 14030 18946 14082 18958
rect 14590 18946 14642 18958
rect 15710 19010 15762 19022
rect 15710 18946 15762 18958
rect 16942 19010 16994 19022
rect 21858 18958 21870 19010
rect 21922 18958 21934 19010
rect 22978 18958 22990 19010
rect 23042 18958 23054 19010
rect 16942 18946 16994 18958
rect 1344 18842 43568 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 43568 18842
rect 1344 18756 43568 18790
rect 2718 18674 2770 18686
rect 10894 18674 10946 18686
rect 21534 18674 21586 18686
rect 22318 18674 22370 18686
rect 7634 18622 7646 18674
rect 7698 18622 7710 18674
rect 13010 18622 13022 18674
rect 13074 18622 13086 18674
rect 17938 18622 17950 18674
rect 18002 18622 18014 18674
rect 20626 18622 20638 18674
rect 20690 18622 20702 18674
rect 21970 18622 21982 18674
rect 22034 18622 22046 18674
rect 2718 18610 2770 18622
rect 10894 18610 10946 18622
rect 21534 18610 21586 18622
rect 22318 18610 22370 18622
rect 23102 18674 23154 18686
rect 23102 18610 23154 18622
rect 34526 18674 34578 18686
rect 38322 18622 38334 18674
rect 38386 18622 38398 18674
rect 34526 18610 34578 18622
rect 2046 18562 2098 18574
rect 21422 18562 21474 18574
rect 6290 18510 6302 18562
rect 6354 18510 6366 18562
rect 7858 18510 7870 18562
rect 7922 18510 7934 18562
rect 11442 18510 11454 18562
rect 11506 18510 11518 18562
rect 13346 18510 13358 18562
rect 13410 18510 13422 18562
rect 17490 18510 17502 18562
rect 17554 18510 17566 18562
rect 36082 18510 36094 18562
rect 36146 18510 36158 18562
rect 2046 18498 2098 18510
rect 21422 18498 21474 18510
rect 1710 18450 1762 18462
rect 1710 18386 1762 18398
rect 2382 18450 2434 18462
rect 2382 18386 2434 18398
rect 3614 18450 3666 18462
rect 9550 18450 9602 18462
rect 4498 18398 4510 18450
rect 4562 18398 4574 18450
rect 5506 18398 5518 18450
rect 5570 18398 5582 18450
rect 5730 18398 5742 18450
rect 5794 18398 5806 18450
rect 6850 18398 6862 18450
rect 6914 18398 6926 18450
rect 7186 18398 7198 18450
rect 7250 18398 7262 18450
rect 3614 18386 3666 18398
rect 9550 18386 9602 18398
rect 10110 18450 10162 18462
rect 12910 18450 12962 18462
rect 11666 18398 11678 18450
rect 11730 18398 11742 18450
rect 12338 18398 12350 18450
rect 12402 18398 12414 18450
rect 10110 18386 10162 18398
rect 12910 18386 12962 18398
rect 13694 18450 13746 18462
rect 13694 18386 13746 18398
rect 14254 18450 14306 18462
rect 19406 18450 19458 18462
rect 20974 18450 21026 18462
rect 17378 18398 17390 18450
rect 17442 18398 17454 18450
rect 18386 18398 18398 18450
rect 18450 18398 18462 18450
rect 18946 18398 18958 18450
rect 19010 18398 19022 18450
rect 19618 18398 19630 18450
rect 19682 18398 19694 18450
rect 14254 18386 14306 18398
rect 19406 18386 19458 18398
rect 20974 18386 21026 18398
rect 22766 18450 22818 18462
rect 22766 18386 22818 18398
rect 23550 18450 23602 18462
rect 34974 18450 35026 18462
rect 25330 18398 25342 18450
rect 25394 18398 25406 18450
rect 26002 18398 26014 18450
rect 26066 18398 26078 18450
rect 30818 18398 30830 18450
rect 30882 18398 30894 18450
rect 31490 18398 31502 18450
rect 31554 18398 31566 18450
rect 35410 18398 35422 18450
rect 35474 18398 35486 18450
rect 23550 18386 23602 18398
rect 34974 18386 35026 18398
rect 3166 18338 3218 18350
rect 3166 18274 3218 18286
rect 4174 18338 4226 18350
rect 4174 18274 4226 18286
rect 14702 18338 14754 18350
rect 14702 18274 14754 18286
rect 16606 18338 16658 18350
rect 16606 18274 16658 18286
rect 20302 18338 20354 18350
rect 20302 18274 20354 18286
rect 28142 18338 28194 18350
rect 32062 18338 32114 18350
rect 28690 18286 28702 18338
rect 28754 18286 28766 18338
rect 28142 18274 28194 18286
rect 32062 18274 32114 18286
rect 19294 18226 19346 18238
rect 5394 18174 5406 18226
rect 5458 18174 5470 18226
rect 14018 18174 14030 18226
rect 14082 18223 14094 18226
rect 14466 18223 14478 18226
rect 14082 18177 14478 18223
rect 14082 18174 14094 18177
rect 14466 18174 14478 18177
rect 14530 18223 14542 18226
rect 14690 18223 14702 18226
rect 14530 18177 14702 18223
rect 14530 18174 14542 18177
rect 14690 18174 14702 18177
rect 14754 18174 14766 18226
rect 19294 18162 19346 18174
rect 21646 18226 21698 18238
rect 21646 18162 21698 18174
rect 1344 18058 43568 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 43568 18058
rect 1344 17972 43568 18006
rect 17838 17890 17890 17902
rect 17838 17826 17890 17838
rect 3166 17778 3218 17790
rect 1922 17726 1934 17778
rect 1986 17726 1998 17778
rect 3166 17714 3218 17726
rect 3278 17778 3330 17790
rect 14142 17778 14194 17790
rect 9650 17726 9662 17778
rect 9714 17726 9726 17778
rect 3278 17714 3330 17726
rect 14142 17714 14194 17726
rect 19294 17778 19346 17790
rect 19294 17714 19346 17726
rect 21870 17778 21922 17790
rect 25566 17778 25618 17790
rect 22978 17726 22990 17778
rect 23042 17726 23054 17778
rect 25106 17726 25118 17778
rect 25170 17726 25182 17778
rect 21870 17714 21922 17726
rect 25566 17714 25618 17726
rect 28590 17778 28642 17790
rect 34190 17778 34242 17790
rect 33730 17726 33742 17778
rect 33794 17726 33806 17778
rect 28590 17714 28642 17726
rect 34190 17714 34242 17726
rect 17390 17666 17442 17678
rect 5058 17614 5070 17666
rect 5122 17614 5134 17666
rect 5842 17614 5854 17666
rect 5906 17614 5918 17666
rect 7858 17614 7870 17666
rect 7922 17614 7934 17666
rect 8306 17614 8318 17666
rect 8370 17614 8382 17666
rect 11442 17614 11454 17666
rect 11506 17614 11518 17666
rect 17390 17602 17442 17614
rect 17726 17666 17778 17678
rect 18510 17666 18562 17678
rect 17938 17614 17950 17666
rect 18002 17614 18014 17666
rect 22306 17614 22318 17666
rect 22370 17614 22382 17666
rect 30818 17614 30830 17666
rect 30882 17614 30894 17666
rect 17726 17602 17778 17614
rect 18510 17602 18562 17614
rect 2158 17554 2210 17566
rect 2158 17490 2210 17502
rect 4510 17554 4562 17566
rect 6402 17502 6414 17554
rect 6466 17502 6478 17554
rect 10098 17502 10110 17554
rect 10162 17502 10174 17554
rect 11666 17502 11678 17554
rect 11730 17502 11742 17554
rect 18834 17502 18846 17554
rect 18898 17502 18910 17554
rect 31602 17502 31614 17554
rect 31666 17502 31678 17554
rect 4510 17490 4562 17502
rect 5854 17442 5906 17454
rect 5854 17378 5906 17390
rect 13582 17442 13634 17454
rect 13582 17378 13634 17390
rect 16606 17442 16658 17454
rect 16606 17378 16658 17390
rect 18174 17442 18226 17454
rect 18174 17378 18226 17390
rect 19742 17442 19794 17454
rect 19742 17378 19794 17390
rect 1344 17274 43568 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 43568 17274
rect 1344 17188 43568 17222
rect 4062 17106 4114 17118
rect 3490 17054 3502 17106
rect 3554 17054 3566 17106
rect 4062 17042 4114 17054
rect 4286 17106 4338 17118
rect 4286 17042 4338 17054
rect 13694 17106 13746 17118
rect 13694 17042 13746 17054
rect 16158 17106 16210 17118
rect 16158 17042 16210 17054
rect 18734 17106 18786 17118
rect 18734 17042 18786 17054
rect 22206 17106 22258 17118
rect 22206 17042 22258 17054
rect 27358 17106 27410 17118
rect 27358 17042 27410 17054
rect 27582 17106 27634 17118
rect 27582 17042 27634 17054
rect 29262 17106 29314 17118
rect 29262 17042 29314 17054
rect 33294 17106 33346 17118
rect 33294 17042 33346 17054
rect 6078 16994 6130 17006
rect 7534 16994 7586 17006
rect 17950 16994 18002 17006
rect 6738 16942 6750 16994
rect 6802 16942 6814 16994
rect 13794 16942 13806 16994
rect 13858 16942 13870 16994
rect 15922 16942 15934 16994
rect 15986 16942 15998 16994
rect 6078 16930 6130 16942
rect 7534 16930 7586 16942
rect 17950 16930 18002 16942
rect 20974 16994 21026 17006
rect 20974 16930 21026 16942
rect 21870 16994 21922 17006
rect 27906 16942 27918 16994
rect 27970 16942 27982 16994
rect 21870 16930 21922 16942
rect 2046 16882 2098 16894
rect 2046 16818 2098 16830
rect 2606 16882 2658 16894
rect 2606 16818 2658 16830
rect 2942 16882 2994 16894
rect 2942 16818 2994 16830
rect 3838 16882 3890 16894
rect 3838 16818 3890 16830
rect 4510 16882 4562 16894
rect 6974 16882 7026 16894
rect 20414 16882 20466 16894
rect 29150 16882 29202 16894
rect 4834 16830 4846 16882
rect 4898 16830 4910 16882
rect 9874 16830 9886 16882
rect 9938 16830 9950 16882
rect 10098 16830 10110 16882
rect 10162 16830 10174 16882
rect 13010 16830 13022 16882
rect 13074 16830 13086 16882
rect 14130 16830 14142 16882
rect 14194 16830 14206 16882
rect 14914 16830 14926 16882
rect 14978 16830 14990 16882
rect 15138 16830 15150 16882
rect 15202 16830 15214 16882
rect 18162 16830 18174 16882
rect 18226 16830 18238 16882
rect 21634 16830 21646 16882
rect 21698 16830 21710 16882
rect 4510 16818 4562 16830
rect 6974 16818 7026 16830
rect 20414 16818 20466 16830
rect 29150 16818 29202 16830
rect 4622 16770 4674 16782
rect 16830 16770 16882 16782
rect 9650 16718 9662 16770
rect 9714 16718 9726 16770
rect 13346 16718 13358 16770
rect 13410 16718 13422 16770
rect 4622 16706 4674 16718
rect 16830 16706 16882 16718
rect 17614 16770 17666 16782
rect 33070 16770 33122 16782
rect 22642 16718 22654 16770
rect 22706 16718 22718 16770
rect 17614 16706 17666 16718
rect 33070 16706 33122 16718
rect 33182 16770 33234 16782
rect 33182 16706 33234 16718
rect 3166 16658 3218 16670
rect 10546 16606 10558 16658
rect 10610 16606 10622 16658
rect 3166 16594 3218 16606
rect 1344 16490 43568 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 43568 16490
rect 1344 16404 43568 16438
rect 4510 16210 4562 16222
rect 17390 16210 17442 16222
rect 2146 16158 2158 16210
rect 2210 16158 2222 16210
rect 8306 16158 8318 16210
rect 8370 16158 8382 16210
rect 11890 16158 11902 16210
rect 11954 16158 11966 16210
rect 15474 16158 15486 16210
rect 15538 16158 15550 16210
rect 4510 16146 4562 16158
rect 17390 16146 17442 16158
rect 17726 16210 17778 16222
rect 17726 16146 17778 16158
rect 18958 16210 19010 16222
rect 18958 16146 19010 16158
rect 22094 16210 22146 16222
rect 22094 16146 22146 16158
rect 28142 16210 28194 16222
rect 35646 16210 35698 16222
rect 32834 16158 32846 16210
rect 32898 16158 32910 16210
rect 35074 16158 35086 16210
rect 35138 16158 35150 16210
rect 28142 16146 28194 16158
rect 35646 16146 35698 16158
rect 3054 16098 3106 16110
rect 3054 16034 3106 16046
rect 3278 16098 3330 16110
rect 3278 16034 3330 16046
rect 3390 16098 3442 16110
rect 3390 16034 3442 16046
rect 4734 16098 4786 16110
rect 16158 16098 16210 16110
rect 17950 16098 18002 16110
rect 5618 16046 5630 16098
rect 5682 16046 5694 16098
rect 7634 16046 7646 16098
rect 7698 16046 7710 16098
rect 10882 16046 10894 16098
rect 10946 16046 10958 16098
rect 14130 16046 14142 16098
rect 14194 16046 14206 16098
rect 14914 16046 14926 16098
rect 14978 16046 14990 16098
rect 15138 16046 15150 16098
rect 15202 16046 15214 16098
rect 16818 16046 16830 16098
rect 16882 16046 16894 16098
rect 4734 16034 4786 16046
rect 16158 16034 16210 16046
rect 17950 16034 18002 16046
rect 29486 16098 29538 16110
rect 29486 16034 29538 16046
rect 29934 16098 29986 16110
rect 29934 16034 29986 16046
rect 30270 16098 30322 16110
rect 32050 16046 32062 16098
rect 32114 16046 32126 16098
rect 30270 16034 30322 16046
rect 2942 15986 2994 15998
rect 6750 15986 6802 15998
rect 5058 15934 5070 15986
rect 5122 15934 5134 15986
rect 2942 15922 2994 15934
rect 6750 15922 6802 15934
rect 8766 15986 8818 15998
rect 11454 15986 11506 15998
rect 19294 15986 19346 15998
rect 11106 15934 11118 15986
rect 11170 15934 11182 15986
rect 13906 15934 13918 15986
rect 13970 15934 13982 15986
rect 15922 15934 15934 15986
rect 15986 15934 15998 15986
rect 16594 15934 16606 15986
rect 16658 15934 16670 15986
rect 8766 15922 8818 15934
rect 11454 15922 11506 15934
rect 19294 15922 19346 15934
rect 19406 15986 19458 15998
rect 19406 15922 19458 15934
rect 29150 15986 29202 15998
rect 29150 15922 29202 15934
rect 29262 15986 29314 15998
rect 29262 15922 29314 15934
rect 29710 15986 29762 15998
rect 29710 15922 29762 15934
rect 2606 15874 2658 15886
rect 19630 15874 19682 15886
rect 18274 15822 18286 15874
rect 18338 15822 18350 15874
rect 2606 15810 2658 15822
rect 19630 15810 19682 15822
rect 26910 15874 26962 15886
rect 26910 15810 26962 15822
rect 29934 15874 29986 15886
rect 29934 15810 29986 15822
rect 1344 15706 43568 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 43568 15706
rect 1344 15620 43568 15654
rect 3390 15538 3442 15550
rect 8542 15538 8594 15550
rect 6290 15486 6302 15538
rect 6354 15486 6366 15538
rect 3390 15474 3442 15486
rect 8542 15474 8594 15486
rect 11454 15538 11506 15550
rect 11454 15474 11506 15486
rect 11678 15538 11730 15550
rect 11678 15474 11730 15486
rect 13134 15538 13186 15550
rect 17502 15538 17554 15550
rect 16258 15486 16270 15538
rect 16322 15486 16334 15538
rect 13134 15474 13186 15486
rect 17502 15474 17554 15486
rect 17726 15538 17778 15550
rect 17726 15474 17778 15486
rect 18510 15538 18562 15550
rect 18510 15474 18562 15486
rect 20190 15538 20242 15550
rect 20190 15474 20242 15486
rect 21534 15538 21586 15550
rect 21534 15474 21586 15486
rect 22878 15538 22930 15550
rect 22878 15474 22930 15486
rect 26350 15538 26402 15550
rect 26350 15474 26402 15486
rect 28926 15538 28978 15550
rect 32386 15486 32398 15538
rect 32450 15486 32462 15538
rect 28926 15474 28978 15486
rect 4622 15426 4674 15438
rect 4622 15362 4674 15374
rect 6638 15426 6690 15438
rect 18062 15426 18114 15438
rect 22094 15426 22146 15438
rect 28702 15426 28754 15438
rect 15586 15374 15598 15426
rect 15650 15374 15662 15426
rect 20514 15374 20526 15426
rect 20578 15374 20590 15426
rect 25666 15374 25678 15426
rect 25730 15374 25742 15426
rect 27570 15374 27582 15426
rect 27634 15374 27646 15426
rect 30146 15374 30158 15426
rect 30210 15374 30222 15426
rect 6638 15362 6690 15374
rect 18062 15362 18114 15374
rect 22094 15362 22146 15374
rect 28702 15362 28754 15374
rect 2382 15314 2434 15326
rect 1922 15262 1934 15314
rect 1986 15262 1998 15314
rect 2382 15250 2434 15262
rect 2830 15314 2882 15326
rect 6078 15314 6130 15326
rect 11230 15314 11282 15326
rect 3938 15262 3950 15314
rect 4002 15262 4014 15314
rect 9762 15262 9774 15314
rect 9826 15262 9838 15314
rect 2830 15250 2882 15262
rect 6078 15250 6130 15262
rect 11230 15250 11282 15262
rect 11342 15314 11394 15326
rect 11342 15250 11394 15262
rect 11566 15314 11618 15326
rect 11566 15250 11618 15262
rect 12462 15314 12514 15326
rect 12462 15250 12514 15262
rect 15934 15314 15986 15326
rect 15934 15250 15986 15262
rect 16606 15314 16658 15326
rect 16606 15250 16658 15262
rect 17390 15314 17442 15326
rect 17390 15250 17442 15262
rect 21646 15314 21698 15326
rect 26910 15314 26962 15326
rect 28590 15314 28642 15326
rect 22306 15262 22318 15314
rect 22370 15262 22382 15314
rect 25890 15262 25902 15314
rect 25954 15262 25966 15314
rect 27346 15262 27358 15314
rect 27410 15262 27422 15314
rect 29362 15262 29374 15314
rect 29426 15262 29438 15314
rect 21646 15250 21698 15262
rect 26910 15250 26962 15262
rect 28590 15250 28642 15262
rect 8766 15202 8818 15214
rect 12686 15202 12738 15214
rect 8418 15150 8430 15202
rect 8482 15150 8494 15202
rect 9986 15150 9998 15202
rect 10050 15150 10062 15202
rect 8766 15138 8818 15150
rect 12686 15138 12738 15150
rect 15038 15202 15090 15214
rect 15038 15138 15090 15150
rect 25342 15202 25394 15214
rect 27794 15150 27806 15202
rect 27858 15150 27870 15202
rect 25342 15138 25394 15150
rect 3054 15090 3106 15102
rect 21534 15090 21586 15102
rect 10210 15038 10222 15090
rect 10274 15038 10286 15090
rect 12114 15038 12126 15090
rect 12178 15038 12190 15090
rect 3054 15026 3106 15038
rect 21534 15026 21586 15038
rect 1344 14922 43568 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 43568 14922
rect 1344 14836 43568 14870
rect 14702 14754 14754 14766
rect 16146 14702 16158 14754
rect 16210 14702 16222 14754
rect 14702 14690 14754 14702
rect 2494 14642 2546 14654
rect 5070 14642 5122 14654
rect 3490 14590 3502 14642
rect 3554 14590 3566 14642
rect 2494 14578 2546 14590
rect 5070 14578 5122 14590
rect 7422 14642 7474 14654
rect 7422 14578 7474 14590
rect 10894 14642 10946 14654
rect 10894 14578 10946 14590
rect 24670 14642 24722 14654
rect 24670 14578 24722 14590
rect 25230 14642 25282 14654
rect 25230 14578 25282 14590
rect 29710 14642 29762 14654
rect 29710 14578 29762 14590
rect 13470 14530 13522 14542
rect 3154 14478 3166 14530
rect 3218 14478 3230 14530
rect 5618 14478 5630 14530
rect 5682 14478 5694 14530
rect 10434 14478 10446 14530
rect 10498 14478 10510 14530
rect 13470 14466 13522 14478
rect 13918 14530 13970 14542
rect 13918 14466 13970 14478
rect 14814 14530 14866 14542
rect 14814 14466 14866 14478
rect 15262 14530 15314 14542
rect 15262 14466 15314 14478
rect 15598 14530 15650 14542
rect 15598 14466 15650 14478
rect 15822 14530 15874 14542
rect 15822 14466 15874 14478
rect 16494 14530 16546 14542
rect 16494 14466 16546 14478
rect 17166 14530 17218 14542
rect 17166 14466 17218 14478
rect 21198 14530 21250 14542
rect 21198 14466 21250 14478
rect 21534 14530 21586 14542
rect 21534 14466 21586 14478
rect 22542 14530 22594 14542
rect 22542 14466 22594 14478
rect 22878 14530 22930 14542
rect 22878 14466 22930 14478
rect 23326 14530 23378 14542
rect 23326 14466 23378 14478
rect 24222 14530 24274 14542
rect 24222 14466 24274 14478
rect 26014 14530 26066 14542
rect 26014 14466 26066 14478
rect 26574 14530 26626 14542
rect 26574 14466 26626 14478
rect 6638 14418 6690 14430
rect 6638 14354 6690 14366
rect 11790 14418 11842 14430
rect 11790 14354 11842 14366
rect 11902 14418 11954 14430
rect 11902 14354 11954 14366
rect 14254 14418 14306 14430
rect 14254 14354 14306 14366
rect 14702 14418 14754 14430
rect 14702 14354 14754 14366
rect 16830 14418 16882 14430
rect 16830 14354 16882 14366
rect 17278 14418 17330 14430
rect 17278 14354 17330 14366
rect 21870 14418 21922 14430
rect 21870 14354 21922 14366
rect 23102 14418 23154 14430
rect 23102 14354 23154 14366
rect 23662 14418 23714 14430
rect 23662 14354 23714 14366
rect 23886 14418 23938 14430
rect 23886 14354 23938 14366
rect 26686 14418 26738 14430
rect 26686 14354 26738 14366
rect 26910 14418 26962 14430
rect 26910 14354 26962 14366
rect 27134 14418 27186 14430
rect 27134 14354 27186 14366
rect 27358 14418 27410 14430
rect 27358 14354 27410 14366
rect 27694 14418 27746 14430
rect 27694 14354 27746 14366
rect 27918 14418 27970 14430
rect 27918 14354 27970 14366
rect 28254 14418 28306 14430
rect 28254 14354 28306 14366
rect 1934 14306 1986 14318
rect 1934 14242 1986 14254
rect 4510 14306 4562 14318
rect 4510 14242 4562 14254
rect 7086 14306 7138 14318
rect 7086 14242 7138 14254
rect 9998 14306 10050 14318
rect 9998 14242 10050 14254
rect 11566 14306 11618 14318
rect 11566 14242 11618 14254
rect 12350 14306 12402 14318
rect 12350 14242 12402 14254
rect 17502 14306 17554 14318
rect 17502 14242 17554 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 22654 14306 22706 14318
rect 22654 14242 22706 14254
rect 23438 14306 23490 14318
rect 23438 14242 23490 14254
rect 24110 14306 24162 14318
rect 24110 14242 24162 14254
rect 25678 14306 25730 14318
rect 25678 14242 25730 14254
rect 26126 14306 26178 14318
rect 26126 14242 26178 14254
rect 26350 14306 26402 14318
rect 26350 14242 26402 14254
rect 27582 14306 27634 14318
rect 27582 14242 27634 14254
rect 28142 14306 28194 14318
rect 28142 14242 28194 14254
rect 29262 14306 29314 14318
rect 29262 14242 29314 14254
rect 1344 14138 43568 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 43568 14138
rect 1344 14052 43568 14086
rect 1710 13970 1762 13982
rect 1710 13906 1762 13918
rect 2718 13970 2770 13982
rect 2718 13906 2770 13918
rect 11902 13970 11954 13982
rect 11902 13906 11954 13918
rect 14590 13970 14642 13982
rect 42814 13970 42866 13982
rect 19058 13918 19070 13970
rect 19122 13918 19134 13970
rect 14590 13906 14642 13918
rect 42814 13906 42866 13918
rect 3614 13858 3666 13870
rect 7758 13858 7810 13870
rect 7410 13806 7422 13858
rect 7474 13806 7486 13858
rect 3614 13794 3666 13806
rect 7758 13794 7810 13806
rect 17726 13858 17778 13870
rect 17726 13794 17778 13806
rect 18062 13858 18114 13870
rect 22542 13858 22594 13870
rect 21298 13806 21310 13858
rect 21362 13806 21374 13858
rect 18062 13794 18114 13806
rect 22542 13794 22594 13806
rect 26014 13858 26066 13870
rect 26014 13794 26066 13806
rect 26350 13858 26402 13870
rect 26350 13794 26402 13806
rect 26462 13858 26514 13870
rect 27682 13806 27694 13858
rect 27746 13806 27758 13858
rect 26462 13794 26514 13806
rect 2270 13746 2322 13758
rect 2270 13682 2322 13694
rect 3054 13746 3106 13758
rect 11006 13746 11058 13758
rect 6402 13694 6414 13746
rect 6466 13694 6478 13746
rect 7074 13694 7086 13746
rect 7138 13694 7150 13746
rect 7522 13694 7534 13746
rect 7586 13694 7598 13746
rect 3054 13682 3106 13694
rect 11006 13682 11058 13694
rect 18622 13746 18674 13758
rect 26686 13746 26738 13758
rect 43150 13746 43202 13758
rect 22082 13694 22094 13746
rect 22146 13694 22158 13746
rect 27010 13694 27022 13746
rect 27074 13694 27086 13746
rect 18622 13682 18674 13694
rect 26686 13682 26738 13694
rect 43150 13682 43202 13694
rect 3950 13634 4002 13646
rect 15262 13634 15314 13646
rect 4162 13582 4174 13634
rect 4226 13582 4238 13634
rect 11218 13582 11230 13634
rect 11282 13582 11294 13634
rect 3950 13570 4002 13582
rect 15262 13570 15314 13582
rect 16606 13634 16658 13646
rect 16606 13570 16658 13582
rect 29822 13634 29874 13646
rect 29822 13570 29874 13582
rect 42590 13634 42642 13646
rect 42590 13570 42642 13582
rect 10770 13470 10782 13522
rect 10834 13470 10846 13522
rect 1344 13354 43568 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 43568 13354
rect 1344 13268 43568 13302
rect 17390 13186 17442 13198
rect 19730 13183 19742 13186
rect 17390 13122 17442 13134
rect 19297 13137 19742 13183
rect 3166 13074 3218 13086
rect 5854 13074 5906 13086
rect 2146 13022 2158 13074
rect 2210 13022 2222 13074
rect 3826 13022 3838 13074
rect 3890 13022 3902 13074
rect 3166 13010 3218 13022
rect 5854 13010 5906 13022
rect 6638 13074 6690 13086
rect 19297 13074 19343 13137
rect 19730 13134 19742 13137
rect 19794 13134 19806 13186
rect 19742 13074 19794 13086
rect 14130 13022 14142 13074
rect 14194 13022 14206 13074
rect 17714 13022 17726 13074
rect 17778 13022 17790 13074
rect 18498 13022 18510 13074
rect 18562 13022 18574 13074
rect 19282 13022 19294 13074
rect 19346 13022 19358 13074
rect 6638 13010 6690 13022
rect 19742 13010 19794 13022
rect 20750 13074 20802 13086
rect 25454 13074 25506 13086
rect 21746 13022 21758 13074
rect 21810 13022 21822 13074
rect 23314 13022 23326 13074
rect 23378 13022 23390 13074
rect 20750 13010 20802 13022
rect 25454 13010 25506 13022
rect 18846 12962 18898 12974
rect 1810 12910 1822 12962
rect 1874 12910 1886 12962
rect 2706 12910 2718 12962
rect 2770 12910 2782 12962
rect 14242 12910 14254 12962
rect 14306 12910 14318 12962
rect 18846 12898 18898 12910
rect 21310 12962 21362 12974
rect 27246 12962 27298 12974
rect 22642 12910 22654 12962
rect 22706 12910 22718 12962
rect 21310 12898 21362 12910
rect 27246 12898 27298 12910
rect 27470 12962 27522 12974
rect 27470 12898 27522 12910
rect 27806 12962 27858 12974
rect 27806 12898 27858 12910
rect 3502 12850 3554 12862
rect 3502 12786 3554 12798
rect 13694 12850 13746 12862
rect 13694 12786 13746 12798
rect 15038 12850 15090 12862
rect 15038 12786 15090 12798
rect 17614 12850 17666 12862
rect 17614 12786 17666 12798
rect 19182 12850 19234 12862
rect 19182 12786 19234 12798
rect 7086 12738 7138 12750
rect 7086 12674 7138 12686
rect 10334 12738 10386 12750
rect 10334 12674 10386 12686
rect 17054 12738 17106 12750
rect 17054 12674 17106 12686
rect 27470 12738 27522 12750
rect 27470 12674 27522 12686
rect 1344 12570 43568 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 43568 12570
rect 1344 12484 43568 12518
rect 2718 12402 2770 12414
rect 2718 12338 2770 12350
rect 4398 12402 4450 12414
rect 4398 12338 4450 12350
rect 5406 12402 5458 12414
rect 5406 12338 5458 12350
rect 5742 12402 5794 12414
rect 5742 12338 5794 12350
rect 6302 12402 6354 12414
rect 6302 12338 6354 12350
rect 7086 12402 7138 12414
rect 7086 12338 7138 12350
rect 7758 12402 7810 12414
rect 7758 12338 7810 12350
rect 10334 12402 10386 12414
rect 10334 12338 10386 12350
rect 10558 12402 10610 12414
rect 10558 12338 10610 12350
rect 11230 12402 11282 12414
rect 11230 12338 11282 12350
rect 14702 12402 14754 12414
rect 14702 12338 14754 12350
rect 18622 12402 18674 12414
rect 18622 12338 18674 12350
rect 26350 12402 26402 12414
rect 26350 12338 26402 12350
rect 5854 12290 5906 12302
rect 5854 12226 5906 12238
rect 6190 12290 6242 12302
rect 6190 12226 6242 12238
rect 8878 12290 8930 12302
rect 8878 12226 8930 12238
rect 9886 12290 9938 12302
rect 9886 12226 9938 12238
rect 16718 12290 16770 12302
rect 29362 12238 29374 12290
rect 29426 12238 29438 12290
rect 16718 12226 16770 12238
rect 1710 12178 1762 12190
rect 1710 12114 1762 12126
rect 2270 12178 2322 12190
rect 2270 12114 2322 12126
rect 5518 12178 5570 12190
rect 5518 12114 5570 12126
rect 7198 12178 7250 12190
rect 7198 12114 7250 12126
rect 8766 12178 8818 12190
rect 8766 12114 8818 12126
rect 9102 12178 9154 12190
rect 9102 12114 9154 12126
rect 9438 12178 9490 12190
rect 9438 12114 9490 12126
rect 10110 12178 10162 12190
rect 10110 12114 10162 12126
rect 10670 12178 10722 12190
rect 10670 12114 10722 12126
rect 13694 12178 13746 12190
rect 16830 12178 16882 12190
rect 17726 12178 17778 12190
rect 13906 12126 13918 12178
rect 13970 12126 13982 12178
rect 17602 12126 17614 12178
rect 17666 12126 17678 12178
rect 13694 12114 13746 12126
rect 16830 12114 16882 12126
rect 17726 12114 17778 12126
rect 17838 12178 17890 12190
rect 17838 12114 17890 12126
rect 18174 12178 18226 12190
rect 27122 12126 27134 12178
rect 27186 12126 27198 12178
rect 18174 12114 18226 12126
rect 3166 12066 3218 12078
rect 3166 12002 3218 12014
rect 4958 12066 5010 12078
rect 4958 12002 5010 12014
rect 9662 12066 9714 12078
rect 9662 12002 9714 12014
rect 18062 12066 18114 12078
rect 18062 12002 18114 12014
rect 6302 11954 6354 11966
rect 6302 11890 6354 11902
rect 7086 11954 7138 11966
rect 13570 11902 13582 11954
rect 13634 11902 13646 11954
rect 7086 11890 7138 11902
rect 1344 11786 43568 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 43568 11786
rect 1344 11700 43568 11734
rect 1822 11506 1874 11518
rect 5058 11454 5070 11506
rect 5122 11454 5134 11506
rect 6738 11454 6750 11506
rect 6802 11454 6814 11506
rect 8306 11454 8318 11506
rect 8370 11454 8382 11506
rect 10434 11454 10446 11506
rect 10498 11454 10510 11506
rect 1822 11442 1874 11454
rect 5630 11394 5682 11406
rect 2258 11342 2270 11394
rect 2322 11342 2334 11394
rect 5630 11330 5682 11342
rect 6078 11394 6130 11406
rect 11230 11394 11282 11406
rect 7074 11342 7086 11394
rect 7138 11342 7150 11394
rect 7522 11342 7534 11394
rect 7586 11342 7598 11394
rect 11666 11342 11678 11394
rect 11730 11342 11742 11394
rect 18722 11342 18734 11394
rect 18786 11342 18798 11394
rect 6078 11330 6130 11342
rect 11230 11330 11282 11342
rect 6302 11282 6354 11294
rect 12238 11282 12290 11294
rect 2930 11230 2942 11282
rect 2994 11230 3006 11282
rect 10882 11230 10894 11282
rect 10946 11230 10958 11282
rect 11890 11230 11902 11282
rect 11954 11230 11966 11282
rect 6302 11218 6354 11230
rect 12238 11218 12290 11230
rect 12350 11282 12402 11294
rect 22318 11282 22370 11294
rect 13682 11230 13694 11282
rect 13746 11230 13758 11282
rect 12350 11218 12402 11230
rect 22318 11218 22370 11230
rect 22430 11282 22482 11294
rect 22430 11218 22482 11230
rect 22990 11282 23042 11294
rect 22990 11218 23042 11230
rect 5854 11170 5906 11182
rect 5854 11106 5906 11118
rect 12574 11170 12626 11182
rect 12574 11106 12626 11118
rect 19182 11170 19234 11182
rect 19182 11106 19234 11118
rect 22654 11170 22706 11182
rect 22654 11106 22706 11118
rect 1344 11002 43568 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 43568 11002
rect 1344 10916 43568 10950
rect 5518 10834 5570 10846
rect 5518 10770 5570 10782
rect 5742 10834 5794 10846
rect 5742 10770 5794 10782
rect 6302 10834 6354 10846
rect 6302 10770 6354 10782
rect 7198 10834 7250 10846
rect 7198 10770 7250 10782
rect 7758 10834 7810 10846
rect 7758 10770 7810 10782
rect 10670 10834 10722 10846
rect 10670 10770 10722 10782
rect 14478 10834 14530 10846
rect 14478 10770 14530 10782
rect 15374 10834 15426 10846
rect 22206 10834 22258 10846
rect 17378 10782 17390 10834
rect 17442 10782 17454 10834
rect 15374 10770 15426 10782
rect 22206 10770 22258 10782
rect 23998 10834 24050 10846
rect 30146 10782 30158 10834
rect 30210 10782 30222 10834
rect 23998 10770 24050 10782
rect 5854 10722 5906 10734
rect 2930 10670 2942 10722
rect 2994 10670 3006 10722
rect 5854 10658 5906 10670
rect 7310 10722 7362 10734
rect 7310 10658 7362 10670
rect 15262 10722 15314 10734
rect 21646 10722 21698 10734
rect 19730 10670 19742 10722
rect 19794 10670 19806 10722
rect 15262 10658 15314 10670
rect 21646 10658 21698 10670
rect 22094 10722 22146 10734
rect 27906 10670 27918 10722
rect 27970 10670 27982 10722
rect 22094 10658 22146 10670
rect 6190 10610 6242 10622
rect 2258 10558 2270 10610
rect 2322 10558 2334 10610
rect 6190 10546 6242 10558
rect 6526 10610 6578 10622
rect 6526 10546 6578 10558
rect 6750 10610 6802 10622
rect 6750 10546 6802 10558
rect 6974 10610 7026 10622
rect 15598 10610 15650 10622
rect 11106 10558 11118 10610
rect 11170 10558 11182 10610
rect 6974 10546 7026 10558
rect 15598 10546 15650 10558
rect 15822 10610 15874 10622
rect 15822 10546 15874 10558
rect 16382 10610 16434 10622
rect 19406 10610 19458 10622
rect 17602 10558 17614 10610
rect 17666 10558 17678 10610
rect 16382 10546 16434 10558
rect 19406 10546 19458 10558
rect 21534 10610 21586 10622
rect 21534 10546 21586 10558
rect 21870 10610 21922 10622
rect 21870 10546 21922 10558
rect 22878 10610 22930 10622
rect 22878 10546 22930 10558
rect 23102 10610 23154 10622
rect 23102 10546 23154 10558
rect 23438 10610 23490 10622
rect 27234 10558 27246 10610
rect 27298 10558 27310 10610
rect 23438 10546 23490 10558
rect 1822 10498 1874 10510
rect 15038 10498 15090 10510
rect 5058 10446 5070 10498
rect 5122 10446 5134 10498
rect 11890 10446 11902 10498
rect 11954 10446 11966 10498
rect 14018 10446 14030 10498
rect 14082 10446 14094 10498
rect 1822 10434 1874 10446
rect 15038 10434 15090 10446
rect 20302 10498 20354 10510
rect 20302 10434 20354 10446
rect 20750 10498 20802 10510
rect 20750 10434 20802 10446
rect 21198 10498 21250 10510
rect 21198 10434 21250 10446
rect 22990 10498 23042 10510
rect 22990 10434 23042 10446
rect 22206 10386 22258 10398
rect 20290 10334 20302 10386
rect 20354 10383 20366 10386
rect 21298 10383 21310 10386
rect 20354 10337 21310 10383
rect 20354 10334 20366 10337
rect 21298 10334 21310 10337
rect 21362 10334 21374 10386
rect 22206 10322 22258 10334
rect 1344 10218 43568 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 43568 10218
rect 1344 10132 43568 10166
rect 12798 10050 12850 10062
rect 12798 9986 12850 9998
rect 2270 9938 2322 9950
rect 2270 9874 2322 9886
rect 5070 9938 5122 9950
rect 5070 9874 5122 9886
rect 5854 9938 5906 9950
rect 5854 9874 5906 9886
rect 6974 9938 7026 9950
rect 6974 9874 7026 9886
rect 7422 9938 7474 9950
rect 7422 9874 7474 9886
rect 12238 9938 12290 9950
rect 12238 9874 12290 9886
rect 13582 9938 13634 9950
rect 27918 9938 27970 9950
rect 15138 9886 15150 9938
rect 15202 9886 15214 9938
rect 15922 9886 15934 9938
rect 15986 9886 15998 9938
rect 18050 9886 18062 9938
rect 18114 9886 18126 9938
rect 26114 9886 26126 9938
rect 26178 9886 26190 9938
rect 13582 9874 13634 9886
rect 27918 9874 27970 9886
rect 30718 9938 30770 9950
rect 30718 9874 30770 9886
rect 6190 9826 6242 9838
rect 6190 9762 6242 9774
rect 6526 9826 6578 9838
rect 6526 9762 6578 9774
rect 11454 9826 11506 9838
rect 11454 9762 11506 9774
rect 12126 9826 12178 9838
rect 12126 9762 12178 9774
rect 12462 9826 12514 9838
rect 12462 9762 12514 9774
rect 12686 9826 12738 9838
rect 20526 9826 20578 9838
rect 18722 9774 18734 9826
rect 18786 9774 18798 9826
rect 12686 9762 12738 9774
rect 20526 9762 20578 9774
rect 22094 9826 22146 9838
rect 22094 9762 22146 9774
rect 22542 9826 22594 9838
rect 29262 9826 29314 9838
rect 23314 9774 23326 9826
rect 23378 9774 23390 9826
rect 22542 9762 22594 9774
rect 29262 9762 29314 9774
rect 1710 9714 1762 9726
rect 1710 9650 1762 9662
rect 11790 9714 11842 9726
rect 11790 9650 11842 9662
rect 21422 9714 21474 9726
rect 21870 9714 21922 9726
rect 21422 9650 21474 9662
rect 21758 9658 21810 9670
rect 6414 9602 6466 9614
rect 12798 9602 12850 9614
rect 11106 9550 11118 9602
rect 11170 9550 11182 9602
rect 6414 9538 6466 9550
rect 12798 9538 12850 9550
rect 14702 9602 14754 9614
rect 14702 9538 14754 9550
rect 19742 9602 19794 9614
rect 19742 9538 19794 9550
rect 20190 9602 20242 9614
rect 20190 9538 20242 9550
rect 20638 9602 20690 9614
rect 20638 9538 20690 9550
rect 20862 9602 20914 9614
rect 21870 9650 21922 9662
rect 22318 9714 22370 9726
rect 22318 9650 22370 9662
rect 22766 9714 22818 9726
rect 22766 9650 22818 9662
rect 22878 9714 22930 9726
rect 28142 9714 28194 9726
rect 23986 9662 23998 9714
rect 24050 9662 24062 9714
rect 22878 9650 22930 9662
rect 28142 9650 28194 9662
rect 28254 9714 28306 9726
rect 28254 9650 28306 9662
rect 29598 9714 29650 9726
rect 29598 9650 29650 9662
rect 29710 9714 29762 9726
rect 29710 9650 29762 9662
rect 21758 9594 21810 9606
rect 28478 9602 28530 9614
rect 20862 9538 20914 9550
rect 28478 9538 28530 9550
rect 29934 9602 29986 9614
rect 29934 9538 29986 9550
rect 30270 9602 30322 9614
rect 30270 9538 30322 9550
rect 1344 9434 43568 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 43568 9434
rect 1344 9348 43568 9382
rect 2046 9266 2098 9278
rect 2046 9202 2098 9214
rect 6078 9266 6130 9278
rect 6078 9202 6130 9214
rect 15374 9266 15426 9278
rect 15374 9202 15426 9214
rect 16158 9266 16210 9278
rect 16158 9202 16210 9214
rect 23998 9266 24050 9278
rect 23998 9202 24050 9214
rect 10558 9154 10610 9166
rect 10558 9090 10610 9102
rect 10670 9154 10722 9166
rect 15822 9154 15874 9166
rect 11218 9102 11230 9154
rect 11282 9102 11294 9154
rect 10670 9090 10722 9102
rect 15822 9090 15874 9102
rect 16718 9154 16770 9166
rect 22990 9154 23042 9166
rect 18722 9102 18734 9154
rect 18786 9102 18798 9154
rect 29250 9102 29262 9154
rect 29314 9102 29326 9154
rect 16718 9090 16770 9102
rect 22990 9090 23042 9102
rect 1710 9042 1762 9054
rect 1710 8978 1762 8990
rect 9550 9042 9602 9054
rect 10334 9042 10386 9054
rect 16270 9042 16322 9054
rect 9986 8990 9998 9042
rect 10050 8990 10062 9042
rect 11442 8990 11454 9042
rect 11506 8990 11518 9042
rect 9550 8978 9602 8990
rect 10334 8978 10386 8990
rect 16270 8978 16322 8990
rect 16606 9042 16658 9054
rect 16606 8978 16658 8990
rect 16942 9042 16994 9054
rect 23214 9042 23266 9054
rect 22642 8990 22654 9042
rect 22706 8990 22718 9042
rect 16942 8978 16994 8990
rect 23214 8978 23266 8990
rect 23438 9042 23490 9054
rect 25330 8990 25342 9042
rect 25394 8990 25406 9042
rect 28578 8990 28590 9042
rect 28642 8990 28654 9042
rect 23438 8978 23490 8990
rect 2494 8930 2546 8942
rect 2494 8866 2546 8878
rect 12014 8930 12066 8942
rect 12014 8866 12066 8878
rect 23102 8930 23154 8942
rect 26002 8878 26014 8930
rect 26066 8878 26078 8930
rect 28130 8878 28142 8930
rect 28194 8878 28206 8930
rect 31378 8878 31390 8930
rect 31442 8878 31454 8930
rect 23102 8866 23154 8878
rect 16158 8818 16210 8830
rect 16158 8754 16210 8766
rect 1344 8650 43568 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 43568 8650
rect 1344 8564 43568 8598
rect 15822 8370 15874 8382
rect 15822 8306 15874 8318
rect 16270 8370 16322 8382
rect 16270 8306 16322 8318
rect 23550 8370 23602 8382
rect 23550 8306 23602 8318
rect 9998 8258 10050 8270
rect 9998 8194 10050 8206
rect 11566 8258 11618 8270
rect 11566 8194 11618 8206
rect 12910 8258 12962 8270
rect 12910 8194 12962 8206
rect 13470 8258 13522 8270
rect 13470 8194 13522 8206
rect 17390 8258 17442 8270
rect 17390 8194 17442 8206
rect 17838 8258 17890 8270
rect 19294 8258 19346 8270
rect 18498 8206 18510 8258
rect 18562 8206 18574 8258
rect 17838 8194 17890 8206
rect 19294 8194 19346 8206
rect 19854 8258 19906 8270
rect 19854 8194 19906 8206
rect 20190 8258 20242 8270
rect 20190 8194 20242 8206
rect 21310 8258 21362 8270
rect 21310 8194 21362 8206
rect 21758 8258 21810 8270
rect 21758 8194 21810 8206
rect 21870 8258 21922 8270
rect 21870 8194 21922 8206
rect 22318 8258 22370 8270
rect 22318 8194 22370 8206
rect 22654 8258 22706 8270
rect 22654 8194 22706 8206
rect 23214 8258 23266 8270
rect 23214 8194 23266 8206
rect 9774 8146 9826 8158
rect 9774 8082 9826 8094
rect 10334 8146 10386 8158
rect 10334 8082 10386 8094
rect 10670 8146 10722 8158
rect 10670 8082 10722 8094
rect 12350 8146 12402 8158
rect 12350 8082 12402 8094
rect 12798 8146 12850 8158
rect 12798 8082 12850 8094
rect 16606 8146 16658 8158
rect 16606 8082 16658 8094
rect 16718 8146 16770 8158
rect 16718 8082 16770 8094
rect 17166 8146 17218 8158
rect 19182 8146 19234 8158
rect 18722 8094 18734 8146
rect 18786 8094 18798 8146
rect 17166 8082 17218 8094
rect 19182 8082 19234 8094
rect 20414 8146 20466 8158
rect 20414 8082 20466 8094
rect 20750 8146 20802 8158
rect 20750 8082 20802 8094
rect 22430 8146 22482 8158
rect 22430 8082 22482 8094
rect 22878 8146 22930 8158
rect 22878 8082 22930 8094
rect 22990 8146 23042 8158
rect 22990 8082 23042 8094
rect 9886 8034 9938 8046
rect 9886 7970 9938 7982
rect 11006 8034 11058 8046
rect 11006 7970 11058 7982
rect 11230 8034 11282 8046
rect 11230 7970 11282 7982
rect 11454 8034 11506 8046
rect 11454 7970 11506 7982
rect 12574 8034 12626 8046
rect 12574 7970 12626 7982
rect 13582 8034 13634 8046
rect 13582 7970 13634 7982
rect 13806 8034 13858 8046
rect 13806 7970 13858 7982
rect 14142 8034 14194 8046
rect 14142 7970 14194 7982
rect 16942 8034 16994 8046
rect 16942 7970 16994 7982
rect 17614 8034 17666 8046
rect 17614 7970 17666 7982
rect 18958 8034 19010 8046
rect 18958 7970 19010 7982
rect 19966 8034 20018 8046
rect 19966 7970 20018 7982
rect 21534 8034 21586 8046
rect 21534 7970 21586 7982
rect 1344 7866 43568 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 43568 7866
rect 1344 7780 43568 7814
rect 2046 7698 2098 7710
rect 2046 7634 2098 7646
rect 10222 7698 10274 7710
rect 10222 7634 10274 7646
rect 10446 7698 10498 7710
rect 10446 7634 10498 7646
rect 13022 7698 13074 7710
rect 13022 7634 13074 7646
rect 15374 7698 15426 7710
rect 15374 7634 15426 7646
rect 15822 7698 15874 7710
rect 15822 7634 15874 7646
rect 19070 7698 19122 7710
rect 19070 7634 19122 7646
rect 19294 7698 19346 7710
rect 19294 7634 19346 7646
rect 20302 7698 20354 7710
rect 20302 7634 20354 7646
rect 21422 7698 21474 7710
rect 21758 7698 21810 7710
rect 21422 7634 21474 7646
rect 21646 7642 21698 7654
rect 10558 7586 10610 7598
rect 10558 7522 10610 7534
rect 12014 7586 12066 7598
rect 12014 7522 12066 7534
rect 12910 7586 12962 7598
rect 12910 7522 12962 7534
rect 15934 7586 15986 7598
rect 15934 7522 15986 7534
rect 17390 7586 17442 7598
rect 17390 7522 17442 7534
rect 17726 7586 17778 7598
rect 17726 7522 17778 7534
rect 18062 7586 18114 7598
rect 18062 7522 18114 7534
rect 18622 7586 18674 7598
rect 18622 7522 18674 7534
rect 19966 7586 20018 7598
rect 19966 7522 20018 7534
rect 20638 7586 20690 7598
rect 21758 7634 21810 7646
rect 21982 7698 22034 7710
rect 21982 7634 22034 7646
rect 22654 7698 22706 7710
rect 22654 7634 22706 7646
rect 22990 7698 23042 7710
rect 22990 7634 23042 7646
rect 21646 7578 21698 7590
rect 20638 7522 20690 7534
rect 1710 7474 1762 7486
rect 1710 7410 1762 7422
rect 12350 7474 12402 7486
rect 12350 7410 12402 7422
rect 12686 7474 12738 7486
rect 12686 7410 12738 7422
rect 16158 7474 16210 7486
rect 16158 7410 16210 7422
rect 16494 7474 16546 7486
rect 16494 7410 16546 7422
rect 16830 7474 16882 7486
rect 16830 7410 16882 7422
rect 18398 7474 18450 7486
rect 18398 7410 18450 7422
rect 18958 7474 19010 7486
rect 18958 7410 19010 7422
rect 2494 7362 2546 7374
rect 2494 7298 2546 7310
rect 11006 7362 11058 7374
rect 11006 7298 11058 7310
rect 12462 7362 12514 7374
rect 12462 7298 12514 7310
rect 16382 7362 16434 7374
rect 16382 7298 16434 7310
rect 18510 7362 18562 7374
rect 18510 7298 18562 7310
rect 13022 7250 13074 7262
rect 13022 7186 13074 7198
rect 15822 7250 15874 7262
rect 15822 7186 15874 7198
rect 1344 7082 43568 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 43568 7082
rect 1344 6996 43568 7030
rect 19630 6802 19682 6814
rect 9986 6750 9998 6802
rect 10050 6750 10062 6802
rect 15810 6750 15822 6802
rect 15874 6750 15886 6802
rect 17938 6750 17950 6802
rect 18002 6750 18014 6802
rect 19630 6738 19682 6750
rect 19966 6802 20018 6814
rect 19966 6738 20018 6750
rect 10334 6690 10386 6702
rect 7074 6638 7086 6690
rect 7138 6638 7150 6690
rect 7858 6638 7870 6690
rect 7922 6638 7934 6690
rect 10334 6626 10386 6638
rect 10670 6690 10722 6702
rect 10670 6626 10722 6638
rect 11454 6690 11506 6702
rect 11454 6626 11506 6638
rect 11902 6690 11954 6702
rect 11902 6626 11954 6638
rect 12686 6690 12738 6702
rect 12686 6626 12738 6638
rect 13022 6690 13074 6702
rect 13022 6626 13074 6638
rect 13470 6690 13522 6702
rect 13470 6626 13522 6638
rect 13806 6690 13858 6702
rect 13806 6626 13858 6638
rect 14142 6690 14194 6702
rect 15138 6638 15150 6690
rect 15202 6638 15214 6690
rect 14142 6626 14194 6638
rect 10894 6578 10946 6590
rect 10894 6514 10946 6526
rect 11118 6578 11170 6590
rect 11118 6514 11170 6526
rect 12798 6578 12850 6590
rect 12798 6514 12850 6526
rect 10670 6466 10722 6478
rect 10670 6402 10722 6414
rect 11342 6466 11394 6478
rect 11342 6402 11394 6414
rect 13806 6466 13858 6478
rect 13806 6402 13858 6414
rect 18846 6466 18898 6478
rect 18846 6402 18898 6414
rect 1344 6298 43568 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 43568 6298
rect 1344 6212 43568 6246
rect 10222 6130 10274 6142
rect 10222 6066 10274 6078
rect 14254 6130 14306 6142
rect 24322 6078 24334 6130
rect 24386 6078 24398 6130
rect 14254 6066 14306 6078
rect 2034 5966 2046 6018
rect 2098 5966 2110 6018
rect 11666 5966 11678 6018
rect 11730 5966 11742 6018
rect 22082 5966 22094 6018
rect 22146 5966 22158 6018
rect 1710 5906 1762 5918
rect 10882 5854 10894 5906
rect 10946 5854 10958 5906
rect 17490 5854 17502 5906
rect 17554 5854 17566 5906
rect 21298 5854 21310 5906
rect 21362 5854 21374 5906
rect 1710 5842 1762 5854
rect 2494 5794 2546 5806
rect 13794 5742 13806 5794
rect 13858 5742 13870 5794
rect 2494 5730 2546 5742
rect 18398 5682 18450 5694
rect 18398 5618 18450 5630
rect 1344 5514 43568 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 43568 5514
rect 1344 5428 43568 5462
rect 11902 5234 11954 5246
rect 8866 5182 8878 5234
rect 8930 5182 8942 5234
rect 10994 5182 11006 5234
rect 11058 5182 11070 5234
rect 11902 5170 11954 5182
rect 12686 5234 12738 5246
rect 13458 5182 13470 5234
rect 13522 5182 13534 5234
rect 15586 5182 15598 5234
rect 15650 5182 15662 5234
rect 18610 5182 18622 5234
rect 18674 5182 18686 5234
rect 20738 5182 20750 5234
rect 20802 5182 20814 5234
rect 12686 5170 12738 5182
rect 1710 5122 1762 5134
rect 1710 5058 1762 5070
rect 2494 5122 2546 5134
rect 11790 5122 11842 5134
rect 42590 5122 42642 5134
rect 8082 5070 8094 5122
rect 8146 5070 8158 5122
rect 16370 5070 16382 5122
rect 16434 5070 16446 5122
rect 17826 5070 17838 5122
rect 17890 5070 17902 5122
rect 2494 5058 2546 5070
rect 11790 5058 11842 5070
rect 42590 5058 42642 5070
rect 43150 5122 43202 5134
rect 43150 5058 43202 5070
rect 2046 5010 2098 5022
rect 2046 4946 2098 4958
rect 12126 5010 12178 5022
rect 42802 4958 42814 5010
rect 42866 4958 42878 5010
rect 12126 4946 12178 4958
rect 1344 4730 43568 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 43568 4730
rect 1344 4644 43568 4678
rect 10558 4562 10610 4574
rect 10558 4498 10610 4510
rect 23886 4562 23938 4574
rect 23886 4498 23938 4510
rect 36654 4562 36706 4574
rect 36654 4498 36706 4510
rect 18162 4398 18174 4450
rect 18226 4398 18238 4450
rect 10110 4338 10162 4350
rect 42366 4338 42418 4350
rect 1810 4286 1822 4338
rect 1874 4286 1886 4338
rect 6066 4286 6078 4338
rect 6130 4286 6142 4338
rect 6402 4286 6414 4338
rect 6466 4286 6478 4338
rect 12898 4286 12910 4338
rect 12962 4286 12974 4338
rect 14130 4286 14142 4338
rect 14194 4286 14206 4338
rect 17490 4286 17502 4338
rect 17554 4286 17566 4338
rect 22978 4286 22990 4338
rect 23042 4286 23054 4338
rect 28802 4286 28814 4338
rect 28866 4286 28878 4338
rect 29922 4286 29934 4338
rect 29986 4286 29998 4338
rect 36978 4286 36990 4338
rect 37042 4286 37054 4338
rect 10110 4274 10162 4286
rect 42366 4274 42418 4286
rect 33294 4226 33346 4238
rect 2146 4174 2158 4226
rect 2210 4174 2222 4226
rect 11666 4174 11678 4226
rect 11730 4174 11742 4226
rect 20290 4174 20302 4226
rect 20354 4174 20366 4226
rect 33294 4162 33346 4174
rect 42142 4226 42194 4238
rect 42802 4174 42814 4226
rect 42866 4174 42878 4226
rect 42142 4162 42194 4174
rect 7422 4114 7474 4126
rect 4162 4062 4174 4114
rect 4226 4062 4238 4114
rect 7422 4050 7474 4062
rect 14702 4114 14754 4126
rect 14702 4050 14754 4062
rect 21086 4114 21138 4126
rect 21086 4050 21138 4062
rect 26462 4114 26514 4126
rect 26462 4050 26514 4062
rect 30830 4114 30882 4126
rect 30830 4050 30882 4062
rect 37998 4114 38050 4126
rect 37998 4050 38050 4062
rect 1344 3946 43568 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 43568 3946
rect 1344 3860 43568 3894
rect 10222 3666 10274 3678
rect 24782 3666 24834 3678
rect 2706 3614 2718 3666
rect 2770 3614 2782 3666
rect 18834 3614 18846 3666
rect 18898 3614 18910 3666
rect 10222 3602 10274 3614
rect 24782 3602 24834 3614
rect 27582 3666 27634 3678
rect 27582 3602 27634 3614
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 32734 3666 32786 3678
rect 32734 3602 32786 3614
rect 35534 3666 35586 3678
rect 35534 3602 35586 3614
rect 36990 3666 37042 3678
rect 36990 3602 37042 3614
rect 39342 3666 39394 3678
rect 39342 3602 39394 3614
rect 40798 3666 40850 3678
rect 40798 3602 40850 3614
rect 4834 3502 4846 3554
rect 4898 3502 4910 3554
rect 8754 3502 8766 3554
rect 8818 3502 8830 3554
rect 12114 3502 12126 3554
rect 12178 3502 12190 3554
rect 15922 3502 15934 3554
rect 15986 3502 15998 3554
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 21410 3502 21422 3554
rect 21474 3502 21486 3554
rect 27122 3502 27134 3554
rect 27186 3502 27198 3554
rect 28466 3502 28478 3554
rect 28530 3502 28542 3554
rect 33618 3502 33630 3554
rect 33682 3502 33694 3554
rect 35970 3502 35982 3554
rect 36034 3502 36046 3554
rect 39778 3502 39790 3554
rect 39842 3502 39854 3554
rect 1822 3442 1874 3454
rect 1822 3378 1874 3390
rect 31726 3442 31778 3454
rect 31726 3378 31778 3390
rect 32174 3442 32226 3454
rect 32174 3378 32226 3390
rect 33406 3442 33458 3454
rect 33406 3378 33458 3390
rect 7758 3330 7810 3342
rect 7758 3266 7810 3278
rect 15374 3330 15426 3342
rect 15374 3266 15426 3278
rect 22430 3330 22482 3342
rect 22430 3266 22482 3278
rect 1344 3162 43568 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 43568 3162
rect 1344 3076 43568 3110
<< via1 >>
rect 8542 41694 8594 41746
rect 9438 41694 9490 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 22430 41358 22482 41410
rect 25566 41358 25618 41410
rect 29374 41358 29426 41410
rect 33182 41358 33234 41410
rect 36990 41358 37042 41410
rect 40798 41358 40850 41410
rect 1934 41246 1986 41298
rect 5630 41246 5682 41298
rect 9438 41246 9490 41298
rect 11230 41246 11282 41298
rect 15038 41246 15090 41298
rect 17278 41246 17330 41298
rect 18398 41246 18450 41298
rect 19518 41246 19570 41298
rect 4286 41134 4338 41186
rect 4734 41134 4786 41186
rect 7870 41134 7922 41186
rect 8542 41134 8594 41186
rect 11678 41134 11730 41186
rect 12126 41134 12178 41186
rect 13134 41134 13186 41186
rect 14366 41134 14418 41186
rect 15262 41134 15314 41186
rect 16158 41134 16210 41186
rect 17726 41134 17778 41186
rect 18846 41134 18898 41186
rect 19966 41134 20018 41186
rect 20974 41134 21026 41186
rect 21422 41134 21474 41186
rect 24558 41134 24610 41186
rect 28366 41134 28418 41186
rect 32174 41134 32226 41186
rect 35982 41134 36034 41186
rect 39790 41134 39842 41186
rect 11454 41022 11506 41074
rect 43150 41022 43202 41074
rect 4958 40910 5010 40962
rect 7646 40910 7698 40962
rect 8766 40910 8818 40962
rect 12462 40910 12514 40962
rect 13470 40910 13522 40962
rect 14142 40910 14194 40962
rect 15598 40910 15650 40962
rect 16382 40910 16434 40962
rect 17502 40910 17554 40962
rect 18622 40910 18674 40962
rect 19742 40910 19794 40962
rect 20750 40910 20802 40962
rect 42814 40910 42866 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 9662 40574 9714 40626
rect 13134 40574 13186 40626
rect 13918 40574 13970 40626
rect 16606 40574 16658 40626
rect 21310 40574 21362 40626
rect 26350 40574 26402 40626
rect 29262 40574 29314 40626
rect 34078 40574 34130 40626
rect 36990 40574 37042 40626
rect 5406 40462 5458 40514
rect 7534 40462 7586 40514
rect 7870 40462 7922 40514
rect 8430 40462 8482 40514
rect 8766 40462 8818 40514
rect 11678 40462 11730 40514
rect 12686 40462 12738 40514
rect 24670 40462 24722 40514
rect 31502 40462 31554 40514
rect 4286 40350 4338 40402
rect 7198 40350 7250 40402
rect 11454 40350 11506 40402
rect 11902 40350 11954 40402
rect 12350 40350 12402 40402
rect 24446 40350 24498 40402
rect 25342 40350 25394 40402
rect 28254 40350 28306 40402
rect 31166 40350 31218 40402
rect 33070 40350 33122 40402
rect 35982 40350 36034 40402
rect 43150 40350 43202 40402
rect 15374 40238 15426 40290
rect 1934 40126 1986 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 6862 39790 6914 39842
rect 7534 39790 7586 39842
rect 24110 39790 24162 39842
rect 29374 39790 29426 39842
rect 33070 39790 33122 39842
rect 37998 39790 38050 39842
rect 40910 39790 40962 39842
rect 4622 39678 4674 39730
rect 6862 39678 6914 39730
rect 7198 39678 7250 39730
rect 11566 39678 11618 39730
rect 13470 39678 13522 39730
rect 20638 39678 20690 39730
rect 26238 39678 26290 39730
rect 1822 39566 1874 39618
rect 8654 39566 8706 39618
rect 16270 39566 16322 39618
rect 17726 39566 17778 39618
rect 23102 39566 23154 39618
rect 26014 39566 26066 39618
rect 27246 39566 27298 39618
rect 31278 39566 31330 39618
rect 32062 39566 32114 39618
rect 36990 39566 37042 39618
rect 39902 39566 39954 39618
rect 2494 39454 2546 39506
rect 8318 39454 8370 39506
rect 9438 39454 9490 39506
rect 15598 39454 15650 39506
rect 18510 39454 18562 39506
rect 21310 39454 21362 39506
rect 21646 39454 21698 39506
rect 22430 39454 22482 39506
rect 22766 39454 22818 39506
rect 27470 39454 27522 39506
rect 27806 39454 27858 39506
rect 28142 39454 28194 39506
rect 34974 39454 35026 39506
rect 35310 39454 35362 39506
rect 35982 39454 36034 39506
rect 36318 39454 36370 39506
rect 5070 39342 5122 39394
rect 5742 39342 5794 39394
rect 7646 39342 7698 39394
rect 7982 39342 8034 39394
rect 12014 39342 12066 39394
rect 12910 39342 12962 39394
rect 17390 39342 17442 39394
rect 26574 39342 26626 39394
rect 28702 39342 28754 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 8318 39006 8370 39058
rect 9662 39006 9714 39058
rect 15710 39006 15762 39058
rect 16830 39006 16882 39058
rect 18286 39006 18338 39058
rect 20414 39006 20466 39058
rect 23886 39006 23938 39058
rect 24670 39006 24722 39058
rect 25790 39006 25842 39058
rect 26686 39006 26738 39058
rect 27918 39006 27970 39058
rect 30830 39006 30882 39058
rect 31502 39006 31554 39058
rect 32174 39006 32226 39058
rect 33406 39006 33458 39058
rect 36430 39006 36482 39058
rect 19630 38894 19682 38946
rect 29150 38894 29202 38946
rect 38334 38894 38386 38946
rect 38670 38894 38722 38946
rect 39118 38894 39170 38946
rect 39454 38894 39506 38946
rect 1934 38782 1986 38834
rect 5182 38782 5234 38834
rect 9438 38782 9490 38834
rect 9886 38782 9938 38834
rect 10110 38782 10162 38834
rect 14926 38782 14978 38834
rect 15486 38782 15538 38834
rect 15598 38782 15650 38834
rect 16046 38782 16098 38834
rect 16494 38782 16546 38834
rect 18062 38782 18114 38834
rect 18286 38782 18338 38834
rect 18622 38782 18674 38834
rect 20190 38782 20242 38834
rect 24334 38782 24386 38834
rect 25230 38782 25282 38834
rect 27582 38782 27634 38834
rect 28926 38782 28978 38834
rect 29710 38782 29762 38834
rect 30046 38782 30098 38834
rect 30606 38782 30658 38834
rect 31166 38782 31218 38834
rect 31950 38782 32002 38834
rect 33070 38782 33122 38834
rect 35646 38782 35698 38834
rect 2606 38670 2658 38722
rect 4734 38670 4786 38722
rect 5854 38670 5906 38722
rect 7982 38670 8034 38722
rect 8766 38670 8818 38722
rect 12126 38670 12178 38722
rect 14254 38670 14306 38722
rect 16270 38670 16322 38722
rect 17614 38670 17666 38722
rect 19518 38670 19570 38722
rect 24110 38670 24162 38722
rect 26238 38670 26290 38722
rect 28366 38670 28418 38722
rect 25454 38558 25506 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 13918 38222 13970 38274
rect 15822 38222 15874 38274
rect 40910 38222 40962 38274
rect 1934 38110 1986 38162
rect 8430 38110 8482 38162
rect 11790 38110 11842 38162
rect 14478 38110 14530 38162
rect 16942 38110 16994 38162
rect 20750 38110 20802 38162
rect 25790 38110 25842 38162
rect 4286 37998 4338 38050
rect 4846 37998 4898 38050
rect 5742 37998 5794 38050
rect 11342 37998 11394 38050
rect 14030 37998 14082 38050
rect 14254 37998 14306 38050
rect 14814 37998 14866 38050
rect 15262 37998 15314 38050
rect 15486 37998 15538 38050
rect 16046 37998 16098 38050
rect 16382 37998 16434 38050
rect 17278 37998 17330 38050
rect 17838 37998 17890 38050
rect 22990 37998 23042 38050
rect 29262 37998 29314 38050
rect 39902 37998 39954 38050
rect 8094 37886 8146 37938
rect 10558 37886 10610 37938
rect 14702 37886 14754 37938
rect 16270 37886 16322 37938
rect 17614 37886 17666 37938
rect 18622 37886 18674 37938
rect 23662 37886 23714 37938
rect 28702 37886 28754 37938
rect 29486 37886 29538 37938
rect 5070 37774 5122 37826
rect 7534 37774 7586 37826
rect 7758 37774 7810 37826
rect 12910 37774 12962 37826
rect 13918 37774 13970 37826
rect 17390 37774 17442 37826
rect 26238 37774 26290 37826
rect 31502 37774 31554 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 7534 37438 7586 37490
rect 9774 37438 9826 37490
rect 15262 37438 15314 37490
rect 15486 37438 15538 37490
rect 15934 37438 15986 37490
rect 16270 37438 16322 37490
rect 17502 37438 17554 37490
rect 18286 37438 18338 37490
rect 18622 37438 18674 37490
rect 6750 37326 6802 37378
rect 8430 37326 8482 37378
rect 8654 37326 8706 37378
rect 10110 37326 10162 37378
rect 10558 37326 10610 37378
rect 12574 37326 12626 37378
rect 14590 37326 14642 37378
rect 17390 37326 17442 37378
rect 18062 37326 18114 37378
rect 19518 37326 19570 37378
rect 4286 37214 4338 37266
rect 6974 37214 7026 37266
rect 7422 37214 7474 37266
rect 7758 37214 7810 37266
rect 7982 37214 8034 37266
rect 8318 37214 8370 37266
rect 9438 37214 9490 37266
rect 9774 37214 9826 37266
rect 10446 37214 10498 37266
rect 12350 37214 12402 37266
rect 13358 37214 13410 37266
rect 13918 37214 13970 37266
rect 14366 37214 14418 37266
rect 15150 37214 15202 37266
rect 17726 37214 17778 37266
rect 17950 37214 18002 37266
rect 18398 37214 18450 37266
rect 18734 37214 18786 37266
rect 19070 37214 19122 37266
rect 6526 37102 6578 37154
rect 8990 37102 9042 37154
rect 11118 37102 11170 37154
rect 13022 37102 13074 37154
rect 1934 36990 1986 37042
rect 10558 36990 10610 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 15374 36654 15426 36706
rect 18286 36654 18338 36706
rect 41582 36654 41634 36706
rect 2046 36542 2098 36594
rect 5854 36542 5906 36594
rect 14926 36542 14978 36594
rect 23214 36542 23266 36594
rect 28590 36542 28642 36594
rect 4062 36430 4114 36482
rect 4846 36430 4898 36482
rect 5630 36430 5682 36482
rect 5966 36430 6018 36482
rect 6526 36430 6578 36482
rect 7310 36430 7362 36482
rect 7646 36430 7698 36482
rect 7758 36430 7810 36482
rect 8094 36430 8146 36482
rect 8430 36430 8482 36482
rect 9438 36430 9490 36482
rect 9774 36430 9826 36482
rect 15486 36430 15538 36482
rect 16830 36430 16882 36482
rect 20526 36430 20578 36482
rect 23326 36430 23378 36482
rect 23662 36430 23714 36482
rect 23886 36430 23938 36482
rect 24446 36430 24498 36482
rect 25678 36430 25730 36482
rect 40574 36430 40626 36482
rect 5070 36318 5122 36370
rect 6302 36318 6354 36370
rect 6750 36318 6802 36370
rect 6862 36318 6914 36370
rect 8766 36318 8818 36370
rect 16494 36318 16546 36370
rect 18174 36318 18226 36370
rect 20302 36318 20354 36370
rect 22542 36318 22594 36370
rect 22654 36318 22706 36370
rect 22878 36318 22930 36370
rect 23102 36318 23154 36370
rect 24334 36318 24386 36370
rect 26462 36318 26514 36370
rect 7422 36206 7474 36258
rect 7982 36206 8034 36258
rect 9550 36206 9602 36258
rect 10222 36206 10274 36258
rect 15374 36206 15426 36258
rect 16046 36206 16098 36258
rect 18286 36206 18338 36258
rect 18958 36206 19010 36258
rect 24222 36206 24274 36258
rect 25006 36206 25058 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 5070 35870 5122 35922
rect 5294 35870 5346 35922
rect 6750 35870 6802 35922
rect 7086 35870 7138 35922
rect 7422 35870 7474 35922
rect 12350 35870 12402 35922
rect 17726 35870 17778 35922
rect 21198 35870 21250 35922
rect 21534 35870 21586 35922
rect 22542 35870 22594 35922
rect 23326 35870 23378 35922
rect 4958 35758 5010 35810
rect 7198 35758 7250 35810
rect 7646 35758 7698 35810
rect 7758 35758 7810 35810
rect 12798 35758 12850 35810
rect 14590 35758 14642 35810
rect 21982 35758 22034 35810
rect 22990 35758 23042 35810
rect 23102 35758 23154 35810
rect 23662 35758 23714 35810
rect 25230 35758 25282 35810
rect 1822 35646 1874 35698
rect 8990 35646 9042 35698
rect 11902 35646 11954 35698
rect 13358 35646 13410 35698
rect 13918 35646 13970 35698
rect 14366 35646 14418 35698
rect 15262 35646 15314 35698
rect 17950 35646 18002 35698
rect 21870 35646 21922 35698
rect 22430 35646 22482 35698
rect 22766 35646 22818 35698
rect 23550 35646 23602 35698
rect 23998 35646 24050 35698
rect 24334 35646 24386 35698
rect 24558 35646 24610 35698
rect 25454 35646 25506 35698
rect 25790 35646 25842 35698
rect 28814 35646 28866 35698
rect 2494 35534 2546 35586
rect 4622 35534 4674 35586
rect 5630 35534 5682 35586
rect 8542 35534 8594 35586
rect 10894 35534 10946 35586
rect 13022 35534 13074 35586
rect 16270 35534 16322 35586
rect 20862 35534 20914 35586
rect 24222 35534 24274 35586
rect 25678 35534 25730 35586
rect 29598 35534 29650 35586
rect 31726 35534 31778 35586
rect 7086 35422 7138 35474
rect 21982 35422 22034 35474
rect 23662 35422 23714 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 15822 35086 15874 35138
rect 1934 34974 1986 35026
rect 4734 34974 4786 35026
rect 11006 34974 11058 35026
rect 11342 34974 11394 35026
rect 13582 34974 13634 35026
rect 21982 34974 22034 35026
rect 22990 34974 23042 35026
rect 23438 34974 23490 35026
rect 26350 34974 26402 35026
rect 28478 34974 28530 35026
rect 4286 34862 4338 34914
rect 5518 34862 5570 34914
rect 5966 34862 6018 34914
rect 6190 34862 6242 34914
rect 7422 34862 7474 34914
rect 10558 34862 10610 34914
rect 11566 34862 11618 34914
rect 11790 34862 11842 34914
rect 14926 34862 14978 34914
rect 15374 34862 15426 34914
rect 16942 34862 16994 34914
rect 22654 34862 22706 34914
rect 23774 34862 23826 34914
rect 24110 34862 24162 34914
rect 24558 34862 24610 34914
rect 25566 34862 25618 34914
rect 6862 34750 6914 34802
rect 7086 34750 7138 34802
rect 10222 34750 10274 34802
rect 14590 34750 14642 34802
rect 15710 34750 15762 34802
rect 20190 34750 20242 34802
rect 20526 34750 20578 34802
rect 22318 34750 22370 34802
rect 22430 34750 22482 34802
rect 24334 34750 24386 34802
rect 4622 34638 4674 34690
rect 5742 34638 5794 34690
rect 7310 34638 7362 34690
rect 11454 34638 11506 34690
rect 12014 34638 12066 34690
rect 12126 34638 12178 34690
rect 12798 34638 12850 34690
rect 15822 34638 15874 34690
rect 16494 34638 16546 34690
rect 17390 34638 17442 34690
rect 17726 34638 17778 34690
rect 23886 34638 23938 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 2830 34302 2882 34354
rect 17950 34302 18002 34354
rect 18734 34302 18786 34354
rect 20638 34302 20690 34354
rect 24110 34302 24162 34354
rect 26910 34302 26962 34354
rect 28254 34302 28306 34354
rect 29934 34302 29986 34354
rect 30830 34302 30882 34354
rect 32510 34302 32562 34354
rect 2046 34190 2098 34242
rect 2718 34190 2770 34242
rect 5742 34190 5794 34242
rect 7646 34190 7698 34242
rect 19630 34190 19682 34242
rect 23774 34190 23826 34242
rect 23886 34190 23938 34242
rect 28926 34190 28978 34242
rect 29150 34190 29202 34242
rect 31726 34190 31778 34242
rect 2158 34078 2210 34130
rect 2494 34078 2546 34130
rect 3278 34078 3330 34130
rect 6526 34078 6578 34130
rect 6974 34078 7026 34130
rect 7422 34078 7474 34130
rect 12798 34078 12850 34130
rect 17390 34078 17442 34130
rect 17614 34078 17666 34130
rect 19518 34078 19570 34130
rect 20302 34078 20354 34130
rect 31950 34078 32002 34130
rect 3614 33966 3666 34018
rect 7758 33966 7810 34018
rect 8318 33966 8370 34018
rect 10558 33966 10610 34018
rect 13358 33966 13410 34018
rect 19070 33966 19122 34018
rect 24446 33966 24498 34018
rect 30382 33966 30434 34018
rect 33182 33966 33234 34018
rect 3054 33854 3106 33906
rect 6750 33854 6802 33906
rect 28590 33854 28642 33906
rect 31166 33854 31218 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 25566 33518 25618 33570
rect 27358 33518 27410 33570
rect 1934 33406 1986 33458
rect 6750 33406 6802 33458
rect 7310 33406 7362 33458
rect 11902 33406 11954 33458
rect 12350 33406 12402 33458
rect 16942 33406 16994 33458
rect 30158 33406 30210 33458
rect 4286 33294 4338 33346
rect 4622 33294 4674 33346
rect 4958 33294 5010 33346
rect 9774 33294 9826 33346
rect 10894 33294 10946 33346
rect 11230 33294 11282 33346
rect 11566 33294 11618 33346
rect 14702 33294 14754 33346
rect 15262 33294 15314 33346
rect 15710 33294 15762 33346
rect 16494 33294 16546 33346
rect 19742 33294 19794 33346
rect 24446 33294 24498 33346
rect 25230 33294 25282 33346
rect 26574 33294 26626 33346
rect 27694 33294 27746 33346
rect 7758 33182 7810 33234
rect 8094 33182 8146 33234
rect 10222 33182 10274 33234
rect 10782 33182 10834 33234
rect 14254 33182 14306 33234
rect 16270 33182 16322 33234
rect 19070 33182 19122 33234
rect 24670 33182 24722 33234
rect 27918 33182 27970 33234
rect 28478 33182 28530 33234
rect 4734 33070 4786 33122
rect 9662 33070 9714 33122
rect 9886 33070 9938 33122
rect 9998 33070 10050 33122
rect 10670 33070 10722 33122
rect 11342 33070 11394 33122
rect 12910 33070 12962 33122
rect 13806 33070 13858 33122
rect 14030 33070 14082 33122
rect 26126 33070 26178 33122
rect 29262 33070 29314 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 2382 32734 2434 32786
rect 5294 32734 5346 32786
rect 6414 32734 6466 32786
rect 8654 32734 8706 32786
rect 10334 32734 10386 32786
rect 14590 32734 14642 32786
rect 16718 32734 16770 32786
rect 18174 32734 18226 32786
rect 2046 32622 2098 32674
rect 2270 32622 2322 32674
rect 6190 32622 6242 32674
rect 8318 32622 8370 32674
rect 10558 32622 10610 32674
rect 12574 32622 12626 32674
rect 14366 32622 14418 32674
rect 16270 32622 16322 32674
rect 2830 32510 2882 32562
rect 5518 32510 5570 32562
rect 6078 32510 6130 32562
rect 6638 32510 6690 32562
rect 7198 32510 7250 32562
rect 7646 32510 7698 32562
rect 7758 32510 7810 32562
rect 8542 32510 8594 32562
rect 8766 32510 8818 32562
rect 8878 32510 8930 32562
rect 11230 32510 11282 32562
rect 11678 32510 11730 32562
rect 12350 32510 12402 32562
rect 13918 32510 13970 32562
rect 14926 32510 14978 32562
rect 15150 32510 15202 32562
rect 15822 32510 15874 32562
rect 17502 32510 17554 32562
rect 18062 32510 18114 32562
rect 18622 32510 18674 32562
rect 26686 32510 26738 32562
rect 3278 32398 3330 32450
rect 3726 32398 3778 32450
rect 7982 32398 8034 32450
rect 11006 32398 11058 32450
rect 13134 32398 13186 32450
rect 13582 32398 13634 32450
rect 17726 32398 17778 32450
rect 24670 32398 24722 32450
rect 27246 32398 27298 32450
rect 2494 32286 2546 32338
rect 6974 32286 7026 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 13806 31950 13858 32002
rect 14478 31950 14530 32002
rect 1934 31838 1986 31890
rect 7086 31838 7138 31890
rect 8094 31838 8146 31890
rect 9886 31838 9938 31890
rect 24222 31838 24274 31890
rect 32062 31838 32114 31890
rect 4062 31726 4114 31778
rect 5966 31726 6018 31778
rect 6526 31726 6578 31778
rect 7310 31726 7362 31778
rect 7870 31726 7922 31778
rect 9550 31726 9602 31778
rect 10222 31726 10274 31778
rect 15374 31726 15426 31778
rect 15822 31726 15874 31778
rect 21310 31726 21362 31778
rect 24558 31726 24610 31778
rect 24782 31726 24834 31778
rect 25118 31726 25170 31778
rect 29262 31726 29314 31778
rect 7646 31614 7698 31666
rect 8318 31614 8370 31666
rect 9998 31614 10050 31666
rect 10558 31614 10610 31666
rect 11342 31614 11394 31666
rect 17054 31614 17106 31666
rect 22094 31614 22146 31666
rect 29934 31614 29986 31666
rect 37326 31614 37378 31666
rect 42814 31614 42866 31666
rect 43150 31614 43202 31666
rect 6190 31502 6242 31554
rect 8206 31502 8258 31554
rect 9214 31502 9266 31554
rect 9774 31502 9826 31554
rect 10894 31502 10946 31554
rect 14030 31502 14082 31554
rect 14478 31502 14530 31554
rect 14926 31502 14978 31554
rect 16158 31502 16210 31554
rect 16494 31502 16546 31554
rect 36990 31502 37042 31554
rect 42590 31502 42642 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4062 31166 4114 31218
rect 5406 31166 5458 31218
rect 20302 31166 20354 31218
rect 20974 31166 21026 31218
rect 23662 31166 23714 31218
rect 27694 31166 27746 31218
rect 28142 31166 28194 31218
rect 28702 31166 28754 31218
rect 31838 31166 31890 31218
rect 2606 31054 2658 31106
rect 3054 31054 3106 31106
rect 9438 31054 9490 31106
rect 9774 31054 9826 31106
rect 10110 31054 10162 31106
rect 20414 31054 20466 31106
rect 23102 31054 23154 31106
rect 28366 31054 28418 31106
rect 32286 31054 32338 31106
rect 3278 30942 3330 30994
rect 3726 30942 3778 30994
rect 9886 30942 9938 30994
rect 10222 30942 10274 30994
rect 12238 30942 12290 30994
rect 14142 30942 14194 30994
rect 20638 30942 20690 30994
rect 20974 30942 21026 30994
rect 21310 30942 21362 30994
rect 21982 30942 22034 30994
rect 22206 30942 22258 30994
rect 22654 30942 22706 30994
rect 28030 30942 28082 30994
rect 28478 30942 28530 30994
rect 28814 30942 28866 30994
rect 29150 30942 29202 30994
rect 31502 30942 31554 30994
rect 1822 30830 1874 30882
rect 2382 30830 2434 30882
rect 4622 30830 4674 30882
rect 14366 30830 14418 30882
rect 16158 30830 16210 30882
rect 22430 30830 22482 30882
rect 24222 30830 24274 30882
rect 31054 30830 31106 30882
rect 31278 30830 31330 30882
rect 2718 30718 2770 30770
rect 10670 30718 10722 30770
rect 11678 30718 11730 30770
rect 12014 30718 12066 30770
rect 20302 30718 20354 30770
rect 23214 30718 23266 30770
rect 23438 30718 23490 30770
rect 24222 30718 24274 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 6078 30382 6130 30434
rect 11790 30382 11842 30434
rect 20078 30382 20130 30434
rect 30494 30382 30546 30434
rect 30942 30382 30994 30434
rect 1934 30270 1986 30322
rect 16270 30270 16322 30322
rect 17614 30270 17666 30322
rect 18062 30270 18114 30322
rect 26462 30270 26514 30322
rect 34078 30270 34130 30322
rect 34638 30270 34690 30322
rect 4846 30158 4898 30210
rect 12014 30158 12066 30210
rect 12238 30158 12290 30210
rect 15486 30158 15538 30210
rect 15710 30158 15762 30210
rect 15934 30158 15986 30210
rect 16158 30158 16210 30210
rect 16718 30158 16770 30210
rect 16942 30158 16994 30210
rect 17054 30158 17106 30210
rect 20862 30158 20914 30210
rect 21758 30158 21810 30210
rect 22654 30158 22706 30210
rect 23550 30158 23602 30210
rect 24334 30158 24386 30210
rect 27918 30158 27970 30210
rect 29486 30158 29538 30210
rect 29710 30158 29762 30210
rect 30046 30158 30098 30210
rect 30270 30158 30322 30210
rect 30830 30158 30882 30210
rect 31166 30158 31218 30210
rect 34414 30158 34466 30210
rect 34974 30158 35026 30210
rect 4062 30046 4114 30098
rect 6302 30046 6354 30098
rect 11118 30046 11170 30098
rect 11342 30046 11394 30098
rect 11566 30046 11618 30098
rect 16382 30046 16434 30098
rect 17390 30046 17442 30098
rect 20190 30046 20242 30098
rect 20526 30046 20578 30098
rect 20638 30046 20690 30098
rect 22318 30046 22370 30098
rect 22990 30046 23042 30098
rect 27582 30046 27634 30098
rect 29150 30046 29202 30098
rect 29934 30046 29986 30098
rect 31950 30046 32002 30098
rect 5742 29934 5794 29986
rect 6750 29934 6802 29986
rect 11678 29934 11730 29986
rect 15150 29934 15202 29986
rect 17502 29934 17554 29986
rect 18398 29934 18450 29986
rect 19630 29934 19682 29986
rect 20078 29934 20130 29986
rect 21982 29934 22034 29986
rect 22430 29934 22482 29986
rect 26798 29934 26850 29986
rect 27134 29934 27186 29986
rect 27694 29934 27746 29986
rect 28254 29934 28306 29986
rect 29262 29934 29314 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 2046 29598 2098 29650
rect 2606 29598 2658 29650
rect 3838 29598 3890 29650
rect 4174 29598 4226 29650
rect 17726 29598 17778 29650
rect 20750 29598 20802 29650
rect 21198 29598 21250 29650
rect 26574 29598 26626 29650
rect 2494 29486 2546 29538
rect 2718 29486 2770 29538
rect 3054 29486 3106 29538
rect 4846 29486 4898 29538
rect 5294 29486 5346 29538
rect 5518 29486 5570 29538
rect 6078 29486 6130 29538
rect 16718 29486 16770 29538
rect 17838 29486 17890 29538
rect 18062 29486 18114 29538
rect 19070 29486 19122 29538
rect 1822 29374 1874 29426
rect 3278 29374 3330 29426
rect 3838 29374 3890 29426
rect 4398 29374 4450 29426
rect 5182 29374 5234 29426
rect 6190 29374 6242 29426
rect 10110 29374 10162 29426
rect 10334 29374 10386 29426
rect 15374 29374 15426 29426
rect 16606 29374 16658 29426
rect 16942 29374 16994 29426
rect 17390 29374 17442 29426
rect 17614 29374 17666 29426
rect 20414 29374 20466 29426
rect 26238 29374 26290 29426
rect 5630 29262 5682 29314
rect 6638 29262 6690 29314
rect 11790 29262 11842 29314
rect 18510 29262 18562 29314
rect 27134 29262 27186 29314
rect 28926 29262 28978 29314
rect 34078 29262 34130 29314
rect 3614 29150 3666 29202
rect 5182 29150 5234 29202
rect 6078 29150 6130 29202
rect 9774 29150 9826 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 4622 28814 4674 28866
rect 11342 28814 11394 28866
rect 17950 28814 18002 28866
rect 30830 28814 30882 28866
rect 1934 28702 1986 28754
rect 6302 28702 6354 28754
rect 26910 28702 26962 28754
rect 33742 28702 33794 28754
rect 4286 28590 4338 28642
rect 8430 28590 8482 28642
rect 9102 28590 9154 28642
rect 10334 28590 10386 28642
rect 10446 28590 10498 28642
rect 10894 28590 10946 28642
rect 11118 28590 11170 28642
rect 11454 28590 11506 28642
rect 11902 28590 11954 28642
rect 13470 28590 13522 28642
rect 13918 28590 13970 28642
rect 14142 28590 14194 28642
rect 17390 28590 17442 28642
rect 17726 28590 17778 28642
rect 18286 28590 18338 28642
rect 20638 28590 20690 28642
rect 25566 28590 25618 28642
rect 26014 28590 26066 28642
rect 27246 28590 27298 28642
rect 29486 28590 29538 28642
rect 29822 28590 29874 28642
rect 30158 28590 30210 28642
rect 30494 28590 30546 28642
rect 32734 28590 32786 28642
rect 32846 28590 32898 28642
rect 4958 28478 5010 28530
rect 12238 28478 12290 28530
rect 14030 28478 14082 28530
rect 16270 28478 16322 28530
rect 16942 28478 16994 28530
rect 25342 28478 25394 28530
rect 26350 28478 26402 28530
rect 27806 28478 27858 28530
rect 29150 28478 29202 28530
rect 30718 28478 30770 28530
rect 4734 28366 4786 28418
rect 10782 28366 10834 28418
rect 15150 28366 15202 28418
rect 15598 28366 15650 28418
rect 15934 28366 15986 28418
rect 16606 28366 16658 28418
rect 20302 28366 20354 28418
rect 27358 28366 27410 28418
rect 27582 28366 27634 28418
rect 27918 28366 27970 28418
rect 28142 28366 28194 28418
rect 28590 28366 28642 28418
rect 29262 28366 29314 28418
rect 30270 28366 30322 28418
rect 30830 28366 30882 28418
rect 31502 28366 31554 28418
rect 33294 28366 33346 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 11678 28030 11730 28082
rect 12910 28030 12962 28082
rect 16270 28030 16322 28082
rect 17502 28030 17554 28082
rect 10782 27918 10834 27970
rect 12462 27918 12514 27970
rect 22206 27918 22258 27970
rect 30942 27918 30994 27970
rect 33854 27918 33906 27970
rect 4286 27806 4338 27858
rect 10558 27806 10610 27858
rect 11118 27806 11170 27858
rect 11790 27806 11842 27858
rect 12126 27806 12178 27858
rect 21646 27806 21698 27858
rect 21870 27806 21922 27858
rect 27246 27806 27298 27858
rect 33070 27806 33122 27858
rect 4734 27694 4786 27746
rect 11342 27694 11394 27746
rect 12350 27694 12402 27746
rect 21758 27694 21810 27746
rect 26910 27694 26962 27746
rect 35982 27694 36034 27746
rect 1934 27582 1986 27634
rect 11566 27582 11618 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 15150 27246 15202 27298
rect 29374 27246 29426 27298
rect 29710 27246 29762 27298
rect 30158 27246 30210 27298
rect 34414 27246 34466 27298
rect 34750 27246 34802 27298
rect 2046 27134 2098 27186
rect 9998 27134 10050 27186
rect 12126 27134 12178 27186
rect 16718 27134 16770 27186
rect 22654 27134 22706 27186
rect 24782 27134 24834 27186
rect 25678 27134 25730 27186
rect 33630 27134 33682 27186
rect 35198 27134 35250 27186
rect 4174 27022 4226 27074
rect 6750 27022 6802 27074
rect 7870 27022 7922 27074
rect 12798 27022 12850 27074
rect 14814 27022 14866 27074
rect 15710 27022 15762 27074
rect 15934 27022 15986 27074
rect 16494 27022 16546 27074
rect 17166 27022 17218 27074
rect 20526 27022 20578 27074
rect 21310 27022 21362 27074
rect 21646 27022 21698 27074
rect 21982 27022 22034 27074
rect 25230 27022 25282 27074
rect 28590 27022 28642 27074
rect 29150 27022 29202 27074
rect 30046 27022 30098 27074
rect 30830 27022 30882 27074
rect 34190 27022 34242 27074
rect 7534 26910 7586 26962
rect 14478 26910 14530 26962
rect 15598 26910 15650 26962
rect 16270 26910 16322 26962
rect 16942 26910 16994 26962
rect 20638 26910 20690 26962
rect 27806 26910 27858 26962
rect 31502 26910 31554 26962
rect 6862 26798 6914 26850
rect 16158 26798 16210 26850
rect 17726 26798 17778 26850
rect 20862 26798 20914 26850
rect 21422 26798 21474 26850
rect 30158 26798 30210 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 6974 26462 7026 26514
rect 15486 26462 15538 26514
rect 16270 26462 16322 26514
rect 25790 26462 25842 26514
rect 27806 26462 27858 26514
rect 28814 26462 28866 26514
rect 29262 26462 29314 26514
rect 34302 26462 34354 26514
rect 5854 26350 5906 26402
rect 7086 26350 7138 26402
rect 7982 26350 8034 26402
rect 15822 26350 15874 26402
rect 16382 26350 16434 26402
rect 18062 26350 18114 26402
rect 27358 26350 27410 26402
rect 27582 26350 27634 26402
rect 6526 26238 6578 26290
rect 7310 26238 7362 26290
rect 7758 26238 7810 26290
rect 11566 26238 11618 26290
rect 11902 26238 11954 26290
rect 12126 26238 12178 26290
rect 12350 26238 12402 26290
rect 12574 26238 12626 26290
rect 16606 26238 16658 26290
rect 16830 26238 16882 26290
rect 22542 26238 22594 26290
rect 22766 26238 22818 26290
rect 23214 26238 23266 26290
rect 23326 26238 23378 26290
rect 25454 26238 25506 26290
rect 28030 26238 28082 26290
rect 3726 26126 3778 26178
rect 11342 26126 11394 26178
rect 12462 26126 12514 26178
rect 13022 26126 13074 26178
rect 16270 26126 16322 26178
rect 17502 26126 17554 26178
rect 19630 26126 19682 26178
rect 21758 26126 21810 26178
rect 22990 26126 23042 26178
rect 25230 26126 25282 26178
rect 33854 26126 33906 26178
rect 7534 26014 7586 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 22318 25678 22370 25730
rect 27134 25678 27186 25730
rect 1710 25566 1762 25618
rect 5854 25566 5906 25618
rect 7310 25566 7362 25618
rect 23102 25566 23154 25618
rect 32174 25566 32226 25618
rect 4622 25454 4674 25506
rect 7086 25454 7138 25506
rect 7534 25454 7586 25506
rect 8094 25454 8146 25506
rect 12350 25454 12402 25506
rect 12462 25454 12514 25506
rect 15598 25454 15650 25506
rect 20526 25454 20578 25506
rect 21646 25454 21698 25506
rect 22094 25454 22146 25506
rect 22654 25454 22706 25506
rect 31614 25454 31666 25506
rect 3838 25342 3890 25394
rect 5742 25342 5794 25394
rect 7758 25342 7810 25394
rect 12574 25342 12626 25394
rect 15710 25342 15762 25394
rect 16718 25342 16770 25394
rect 21310 25342 21362 25394
rect 21422 25342 21474 25394
rect 27022 25342 27074 25394
rect 6974 25230 7026 25282
rect 10558 25230 10610 25282
rect 11902 25230 11954 25282
rect 15262 25230 15314 25282
rect 16494 25230 16546 25282
rect 17054 25230 17106 25282
rect 17502 25230 17554 25282
rect 19854 25230 19906 25282
rect 20302 25230 20354 25282
rect 20638 25230 20690 25282
rect 20862 25230 20914 25282
rect 31726 25230 31778 25282
rect 33854 25230 33906 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 10558 24894 10610 24946
rect 12686 24894 12738 24946
rect 12798 24894 12850 24946
rect 13470 24894 13522 24946
rect 15150 24894 15202 24946
rect 15262 24894 15314 24946
rect 16606 24894 16658 24946
rect 17614 24894 17666 24946
rect 20078 24894 20130 24946
rect 23438 24894 23490 24946
rect 23886 24894 23938 24946
rect 28926 24894 28978 24946
rect 33182 24894 33234 24946
rect 6750 24782 6802 24834
rect 7646 24782 7698 24834
rect 9550 24782 9602 24834
rect 9998 24782 10050 24834
rect 15486 24782 15538 24834
rect 16830 24782 16882 24834
rect 19294 24782 19346 24834
rect 19630 24782 19682 24834
rect 34302 24782 34354 24834
rect 4286 24670 4338 24722
rect 7310 24670 7362 24722
rect 9774 24670 9826 24722
rect 10110 24670 10162 24722
rect 10894 24670 10946 24722
rect 12238 24670 12290 24722
rect 12462 24670 12514 24722
rect 12574 24670 12626 24722
rect 14814 24670 14866 24722
rect 15038 24670 15090 24722
rect 16158 24670 16210 24722
rect 16382 24670 16434 24722
rect 17950 24670 18002 24722
rect 18286 24670 18338 24722
rect 23326 24670 23378 24722
rect 28478 24670 28530 24722
rect 29374 24670 29426 24722
rect 6862 24558 6914 24610
rect 6974 24558 7026 24610
rect 9886 24558 9938 24610
rect 11118 24558 11170 24610
rect 11902 24558 11954 24610
rect 14590 24558 14642 24610
rect 16494 24558 16546 24610
rect 18846 24558 18898 24610
rect 25566 24558 25618 24610
rect 27694 24558 27746 24610
rect 30158 24558 30210 24610
rect 32286 24558 32338 24610
rect 33630 24558 33682 24610
rect 1934 24446 1986 24498
rect 7198 24446 7250 24498
rect 33630 24446 33682 24498
rect 33966 24670 34018 24722
rect 34078 24446 34130 24498
rect 34414 24446 34466 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 5742 24110 5794 24162
rect 1710 23998 1762 24050
rect 3838 23998 3890 24050
rect 11118 23998 11170 24050
rect 11678 23998 11730 24050
rect 16494 23998 16546 24050
rect 29374 23998 29426 24050
rect 32958 23998 33010 24050
rect 36206 23998 36258 24050
rect 4622 23886 4674 23938
rect 9886 23886 9938 23938
rect 10110 23886 10162 23938
rect 10334 23886 10386 23938
rect 10558 23886 10610 23938
rect 11454 23886 11506 23938
rect 16046 23886 16098 23938
rect 17166 23886 17218 23938
rect 17502 23886 17554 23938
rect 18622 23886 18674 23938
rect 29710 23886 29762 23938
rect 33294 23886 33346 23938
rect 5630 23774 5682 23826
rect 10782 23774 10834 23826
rect 15486 23774 15538 23826
rect 16830 23774 16882 23826
rect 34078 23774 34130 23826
rect 9774 23662 9826 23714
rect 15150 23662 15202 23714
rect 17614 23662 17666 23714
rect 17838 23662 17890 23714
rect 18286 23662 18338 23714
rect 30046 23662 30098 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 8430 23326 8482 23378
rect 20190 23326 20242 23378
rect 29486 23326 29538 23378
rect 30942 23326 30994 23378
rect 32510 23326 32562 23378
rect 33294 23326 33346 23378
rect 42814 23326 42866 23378
rect 5742 23214 5794 23266
rect 20078 23214 20130 23266
rect 34526 23214 34578 23266
rect 6526 23102 6578 23154
rect 28702 23102 28754 23154
rect 29038 23102 29090 23154
rect 29598 23102 29650 23154
rect 29822 23102 29874 23154
rect 30158 23102 30210 23154
rect 30494 23102 30546 23154
rect 30718 23102 30770 23154
rect 33070 23102 33122 23154
rect 33742 23102 33794 23154
rect 43150 23102 43202 23154
rect 3614 22990 3666 23042
rect 8318 22990 8370 23042
rect 10670 22990 10722 23042
rect 27358 22990 27410 23042
rect 28030 22990 28082 23042
rect 31390 22990 31442 23042
rect 36654 22990 36706 23042
rect 42590 22990 42642 23042
rect 28366 22878 28418 22930
rect 28702 22878 28754 22930
rect 29262 22878 29314 22930
rect 30606 22878 30658 22930
rect 33406 22878 33458 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 1934 22542 1986 22594
rect 29486 22542 29538 22594
rect 9326 22430 9378 22482
rect 10222 22430 10274 22482
rect 11118 22430 11170 22482
rect 12014 22430 12066 22482
rect 20750 22430 20802 22482
rect 25566 22430 25618 22482
rect 27694 22430 27746 22482
rect 29934 22430 29986 22482
rect 33742 22430 33794 22482
rect 34750 22430 34802 22482
rect 4286 22318 4338 22370
rect 9662 22318 9714 22370
rect 10110 22318 10162 22370
rect 10334 22318 10386 22370
rect 10670 22318 10722 22370
rect 10894 22318 10946 22370
rect 11678 22318 11730 22370
rect 21422 22318 21474 22370
rect 22766 22318 22818 22370
rect 26798 22318 26850 22370
rect 26910 22318 26962 22370
rect 27134 22318 27186 22370
rect 27358 22318 27410 22370
rect 33854 22318 33906 22370
rect 34190 22318 34242 22370
rect 34974 22318 35026 22370
rect 35422 22318 35474 22370
rect 11342 22206 11394 22258
rect 14926 22206 14978 22258
rect 21310 22206 21362 22258
rect 21758 22206 21810 22258
rect 23438 22206 23490 22258
rect 28030 22206 28082 22258
rect 28590 22206 28642 22258
rect 29150 22206 29202 22258
rect 33630 22206 33682 22258
rect 34638 22206 34690 22258
rect 9886 22094 9938 22146
rect 10558 22094 10610 22146
rect 14590 22094 14642 22146
rect 15038 22094 15090 22146
rect 15262 22094 15314 22146
rect 26014 22094 26066 22146
rect 27022 22094 27074 22146
rect 27806 22094 27858 22146
rect 29374 22094 29426 22146
rect 30382 22094 30434 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 10110 21758 10162 21810
rect 11342 21758 11394 21810
rect 11790 21758 11842 21810
rect 17614 21758 17666 21810
rect 18174 21758 18226 21810
rect 27022 21758 27074 21810
rect 27694 21758 27746 21810
rect 34414 21758 34466 21810
rect 9998 21646 10050 21698
rect 10894 21646 10946 21698
rect 16270 21646 16322 21698
rect 19294 21646 19346 21698
rect 25902 21646 25954 21698
rect 27358 21646 27410 21698
rect 28142 21646 28194 21698
rect 28366 21646 28418 21698
rect 4174 21534 4226 21586
rect 8990 21534 9042 21586
rect 10670 21534 10722 21586
rect 12798 21534 12850 21586
rect 15934 21534 15986 21586
rect 17502 21534 17554 21586
rect 24334 21534 24386 21586
rect 25342 21534 25394 21586
rect 26686 21534 26738 21586
rect 28814 21534 28866 21586
rect 1934 21422 1986 21474
rect 5070 21422 5122 21474
rect 5182 21422 5234 21474
rect 6078 21422 6130 21474
rect 8206 21422 8258 21474
rect 10222 21422 10274 21474
rect 11230 21422 11282 21474
rect 13470 21422 13522 21474
rect 15598 21422 15650 21474
rect 16830 21422 16882 21474
rect 29374 21422 29426 21474
rect 31838 21422 31890 21474
rect 10446 21310 10498 21362
rect 17614 21310 17666 21362
rect 25790 21310 25842 21362
rect 28030 21310 28082 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 27470 20974 27522 21026
rect 29934 20974 29986 21026
rect 31838 20974 31890 21026
rect 32174 20974 32226 21026
rect 1710 20862 1762 20914
rect 3838 20862 3890 20914
rect 12910 20862 12962 20914
rect 14254 20862 14306 20914
rect 18286 20862 18338 20914
rect 25230 20862 25282 20914
rect 25678 20862 25730 20914
rect 28366 20862 28418 20914
rect 30942 20862 30994 20914
rect 31502 20862 31554 20914
rect 35086 20862 35138 20914
rect 4622 20750 4674 20802
rect 12574 20750 12626 20802
rect 14926 20750 14978 20802
rect 15710 20750 15762 20802
rect 15934 20750 15986 20802
rect 16942 20750 16994 20802
rect 17838 20750 17890 20802
rect 18846 20750 18898 20802
rect 21534 20750 21586 20802
rect 21646 20750 21698 20802
rect 21870 20750 21922 20802
rect 22990 20750 23042 20802
rect 23102 20750 23154 20802
rect 23326 20750 23378 20802
rect 24110 20750 24162 20802
rect 24558 20750 24610 20802
rect 27134 20750 27186 20802
rect 27694 20750 27746 20802
rect 27918 20750 27970 20802
rect 29262 20750 29314 20802
rect 30270 20750 30322 20802
rect 33854 20750 33906 20802
rect 34190 20750 34242 20802
rect 7758 20638 7810 20690
rect 10110 20638 10162 20690
rect 13470 20638 13522 20690
rect 13582 20638 13634 20690
rect 14590 20638 14642 20690
rect 16494 20638 16546 20690
rect 18398 20638 18450 20690
rect 22094 20638 22146 20690
rect 22654 20638 22706 20690
rect 23774 20638 23826 20690
rect 24446 20638 24498 20690
rect 29598 20638 29650 20690
rect 29822 20638 29874 20690
rect 31614 20638 31666 20690
rect 34526 20638 34578 20690
rect 5070 20526 5122 20578
rect 8094 20526 8146 20578
rect 13806 20526 13858 20578
rect 14478 20526 14530 20578
rect 21310 20526 21362 20578
rect 23438 20526 23490 20578
rect 24670 20526 24722 20578
rect 27806 20526 27858 20578
rect 32286 20526 32338 20578
rect 32398 20526 32450 20578
rect 32958 20526 33010 20578
rect 34190 20526 34242 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 10446 20190 10498 20242
rect 12014 20190 12066 20242
rect 14814 20190 14866 20242
rect 15598 20190 15650 20242
rect 29262 20190 29314 20242
rect 30046 20190 30098 20242
rect 30382 20190 30434 20242
rect 31278 20190 31330 20242
rect 13246 20078 13298 20130
rect 13918 20078 13970 20130
rect 21422 20078 21474 20130
rect 23886 20078 23938 20130
rect 24110 20078 24162 20130
rect 28030 20078 28082 20130
rect 29038 20078 29090 20130
rect 30270 20078 30322 20130
rect 30718 20078 30770 20130
rect 32062 20078 32114 20130
rect 4286 19966 4338 20018
rect 5966 19966 6018 20018
rect 9550 19966 9602 20018
rect 10110 19966 10162 20018
rect 11006 19966 11058 20018
rect 12574 19966 12626 20018
rect 13134 19966 13186 20018
rect 14254 19966 14306 20018
rect 15262 19966 15314 20018
rect 15710 19966 15762 20018
rect 16046 19966 16098 20018
rect 16382 19966 16434 20018
rect 22206 19966 22258 20018
rect 23102 19966 23154 20018
rect 29486 19966 29538 20018
rect 29710 19966 29762 20018
rect 31502 19966 31554 20018
rect 31726 19966 31778 20018
rect 32510 19966 32562 20018
rect 33182 19966 33234 20018
rect 1934 19854 1986 19906
rect 6414 19854 6466 19906
rect 16830 19854 16882 19906
rect 17502 19854 17554 19906
rect 19294 19854 19346 19906
rect 22766 19854 22818 19906
rect 24558 19854 24610 19906
rect 25342 19854 25394 19906
rect 28478 19854 28530 19906
rect 29374 19854 29426 19906
rect 31614 19854 31666 19906
rect 33966 19854 34018 19906
rect 36094 19854 36146 19906
rect 36542 19854 36594 19906
rect 10782 19742 10834 19794
rect 15934 19742 15986 19794
rect 23102 19742 23154 19794
rect 23438 19742 23490 19794
rect 23774 19742 23826 19794
rect 27918 19742 27970 19794
rect 28366 19742 28418 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 16046 19406 16098 19458
rect 21758 19406 21810 19458
rect 23102 19406 23154 19458
rect 34750 19406 34802 19458
rect 35086 19406 35138 19458
rect 35422 19406 35474 19458
rect 1934 19294 1986 19346
rect 12238 19294 12290 19346
rect 14030 19294 14082 19346
rect 15038 19294 15090 19346
rect 17054 19294 17106 19346
rect 17390 19294 17442 19346
rect 20750 19294 20802 19346
rect 24334 19294 24386 19346
rect 28590 19294 28642 19346
rect 35758 19294 35810 19346
rect 36206 19294 36258 19346
rect 36430 19294 36482 19346
rect 3950 19182 4002 19234
rect 5742 19182 5794 19234
rect 6638 19182 6690 19234
rect 6974 19182 7026 19234
rect 7310 19182 7362 19234
rect 10110 19182 10162 19234
rect 10558 19182 10610 19234
rect 11230 19182 11282 19234
rect 11566 19182 11618 19234
rect 12350 19182 12402 19234
rect 13582 19182 13634 19234
rect 13918 19182 13970 19234
rect 16046 19182 16098 19234
rect 20302 19182 20354 19234
rect 21534 19182 21586 19234
rect 22318 19182 22370 19234
rect 22654 19182 22706 19234
rect 22878 19182 22930 19234
rect 23326 19182 23378 19234
rect 23886 19182 23938 19234
rect 24782 19182 24834 19234
rect 29150 19182 29202 19234
rect 36094 19182 36146 19234
rect 37102 19182 37154 19234
rect 5854 19070 5906 19122
rect 12686 19070 12738 19122
rect 14254 19070 14306 19122
rect 4734 18958 4786 19010
rect 13694 18958 13746 19010
rect 16382 19070 16434 19122
rect 16718 19070 16770 19122
rect 19518 19070 19570 19122
rect 22094 19070 22146 19122
rect 23774 19070 23826 19122
rect 32062 19070 32114 19122
rect 34862 19070 34914 19122
rect 35646 19070 35698 19122
rect 14030 18958 14082 19010
rect 14478 18958 14530 19010
rect 14590 18958 14642 19010
rect 15710 18958 15762 19010
rect 16942 18958 16994 19010
rect 21870 18958 21922 19010
rect 22990 18958 23042 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 2718 18622 2770 18674
rect 7646 18622 7698 18674
rect 10894 18622 10946 18674
rect 13022 18622 13074 18674
rect 17950 18622 18002 18674
rect 20638 18622 20690 18674
rect 21534 18622 21586 18674
rect 21982 18622 22034 18674
rect 22318 18622 22370 18674
rect 23102 18622 23154 18674
rect 34526 18622 34578 18674
rect 38334 18622 38386 18674
rect 2046 18510 2098 18562
rect 6302 18510 6354 18562
rect 7870 18510 7922 18562
rect 11454 18510 11506 18562
rect 13358 18510 13410 18562
rect 17502 18510 17554 18562
rect 21422 18510 21474 18562
rect 36094 18510 36146 18562
rect 1710 18398 1762 18450
rect 2382 18398 2434 18450
rect 3614 18398 3666 18450
rect 4510 18398 4562 18450
rect 5518 18398 5570 18450
rect 5742 18398 5794 18450
rect 6862 18398 6914 18450
rect 7198 18398 7250 18450
rect 9550 18398 9602 18450
rect 10110 18398 10162 18450
rect 11678 18398 11730 18450
rect 12350 18398 12402 18450
rect 12910 18398 12962 18450
rect 13694 18398 13746 18450
rect 14254 18398 14306 18450
rect 17390 18398 17442 18450
rect 18398 18398 18450 18450
rect 18958 18398 19010 18450
rect 19406 18398 19458 18450
rect 19630 18398 19682 18450
rect 20974 18398 21026 18450
rect 22766 18398 22818 18450
rect 23550 18398 23602 18450
rect 25342 18398 25394 18450
rect 26014 18398 26066 18450
rect 30830 18398 30882 18450
rect 31502 18398 31554 18450
rect 34974 18398 35026 18450
rect 35422 18398 35474 18450
rect 3166 18286 3218 18338
rect 4174 18286 4226 18338
rect 14702 18286 14754 18338
rect 16606 18286 16658 18338
rect 20302 18286 20354 18338
rect 28142 18286 28194 18338
rect 28702 18286 28754 18338
rect 32062 18286 32114 18338
rect 5406 18174 5458 18226
rect 14030 18174 14082 18226
rect 14478 18174 14530 18226
rect 14702 18174 14754 18226
rect 19294 18174 19346 18226
rect 21646 18174 21698 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 17838 17838 17890 17890
rect 1934 17726 1986 17778
rect 3166 17726 3218 17778
rect 3278 17726 3330 17778
rect 9662 17726 9714 17778
rect 14142 17726 14194 17778
rect 19294 17726 19346 17778
rect 21870 17726 21922 17778
rect 22990 17726 23042 17778
rect 25118 17726 25170 17778
rect 25566 17726 25618 17778
rect 28590 17726 28642 17778
rect 33742 17726 33794 17778
rect 34190 17726 34242 17778
rect 5070 17614 5122 17666
rect 5854 17614 5906 17666
rect 7870 17614 7922 17666
rect 8318 17614 8370 17666
rect 11454 17614 11506 17666
rect 17390 17614 17442 17666
rect 17726 17614 17778 17666
rect 17950 17614 18002 17666
rect 18510 17614 18562 17666
rect 22318 17614 22370 17666
rect 30830 17614 30882 17666
rect 2158 17502 2210 17554
rect 4510 17502 4562 17554
rect 6414 17502 6466 17554
rect 10110 17502 10162 17554
rect 11678 17502 11730 17554
rect 18846 17502 18898 17554
rect 31614 17502 31666 17554
rect 5854 17390 5906 17442
rect 13582 17390 13634 17442
rect 16606 17390 16658 17442
rect 18174 17390 18226 17442
rect 19742 17390 19794 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 3502 17054 3554 17106
rect 4062 17054 4114 17106
rect 4286 17054 4338 17106
rect 13694 17054 13746 17106
rect 16158 17054 16210 17106
rect 18734 17054 18786 17106
rect 22206 17054 22258 17106
rect 27358 17054 27410 17106
rect 27582 17054 27634 17106
rect 29262 17054 29314 17106
rect 33294 17054 33346 17106
rect 6078 16942 6130 16994
rect 6750 16942 6802 16994
rect 7534 16942 7586 16994
rect 13806 16942 13858 16994
rect 15934 16942 15986 16994
rect 17950 16942 18002 16994
rect 20974 16942 21026 16994
rect 21870 16942 21922 16994
rect 27918 16942 27970 16994
rect 2046 16830 2098 16882
rect 2606 16830 2658 16882
rect 2942 16830 2994 16882
rect 3838 16830 3890 16882
rect 4510 16830 4562 16882
rect 4846 16830 4898 16882
rect 6974 16830 7026 16882
rect 9886 16830 9938 16882
rect 10110 16830 10162 16882
rect 13022 16830 13074 16882
rect 14142 16830 14194 16882
rect 14926 16830 14978 16882
rect 15150 16830 15202 16882
rect 18174 16830 18226 16882
rect 20414 16830 20466 16882
rect 21646 16830 21698 16882
rect 29150 16830 29202 16882
rect 4622 16718 4674 16770
rect 9662 16718 9714 16770
rect 13358 16718 13410 16770
rect 16830 16718 16882 16770
rect 17614 16718 17666 16770
rect 22654 16718 22706 16770
rect 33070 16718 33122 16770
rect 33182 16718 33234 16770
rect 3166 16606 3218 16658
rect 10558 16606 10610 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 2158 16158 2210 16210
rect 4510 16158 4562 16210
rect 8318 16158 8370 16210
rect 11902 16158 11954 16210
rect 15486 16158 15538 16210
rect 17390 16158 17442 16210
rect 17726 16158 17778 16210
rect 18958 16158 19010 16210
rect 22094 16158 22146 16210
rect 28142 16158 28194 16210
rect 32846 16158 32898 16210
rect 35086 16158 35138 16210
rect 35646 16158 35698 16210
rect 3054 16046 3106 16098
rect 3278 16046 3330 16098
rect 3390 16046 3442 16098
rect 4734 16046 4786 16098
rect 5630 16046 5682 16098
rect 7646 16046 7698 16098
rect 10894 16046 10946 16098
rect 14142 16046 14194 16098
rect 14926 16046 14978 16098
rect 15150 16046 15202 16098
rect 16158 16046 16210 16098
rect 16830 16046 16882 16098
rect 17950 16046 18002 16098
rect 29486 16046 29538 16098
rect 29934 16046 29986 16098
rect 30270 16046 30322 16098
rect 32062 16046 32114 16098
rect 2942 15934 2994 15986
rect 5070 15934 5122 15986
rect 6750 15934 6802 15986
rect 8766 15934 8818 15986
rect 11118 15934 11170 15986
rect 11454 15934 11506 15986
rect 13918 15934 13970 15986
rect 15934 15934 15986 15986
rect 16606 15934 16658 15986
rect 19294 15934 19346 15986
rect 19406 15934 19458 15986
rect 29150 15934 29202 15986
rect 29262 15934 29314 15986
rect 29710 15934 29762 15986
rect 2606 15822 2658 15874
rect 18286 15822 18338 15874
rect 19630 15822 19682 15874
rect 26910 15822 26962 15874
rect 29934 15822 29986 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 3390 15486 3442 15538
rect 6302 15486 6354 15538
rect 8542 15486 8594 15538
rect 11454 15486 11506 15538
rect 11678 15486 11730 15538
rect 13134 15486 13186 15538
rect 16270 15486 16322 15538
rect 17502 15486 17554 15538
rect 17726 15486 17778 15538
rect 18510 15486 18562 15538
rect 20190 15486 20242 15538
rect 21534 15486 21586 15538
rect 22878 15486 22930 15538
rect 26350 15486 26402 15538
rect 28926 15486 28978 15538
rect 32398 15486 32450 15538
rect 4622 15374 4674 15426
rect 6638 15374 6690 15426
rect 15598 15374 15650 15426
rect 18062 15374 18114 15426
rect 20526 15374 20578 15426
rect 22094 15374 22146 15426
rect 25678 15374 25730 15426
rect 27582 15374 27634 15426
rect 28702 15374 28754 15426
rect 30158 15374 30210 15426
rect 1934 15262 1986 15314
rect 2382 15262 2434 15314
rect 2830 15262 2882 15314
rect 3950 15262 4002 15314
rect 6078 15262 6130 15314
rect 9774 15262 9826 15314
rect 11230 15262 11282 15314
rect 11342 15262 11394 15314
rect 11566 15262 11618 15314
rect 12462 15262 12514 15314
rect 15934 15262 15986 15314
rect 16606 15262 16658 15314
rect 17390 15262 17442 15314
rect 21646 15262 21698 15314
rect 22318 15262 22370 15314
rect 25902 15262 25954 15314
rect 26910 15262 26962 15314
rect 27358 15262 27410 15314
rect 28590 15262 28642 15314
rect 29374 15262 29426 15314
rect 8430 15150 8482 15202
rect 8766 15150 8818 15202
rect 9998 15150 10050 15202
rect 12686 15150 12738 15202
rect 15038 15150 15090 15202
rect 25342 15150 25394 15202
rect 27806 15150 27858 15202
rect 3054 15038 3106 15090
rect 10222 15038 10274 15090
rect 12126 15038 12178 15090
rect 21534 15038 21586 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 14702 14702 14754 14754
rect 16158 14702 16210 14754
rect 2494 14590 2546 14642
rect 3502 14590 3554 14642
rect 5070 14590 5122 14642
rect 7422 14590 7474 14642
rect 10894 14590 10946 14642
rect 24670 14590 24722 14642
rect 25230 14590 25282 14642
rect 29710 14590 29762 14642
rect 3166 14478 3218 14530
rect 5630 14478 5682 14530
rect 10446 14478 10498 14530
rect 13470 14478 13522 14530
rect 13918 14478 13970 14530
rect 14814 14478 14866 14530
rect 15262 14478 15314 14530
rect 15598 14478 15650 14530
rect 15822 14478 15874 14530
rect 16494 14478 16546 14530
rect 17166 14478 17218 14530
rect 21198 14478 21250 14530
rect 21534 14478 21586 14530
rect 22542 14478 22594 14530
rect 22878 14478 22930 14530
rect 23326 14478 23378 14530
rect 24222 14478 24274 14530
rect 26014 14478 26066 14530
rect 26574 14478 26626 14530
rect 6638 14366 6690 14418
rect 11790 14366 11842 14418
rect 11902 14366 11954 14418
rect 14254 14366 14306 14418
rect 14702 14366 14754 14418
rect 16830 14366 16882 14418
rect 17278 14366 17330 14418
rect 21870 14366 21922 14418
rect 23102 14366 23154 14418
rect 23662 14366 23714 14418
rect 23886 14366 23938 14418
rect 26686 14366 26738 14418
rect 26910 14366 26962 14418
rect 27134 14366 27186 14418
rect 27358 14366 27410 14418
rect 27694 14366 27746 14418
rect 27918 14366 27970 14418
rect 28254 14366 28306 14418
rect 1934 14254 1986 14306
rect 4510 14254 4562 14306
rect 7086 14254 7138 14306
rect 9998 14254 10050 14306
rect 11566 14254 11618 14306
rect 12350 14254 12402 14306
rect 17502 14254 17554 14306
rect 21422 14254 21474 14306
rect 22654 14254 22706 14306
rect 23438 14254 23490 14306
rect 24110 14254 24162 14306
rect 25678 14254 25730 14306
rect 26126 14254 26178 14306
rect 26350 14254 26402 14306
rect 27582 14254 27634 14306
rect 28142 14254 28194 14306
rect 29262 14254 29314 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 1710 13918 1762 13970
rect 2718 13918 2770 13970
rect 11902 13918 11954 13970
rect 14590 13918 14642 13970
rect 19070 13918 19122 13970
rect 42814 13918 42866 13970
rect 3614 13806 3666 13858
rect 7422 13806 7474 13858
rect 7758 13806 7810 13858
rect 17726 13806 17778 13858
rect 18062 13806 18114 13858
rect 21310 13806 21362 13858
rect 22542 13806 22594 13858
rect 26014 13806 26066 13858
rect 26350 13806 26402 13858
rect 26462 13806 26514 13858
rect 27694 13806 27746 13858
rect 2270 13694 2322 13746
rect 3054 13694 3106 13746
rect 6414 13694 6466 13746
rect 7086 13694 7138 13746
rect 7534 13694 7586 13746
rect 11006 13694 11058 13746
rect 18622 13694 18674 13746
rect 22094 13694 22146 13746
rect 26686 13694 26738 13746
rect 27022 13694 27074 13746
rect 43150 13694 43202 13746
rect 3950 13582 4002 13634
rect 4174 13582 4226 13634
rect 11230 13582 11282 13634
rect 15262 13582 15314 13634
rect 16606 13582 16658 13634
rect 29822 13582 29874 13634
rect 42590 13582 42642 13634
rect 10782 13470 10834 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 17390 13134 17442 13186
rect 2158 13022 2210 13074
rect 3166 13022 3218 13074
rect 3838 13022 3890 13074
rect 5854 13022 5906 13074
rect 19742 13134 19794 13186
rect 6638 13022 6690 13074
rect 14142 13022 14194 13074
rect 17726 13022 17778 13074
rect 18510 13022 18562 13074
rect 19294 13022 19346 13074
rect 19742 13022 19794 13074
rect 20750 13022 20802 13074
rect 21758 13022 21810 13074
rect 23326 13022 23378 13074
rect 25454 13022 25506 13074
rect 1822 12910 1874 12962
rect 2718 12910 2770 12962
rect 14254 12910 14306 12962
rect 18846 12910 18898 12962
rect 21310 12910 21362 12962
rect 22654 12910 22706 12962
rect 27246 12910 27298 12962
rect 27470 12910 27522 12962
rect 27806 12910 27858 12962
rect 3502 12798 3554 12850
rect 13694 12798 13746 12850
rect 15038 12798 15090 12850
rect 17614 12798 17666 12850
rect 19182 12798 19234 12850
rect 7086 12686 7138 12738
rect 10334 12686 10386 12738
rect 17054 12686 17106 12738
rect 27470 12686 27522 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 2718 12350 2770 12402
rect 4398 12350 4450 12402
rect 5406 12350 5458 12402
rect 5742 12350 5794 12402
rect 6302 12350 6354 12402
rect 7086 12350 7138 12402
rect 7758 12350 7810 12402
rect 10334 12350 10386 12402
rect 10558 12350 10610 12402
rect 11230 12350 11282 12402
rect 14702 12350 14754 12402
rect 18622 12350 18674 12402
rect 26350 12350 26402 12402
rect 5854 12238 5906 12290
rect 6190 12238 6242 12290
rect 8878 12238 8930 12290
rect 9886 12238 9938 12290
rect 16718 12238 16770 12290
rect 29374 12238 29426 12290
rect 1710 12126 1762 12178
rect 2270 12126 2322 12178
rect 5518 12126 5570 12178
rect 7198 12126 7250 12178
rect 8766 12126 8818 12178
rect 9102 12126 9154 12178
rect 9438 12126 9490 12178
rect 10110 12126 10162 12178
rect 10670 12126 10722 12178
rect 13694 12126 13746 12178
rect 13918 12126 13970 12178
rect 16830 12126 16882 12178
rect 17614 12126 17666 12178
rect 17726 12126 17778 12178
rect 17838 12126 17890 12178
rect 18174 12126 18226 12178
rect 27134 12126 27186 12178
rect 3166 12014 3218 12066
rect 4958 12014 5010 12066
rect 9662 12014 9714 12066
rect 18062 12014 18114 12066
rect 6302 11902 6354 11954
rect 7086 11902 7138 11954
rect 13582 11902 13634 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 1822 11454 1874 11506
rect 5070 11454 5122 11506
rect 6750 11454 6802 11506
rect 8318 11454 8370 11506
rect 10446 11454 10498 11506
rect 2270 11342 2322 11394
rect 5630 11342 5682 11394
rect 6078 11342 6130 11394
rect 7086 11342 7138 11394
rect 7534 11342 7586 11394
rect 11230 11342 11282 11394
rect 11678 11342 11730 11394
rect 18734 11342 18786 11394
rect 2942 11230 2994 11282
rect 6302 11230 6354 11282
rect 10894 11230 10946 11282
rect 11902 11230 11954 11282
rect 12238 11230 12290 11282
rect 12350 11230 12402 11282
rect 13694 11230 13746 11282
rect 22318 11230 22370 11282
rect 22430 11230 22482 11282
rect 22990 11230 23042 11282
rect 5854 11118 5906 11170
rect 12574 11118 12626 11170
rect 19182 11118 19234 11170
rect 22654 11118 22706 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 5518 10782 5570 10834
rect 5742 10782 5794 10834
rect 6302 10782 6354 10834
rect 7198 10782 7250 10834
rect 7758 10782 7810 10834
rect 10670 10782 10722 10834
rect 14478 10782 14530 10834
rect 15374 10782 15426 10834
rect 17390 10782 17442 10834
rect 22206 10782 22258 10834
rect 23998 10782 24050 10834
rect 30158 10782 30210 10834
rect 2942 10670 2994 10722
rect 5854 10670 5906 10722
rect 7310 10670 7362 10722
rect 15262 10670 15314 10722
rect 19742 10670 19794 10722
rect 21646 10670 21698 10722
rect 22094 10670 22146 10722
rect 27918 10670 27970 10722
rect 2270 10558 2322 10610
rect 6190 10558 6242 10610
rect 6526 10558 6578 10610
rect 6750 10558 6802 10610
rect 6974 10558 7026 10610
rect 11118 10558 11170 10610
rect 15598 10558 15650 10610
rect 15822 10558 15874 10610
rect 16382 10558 16434 10610
rect 17614 10558 17666 10610
rect 19406 10558 19458 10610
rect 21534 10558 21586 10610
rect 21870 10558 21922 10610
rect 22878 10558 22930 10610
rect 23102 10558 23154 10610
rect 23438 10558 23490 10610
rect 27246 10558 27298 10610
rect 1822 10446 1874 10498
rect 5070 10446 5122 10498
rect 11902 10446 11954 10498
rect 14030 10446 14082 10498
rect 15038 10446 15090 10498
rect 20302 10446 20354 10498
rect 20750 10446 20802 10498
rect 21198 10446 21250 10498
rect 22990 10446 23042 10498
rect 20302 10334 20354 10386
rect 21310 10334 21362 10386
rect 22206 10334 22258 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 12798 9998 12850 10050
rect 2270 9886 2322 9938
rect 5070 9886 5122 9938
rect 5854 9886 5906 9938
rect 6974 9886 7026 9938
rect 7422 9886 7474 9938
rect 12238 9886 12290 9938
rect 13582 9886 13634 9938
rect 15150 9886 15202 9938
rect 15934 9886 15986 9938
rect 18062 9886 18114 9938
rect 26126 9886 26178 9938
rect 27918 9886 27970 9938
rect 30718 9886 30770 9938
rect 6190 9774 6242 9826
rect 6526 9774 6578 9826
rect 11454 9774 11506 9826
rect 12126 9774 12178 9826
rect 12462 9774 12514 9826
rect 12686 9774 12738 9826
rect 18734 9774 18786 9826
rect 20526 9774 20578 9826
rect 22094 9774 22146 9826
rect 22542 9774 22594 9826
rect 23326 9774 23378 9826
rect 29262 9774 29314 9826
rect 1710 9662 1762 9714
rect 11790 9662 11842 9714
rect 21422 9662 21474 9714
rect 6414 9550 6466 9602
rect 11118 9550 11170 9602
rect 12798 9550 12850 9602
rect 14702 9550 14754 9602
rect 19742 9550 19794 9602
rect 20190 9550 20242 9602
rect 20638 9550 20690 9602
rect 20862 9550 20914 9602
rect 21758 9606 21810 9658
rect 21870 9662 21922 9714
rect 22318 9662 22370 9714
rect 22766 9662 22818 9714
rect 22878 9662 22930 9714
rect 23998 9662 24050 9714
rect 28142 9662 28194 9714
rect 28254 9662 28306 9714
rect 29598 9662 29650 9714
rect 29710 9662 29762 9714
rect 28478 9550 28530 9602
rect 29934 9550 29986 9602
rect 30270 9550 30322 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 2046 9214 2098 9266
rect 6078 9214 6130 9266
rect 15374 9214 15426 9266
rect 16158 9214 16210 9266
rect 23998 9214 24050 9266
rect 10558 9102 10610 9154
rect 10670 9102 10722 9154
rect 11230 9102 11282 9154
rect 15822 9102 15874 9154
rect 16718 9102 16770 9154
rect 18734 9102 18786 9154
rect 22990 9102 23042 9154
rect 29262 9102 29314 9154
rect 1710 8990 1762 9042
rect 9550 8990 9602 9042
rect 9998 8990 10050 9042
rect 10334 8990 10386 9042
rect 11454 8990 11506 9042
rect 16270 8990 16322 9042
rect 16606 8990 16658 9042
rect 16942 8990 16994 9042
rect 22654 8990 22706 9042
rect 23214 8990 23266 9042
rect 23438 8990 23490 9042
rect 25342 8990 25394 9042
rect 28590 8990 28642 9042
rect 2494 8878 2546 8930
rect 12014 8878 12066 8930
rect 23102 8878 23154 8930
rect 26014 8878 26066 8930
rect 28142 8878 28194 8930
rect 31390 8878 31442 8930
rect 16158 8766 16210 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 15822 8318 15874 8370
rect 16270 8318 16322 8370
rect 23550 8318 23602 8370
rect 9998 8206 10050 8258
rect 11566 8206 11618 8258
rect 12910 8206 12962 8258
rect 13470 8206 13522 8258
rect 17390 8206 17442 8258
rect 17838 8206 17890 8258
rect 18510 8206 18562 8258
rect 19294 8206 19346 8258
rect 19854 8206 19906 8258
rect 20190 8206 20242 8258
rect 21310 8206 21362 8258
rect 21758 8206 21810 8258
rect 21870 8206 21922 8258
rect 22318 8206 22370 8258
rect 22654 8206 22706 8258
rect 23214 8206 23266 8258
rect 9774 8094 9826 8146
rect 10334 8094 10386 8146
rect 10670 8094 10722 8146
rect 12350 8094 12402 8146
rect 12798 8094 12850 8146
rect 16606 8094 16658 8146
rect 16718 8094 16770 8146
rect 17166 8094 17218 8146
rect 18734 8094 18786 8146
rect 19182 8094 19234 8146
rect 20414 8094 20466 8146
rect 20750 8094 20802 8146
rect 22430 8094 22482 8146
rect 22878 8094 22930 8146
rect 22990 8094 23042 8146
rect 9886 7982 9938 8034
rect 11006 7982 11058 8034
rect 11230 7982 11282 8034
rect 11454 7982 11506 8034
rect 12574 7982 12626 8034
rect 13582 7982 13634 8034
rect 13806 7982 13858 8034
rect 14142 7982 14194 8034
rect 16942 7982 16994 8034
rect 17614 7982 17666 8034
rect 18958 7982 19010 8034
rect 19966 7982 20018 8034
rect 21534 7982 21586 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 2046 7646 2098 7698
rect 10222 7646 10274 7698
rect 10446 7646 10498 7698
rect 13022 7646 13074 7698
rect 15374 7646 15426 7698
rect 15822 7646 15874 7698
rect 19070 7646 19122 7698
rect 19294 7646 19346 7698
rect 20302 7646 20354 7698
rect 21422 7646 21474 7698
rect 10558 7534 10610 7586
rect 12014 7534 12066 7586
rect 12910 7534 12962 7586
rect 15934 7534 15986 7586
rect 17390 7534 17442 7586
rect 17726 7534 17778 7586
rect 18062 7534 18114 7586
rect 18622 7534 18674 7586
rect 19966 7534 20018 7586
rect 20638 7534 20690 7586
rect 21646 7590 21698 7642
rect 21758 7646 21810 7698
rect 21982 7646 22034 7698
rect 22654 7646 22706 7698
rect 22990 7646 23042 7698
rect 1710 7422 1762 7474
rect 12350 7422 12402 7474
rect 12686 7422 12738 7474
rect 16158 7422 16210 7474
rect 16494 7422 16546 7474
rect 16830 7422 16882 7474
rect 18398 7422 18450 7474
rect 18958 7422 19010 7474
rect 2494 7310 2546 7362
rect 11006 7310 11058 7362
rect 12462 7310 12514 7362
rect 16382 7310 16434 7362
rect 18510 7310 18562 7362
rect 13022 7198 13074 7250
rect 15822 7198 15874 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 9998 6750 10050 6802
rect 15822 6750 15874 6802
rect 17950 6750 18002 6802
rect 19630 6750 19682 6802
rect 19966 6750 20018 6802
rect 7086 6638 7138 6690
rect 7870 6638 7922 6690
rect 10334 6638 10386 6690
rect 10670 6638 10722 6690
rect 11454 6638 11506 6690
rect 11902 6638 11954 6690
rect 12686 6638 12738 6690
rect 13022 6638 13074 6690
rect 13470 6638 13522 6690
rect 13806 6638 13858 6690
rect 14142 6638 14194 6690
rect 15150 6638 15202 6690
rect 10894 6526 10946 6578
rect 11118 6526 11170 6578
rect 12798 6526 12850 6578
rect 10670 6414 10722 6466
rect 11342 6414 11394 6466
rect 13806 6414 13858 6466
rect 18846 6414 18898 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 10222 6078 10274 6130
rect 14254 6078 14306 6130
rect 24334 6078 24386 6130
rect 2046 5966 2098 6018
rect 11678 5966 11730 6018
rect 22094 5966 22146 6018
rect 1710 5854 1762 5906
rect 10894 5854 10946 5906
rect 17502 5854 17554 5906
rect 21310 5854 21362 5906
rect 2494 5742 2546 5794
rect 13806 5742 13858 5794
rect 18398 5630 18450 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 8878 5182 8930 5234
rect 11006 5182 11058 5234
rect 11902 5182 11954 5234
rect 12686 5182 12738 5234
rect 13470 5182 13522 5234
rect 15598 5182 15650 5234
rect 18622 5182 18674 5234
rect 20750 5182 20802 5234
rect 1710 5070 1762 5122
rect 2494 5070 2546 5122
rect 8094 5070 8146 5122
rect 11790 5070 11842 5122
rect 16382 5070 16434 5122
rect 17838 5070 17890 5122
rect 42590 5070 42642 5122
rect 43150 5070 43202 5122
rect 2046 4958 2098 5010
rect 12126 4958 12178 5010
rect 42814 4958 42866 5010
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 10558 4510 10610 4562
rect 23886 4510 23938 4562
rect 36654 4510 36706 4562
rect 18174 4398 18226 4450
rect 1822 4286 1874 4338
rect 6078 4286 6130 4338
rect 6414 4286 6466 4338
rect 10110 4286 10162 4338
rect 12910 4286 12962 4338
rect 14142 4286 14194 4338
rect 17502 4286 17554 4338
rect 22990 4286 23042 4338
rect 28814 4286 28866 4338
rect 29934 4286 29986 4338
rect 36990 4286 37042 4338
rect 42366 4286 42418 4338
rect 2158 4174 2210 4226
rect 11678 4174 11730 4226
rect 20302 4174 20354 4226
rect 33294 4174 33346 4226
rect 42142 4174 42194 4226
rect 42814 4174 42866 4226
rect 4174 4062 4226 4114
rect 7422 4062 7474 4114
rect 14702 4062 14754 4114
rect 21086 4062 21138 4114
rect 26462 4062 26514 4114
rect 30830 4062 30882 4114
rect 37998 4062 38050 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 2718 3614 2770 3666
rect 10222 3614 10274 3666
rect 18846 3614 18898 3666
rect 24782 3614 24834 3666
rect 27582 3614 27634 3666
rect 29374 3614 29426 3666
rect 32734 3614 32786 3666
rect 35534 3614 35586 3666
rect 36990 3614 37042 3666
rect 39342 3614 39394 3666
rect 40798 3614 40850 3666
rect 4846 3502 4898 3554
rect 8766 3502 8818 3554
rect 12126 3502 12178 3554
rect 15934 3502 15986 3554
rect 19742 3502 19794 3554
rect 21422 3502 21474 3554
rect 27134 3502 27186 3554
rect 28478 3502 28530 3554
rect 33630 3502 33682 3554
rect 35982 3502 36034 3554
rect 39790 3502 39842 3554
rect 1822 3390 1874 3442
rect 31726 3390 31778 3442
rect 32174 3390 32226 3442
rect 33406 3390 33458 3442
rect 7758 3278 7810 3330
rect 15374 3278 15426 3330
rect 22430 3278 22482 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 3808 44200 3920 45000
rect 4928 44200 5040 45000
rect 6048 44200 6160 45000
rect 7168 44200 7280 45000
rect 8288 44200 8400 45000
rect 9408 44200 9520 45000
rect 10528 44200 10640 45000
rect 11648 44200 11760 45000
rect 12768 44200 12880 45000
rect 13888 44200 14000 45000
rect 15008 44200 15120 45000
rect 16128 44200 16240 45000
rect 17248 44200 17360 45000
rect 18368 44200 18480 45000
rect 19488 44200 19600 45000
rect 20608 44200 20720 45000
rect 21728 44200 21840 45000
rect 22848 44200 22960 45000
rect 23968 44200 24080 45000
rect 25088 44200 25200 45000
rect 26208 44200 26320 45000
rect 27328 44200 27440 45000
rect 28448 44200 28560 45000
rect 29568 44200 29680 45000
rect 30688 44200 30800 45000
rect 31808 44200 31920 45000
rect 32928 44200 33040 45000
rect 34048 44200 34160 45000
rect 35168 44200 35280 45000
rect 36288 44200 36400 45000
rect 37408 44200 37520 45000
rect 38528 44200 38640 45000
rect 39648 44200 39760 45000
rect 40768 44200 40880 45000
rect 41132 44268 41636 44324
rect 1932 41298 1988 41310
rect 1932 41246 1934 41298
rect 1986 41246 1988 41298
rect 1932 40628 1988 41246
rect 1932 40562 1988 40572
rect 1932 40178 1988 40190
rect 1932 40126 1934 40178
rect 1986 40126 1988 40178
rect 1820 39618 1876 39630
rect 1820 39566 1822 39618
rect 1874 39566 1876 39618
rect 1820 38836 1876 39566
rect 1932 39620 1988 40126
rect 3836 39732 3892 44200
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4732 41300 4788 41310
rect 4284 41186 4340 41198
rect 4284 41134 4286 41186
rect 4338 41134 4340 41186
rect 4284 41076 4340 41134
rect 4732 41186 4788 41244
rect 4956 41188 5012 44200
rect 6076 42084 6132 44200
rect 5628 42028 6132 42084
rect 4732 41134 4734 41186
rect 4786 41134 4788 41186
rect 4732 41122 4788 41134
rect 4844 41132 5012 41188
rect 5404 41972 5460 41982
rect 4284 41010 4340 41020
rect 4396 40964 4452 40974
rect 3836 39666 3892 39676
rect 4172 40740 4228 40750
rect 1932 39554 1988 39564
rect 2492 39506 2548 39518
rect 2492 39454 2494 39506
rect 2546 39454 2548 39506
rect 1932 38836 1988 38846
rect 1820 38780 1932 38836
rect 1372 38724 1428 38734
rect 1260 30100 1316 30110
rect 1260 13076 1316 30044
rect 1372 21924 1428 38668
rect 1820 35698 1876 38780
rect 1932 38742 1988 38780
rect 1932 38164 1988 38174
rect 1932 38070 1988 38108
rect 1932 37042 1988 37054
rect 1932 36990 1934 37042
rect 1986 36990 1988 37042
rect 1932 36596 1988 36990
rect 2492 36932 2548 39454
rect 4172 39172 4228 40684
rect 4284 40404 4340 40414
rect 4396 40404 4452 40908
rect 4284 40402 4452 40404
rect 4284 40350 4286 40402
rect 4338 40350 4452 40402
rect 4284 40348 4452 40350
rect 4284 40338 4340 40348
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4620 39730 4676 39742
rect 4620 39678 4622 39730
rect 4674 39678 4676 39730
rect 4620 39172 4676 39678
rect 4172 39116 4676 39172
rect 2604 38724 2660 38734
rect 2604 38722 2996 38724
rect 2604 38670 2606 38722
rect 2658 38670 2996 38722
rect 2604 38668 2996 38670
rect 2604 38658 2660 38668
rect 2492 36876 2884 36932
rect 1932 36530 1988 36540
rect 2044 36594 2100 36606
rect 2044 36542 2046 36594
rect 2098 36542 2100 36594
rect 1820 35646 1822 35698
rect 1874 35646 1876 35698
rect 1820 35634 1876 35646
rect 1596 35588 1652 35598
rect 1484 35028 1540 35038
rect 1484 29652 1540 34972
rect 1484 29586 1540 29596
rect 1372 21858 1428 21868
rect 1260 13010 1316 13020
rect 1596 11620 1652 35532
rect 2044 35252 2100 36542
rect 2492 35588 2548 35598
rect 2044 35186 2100 35196
rect 2380 35586 2548 35588
rect 2380 35534 2494 35586
rect 2546 35534 2548 35586
rect 2380 35532 2548 35534
rect 1932 35026 1988 35038
rect 1932 34974 1934 35026
rect 1986 34974 1988 35026
rect 1932 33908 1988 34974
rect 2044 34804 2100 34814
rect 2044 34242 2100 34748
rect 2044 34190 2046 34242
rect 2098 34190 2100 34242
rect 2044 34178 2100 34190
rect 2156 34132 2212 34142
rect 2156 34038 2212 34076
rect 1932 33842 1988 33852
rect 2268 33908 2324 33918
rect 1932 33458 1988 33470
rect 1932 33406 1934 33458
rect 1986 33406 1988 33458
rect 1932 32564 1988 33406
rect 2044 33460 2100 33470
rect 2044 32674 2100 33404
rect 2044 32622 2046 32674
rect 2098 32622 2100 32674
rect 2044 32610 2100 32622
rect 2268 32674 2324 33852
rect 2380 32786 2436 35532
rect 2492 35522 2548 35532
rect 2828 34354 2884 36876
rect 2940 36596 2996 38668
rect 2940 36530 2996 36540
rect 4060 37828 4116 37838
rect 4060 36482 4116 37772
rect 4060 36430 4062 36482
rect 4114 36430 4116 36482
rect 4060 36418 4116 36430
rect 4172 36148 4228 39116
rect 4284 38948 4340 38958
rect 4284 38050 4340 38892
rect 4732 38722 4788 38734
rect 4732 38670 4734 38722
rect 4786 38670 4788 38722
rect 4732 38612 4788 38670
rect 4732 38546 4788 38556
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4284 37998 4286 38050
rect 4338 37998 4340 38050
rect 4284 37986 4340 37998
rect 4844 38052 4900 41132
rect 4956 40962 5012 40974
rect 4956 40910 4958 40962
rect 5010 40910 5012 40962
rect 4956 40404 5012 40910
rect 5404 40514 5460 41916
rect 5628 41300 5684 42028
rect 7196 41412 7252 44200
rect 7196 41356 7588 41412
rect 5628 41206 5684 41244
rect 5404 40462 5406 40514
rect 5458 40462 5460 40514
rect 5404 40450 5460 40462
rect 7532 40514 7588 41356
rect 7868 41186 7924 41198
rect 7868 41134 7870 41186
rect 7922 41134 7924 41186
rect 7644 40964 7700 40974
rect 7644 40870 7700 40908
rect 7868 40740 7924 41134
rect 8204 40740 8260 40750
rect 7868 40674 7924 40684
rect 8092 40684 8204 40740
rect 7532 40462 7534 40514
rect 7586 40462 7588 40514
rect 4956 40338 5012 40348
rect 5964 40404 6020 40414
rect 5068 39394 5124 39406
rect 5068 39342 5070 39394
rect 5122 39342 5124 39394
rect 5068 38836 5124 39342
rect 5740 39394 5796 39406
rect 5740 39342 5742 39394
rect 5794 39342 5796 39394
rect 5180 38836 5236 38846
rect 5068 38780 5180 38836
rect 5180 38742 5236 38780
rect 5740 38836 5796 39342
rect 5740 38770 5796 38780
rect 5852 38722 5908 38734
rect 5852 38670 5854 38722
rect 5906 38670 5908 38722
rect 4844 37958 4900 37996
rect 5740 38052 5796 38062
rect 5740 37958 5796 37996
rect 5068 37828 5124 37838
rect 5068 37826 5236 37828
rect 5068 37774 5070 37826
rect 5122 37774 5236 37826
rect 5068 37772 5236 37774
rect 5068 37762 5124 37772
rect 4284 37380 4340 37390
rect 4284 37266 4340 37324
rect 4956 37268 5012 37278
rect 4284 37214 4286 37266
rect 4338 37214 4340 37266
rect 4284 37202 4340 37214
rect 4844 37212 4956 37268
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4844 36708 4900 37212
rect 4956 37202 5012 37212
rect 4060 36092 4228 36148
rect 4620 36652 4900 36708
rect 5068 36932 5124 36942
rect 4060 34804 4116 36092
rect 4620 35588 4676 36652
rect 4284 35586 4676 35588
rect 4284 35534 4622 35586
rect 4674 35534 4676 35586
rect 4284 35532 4676 35534
rect 4284 35140 4340 35532
rect 4620 35522 4676 35532
rect 4844 36482 4900 36494
rect 4844 36430 4846 36482
rect 4898 36430 4900 36482
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4060 34738 4116 34748
rect 4172 35084 4788 35140
rect 2828 34302 2830 34354
rect 2882 34302 2884 34354
rect 2828 34290 2884 34302
rect 2716 34242 2772 34254
rect 2716 34190 2718 34242
rect 2770 34190 2772 34242
rect 2492 34130 2548 34142
rect 2492 34078 2494 34130
rect 2546 34078 2548 34130
rect 2492 33460 2548 34078
rect 2604 34132 2660 34142
rect 2716 34132 2772 34190
rect 2660 34076 2772 34132
rect 3276 34130 3332 34142
rect 3276 34078 3278 34130
rect 3330 34078 3332 34130
rect 2604 34066 2660 34076
rect 3052 33906 3108 33918
rect 3052 33854 3054 33906
rect 3106 33854 3108 33906
rect 2548 33404 2660 33460
rect 2492 33394 2548 33404
rect 2380 32734 2382 32786
rect 2434 32734 2436 32786
rect 2380 32722 2436 32734
rect 2268 32622 2270 32674
rect 2322 32622 2324 32674
rect 2268 32610 2324 32622
rect 1932 32498 1988 32508
rect 2492 32338 2548 32350
rect 2492 32286 2494 32338
rect 2546 32286 2548 32338
rect 1932 31890 1988 31902
rect 1932 31838 1934 31890
rect 1986 31838 1988 31890
rect 1932 31220 1988 31838
rect 1932 31154 1988 31164
rect 1820 30882 1876 30894
rect 1820 30830 1822 30882
rect 1874 30830 1876 30882
rect 1820 29876 1876 30830
rect 2380 30882 2436 30894
rect 2380 30830 2382 30882
rect 2434 30830 2436 30882
rect 1932 30324 1988 30334
rect 1932 30230 1988 30268
rect 1820 29426 1876 29820
rect 2044 29652 2100 29662
rect 2044 29558 2100 29596
rect 2380 29540 2436 30830
rect 2492 29988 2548 32286
rect 2604 31948 2660 33404
rect 3052 33012 3108 33854
rect 3052 32946 3108 32956
rect 2828 32562 2884 32574
rect 2828 32510 2830 32562
rect 2882 32510 2884 32562
rect 2828 32452 2884 32510
rect 3276 32452 3332 34078
rect 3612 34018 3668 34030
rect 3612 33966 3614 34018
rect 3666 33966 3668 34018
rect 3612 32900 3668 33966
rect 3612 32834 3668 32844
rect 4172 32676 4228 35084
rect 4732 35026 4788 35084
rect 4732 34974 4734 35026
rect 4786 34974 4788 35026
rect 4732 34962 4788 34974
rect 4284 34914 4340 34926
rect 4284 34862 4286 34914
rect 4338 34862 4340 34914
rect 4284 33572 4340 34862
rect 4620 34690 4676 34702
rect 4620 34638 4622 34690
rect 4674 34638 4676 34690
rect 4620 33908 4676 34638
rect 4620 33842 4676 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4284 33506 4340 33516
rect 4284 33346 4340 33358
rect 4284 33294 4286 33346
rect 4338 33294 4340 33346
rect 4284 33236 4340 33294
rect 4620 33348 4676 33358
rect 4620 33254 4676 33292
rect 4284 33170 4340 33180
rect 4732 33122 4788 33134
rect 4732 33070 4734 33122
rect 4786 33070 4788 33122
rect 4732 32900 4788 33070
rect 4732 32834 4788 32844
rect 4172 32610 4228 32620
rect 3724 32452 3780 32462
rect 2828 32450 3780 32452
rect 2828 32398 3278 32450
rect 3330 32398 3726 32450
rect 3778 32398 3780 32450
rect 2828 32396 3780 32398
rect 3276 32386 3332 32396
rect 2604 31892 2996 31948
rect 2604 31444 2660 31454
rect 2604 31106 2660 31388
rect 2604 31054 2606 31106
rect 2658 31054 2660 31106
rect 2604 30324 2660 31054
rect 2940 31108 2996 31892
rect 3052 31108 3108 31118
rect 2940 31106 3108 31108
rect 2940 31054 3054 31106
rect 3106 31054 3108 31106
rect 2940 31052 3108 31054
rect 2716 30772 2772 30782
rect 2716 30770 2996 30772
rect 2716 30718 2718 30770
rect 2770 30718 2996 30770
rect 2716 30716 2996 30718
rect 2716 30706 2772 30716
rect 2604 30258 2660 30268
rect 2492 29932 2660 29988
rect 2604 29650 2660 29932
rect 2604 29598 2606 29650
rect 2658 29598 2660 29650
rect 2604 29586 2660 29598
rect 2716 29652 2772 29662
rect 2492 29540 2548 29550
rect 2380 29538 2548 29540
rect 2380 29486 2494 29538
rect 2546 29486 2548 29538
rect 2380 29484 2548 29486
rect 1820 29374 1822 29426
rect 1874 29374 1876 29426
rect 1820 29362 1876 29374
rect 1932 28754 1988 28766
rect 1932 28702 1934 28754
rect 1986 28702 1988 28754
rect 1932 28532 1988 28702
rect 1932 28466 1988 28476
rect 1932 27634 1988 27646
rect 1932 27582 1934 27634
rect 1986 27582 1988 27634
rect 1932 27188 1988 27582
rect 1932 27122 1988 27132
rect 2044 27186 2100 27198
rect 2044 27134 2046 27186
rect 2098 27134 2100 27186
rect 2044 25844 2100 27134
rect 2044 25778 2100 25788
rect 1708 25620 1764 25630
rect 1708 25526 1764 25564
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 1708 24050 1764 24062
rect 1708 23998 1710 24050
rect 1762 23998 1764 24050
rect 1708 23604 1764 23998
rect 1708 23538 1764 23548
rect 1932 23156 1988 23166
rect 1932 22594 1988 23100
rect 1932 22542 1934 22594
rect 1986 22542 1988 22594
rect 1932 22530 1988 22542
rect 1932 21812 1988 21822
rect 1932 21474 1988 21756
rect 1932 21422 1934 21474
rect 1986 21422 1988 21474
rect 1932 21410 1988 21422
rect 1708 21028 1764 21038
rect 1708 20914 1764 20972
rect 1708 20862 1710 20914
rect 1762 20862 1764 20914
rect 1708 20850 1764 20862
rect 1932 20468 1988 20478
rect 1932 19906 1988 20412
rect 1932 19854 1934 19906
rect 1986 19854 1988 19906
rect 1932 19842 1988 19854
rect 1932 19348 1988 19358
rect 1932 19254 1988 19292
rect 2044 18562 2100 18574
rect 2044 18510 2046 18562
rect 2098 18510 2100 18562
rect 1708 18452 1764 18462
rect 1708 17780 1764 18396
rect 2044 18228 2100 18510
rect 2044 18162 2100 18172
rect 2380 18450 2436 18462
rect 2380 18398 2382 18450
rect 2434 18398 2436 18450
rect 2380 18340 2436 18398
rect 1708 17714 1764 17724
rect 1932 17780 1988 17790
rect 1932 17686 1988 17724
rect 2156 17556 2212 17566
rect 1932 17554 2212 17556
rect 1932 17502 2158 17554
rect 2210 17502 2212 17554
rect 1932 17500 2212 17502
rect 1932 16100 1988 17500
rect 2156 17490 2212 17500
rect 2268 17556 2324 17566
rect 2268 17108 2324 17500
rect 2044 17052 2324 17108
rect 2044 16882 2100 17052
rect 2044 16830 2046 16882
rect 2098 16830 2100 16882
rect 2044 16818 2100 16830
rect 2268 16884 2324 16894
rect 2156 16772 2212 16782
rect 2156 16210 2212 16716
rect 2156 16158 2158 16210
rect 2210 16158 2212 16210
rect 2156 16146 2212 16158
rect 1932 16034 1988 16044
rect 1932 15314 1988 15326
rect 1932 15262 1934 15314
rect 1986 15262 1988 15314
rect 1708 15092 1764 15102
rect 1708 13972 1764 15036
rect 1708 13878 1764 13916
rect 1932 15092 1988 15262
rect 2268 15316 2324 16828
rect 2380 16436 2436 18284
rect 2380 16370 2436 16380
rect 2380 15316 2436 15326
rect 2268 15314 2436 15316
rect 2268 15262 2382 15314
rect 2434 15262 2436 15314
rect 2268 15260 2436 15262
rect 2380 15250 2436 15260
rect 1932 14306 1988 15036
rect 2492 14868 2548 29484
rect 2716 29538 2772 29596
rect 2716 29486 2718 29538
rect 2770 29486 2772 29538
rect 2716 29474 2772 29486
rect 2940 29316 2996 30716
rect 3052 29538 3108 31052
rect 3276 30994 3332 31006
rect 3276 30942 3278 30994
rect 3330 30942 3332 30994
rect 3276 29652 3332 30942
rect 3276 29586 3332 29596
rect 3052 29486 3054 29538
rect 3106 29486 3108 29538
rect 3052 29474 3108 29486
rect 3276 29426 3332 29438
rect 3276 29374 3278 29426
rect 3330 29374 3332 29426
rect 3276 29316 3332 29374
rect 2940 29260 3332 29316
rect 3052 27300 3108 27310
rect 2716 21812 2772 21822
rect 2716 18674 2772 21756
rect 2716 18622 2718 18674
rect 2770 18622 2772 18674
rect 2716 18610 2772 18622
rect 3052 17780 3108 27244
rect 3500 23548 3556 32396
rect 3724 32386 3780 32396
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4060 31778 4116 31790
rect 4060 31726 4062 31778
rect 4114 31726 4116 31778
rect 4060 31218 4116 31726
rect 4844 31668 4900 36430
rect 5068 36372 5124 36876
rect 4956 36370 5124 36372
rect 4956 36318 5070 36370
rect 5122 36318 5124 36370
rect 4956 36316 5124 36318
rect 4956 35810 5012 36316
rect 5068 36306 5124 36316
rect 5068 35924 5124 35934
rect 5068 35830 5124 35868
rect 4956 35758 4958 35810
rect 5010 35758 5012 35810
rect 4956 35746 5012 35758
rect 4956 34916 5012 34926
rect 4956 33346 5012 34860
rect 5180 34692 5236 37772
rect 5852 37492 5908 38670
rect 5852 37426 5908 37436
rect 5964 36820 6020 40348
rect 7196 40404 7252 40414
rect 7196 40310 7252 40348
rect 6860 39842 6916 39854
rect 6860 39790 6862 39842
rect 6914 39790 6916 39842
rect 6860 39730 6916 39790
rect 7532 39842 7588 40462
rect 7532 39790 7534 39842
rect 7586 39790 7588 39842
rect 7532 39778 7588 39790
rect 7868 40514 7924 40526
rect 7868 40462 7870 40514
rect 7922 40462 7924 40514
rect 6860 39678 6862 39730
rect 6914 39678 6916 39730
rect 6860 39666 6916 39678
rect 7196 39732 7252 39742
rect 7196 39638 7252 39676
rect 5740 36764 6020 36820
rect 6412 39396 6468 39406
rect 6412 38836 6468 39340
rect 7644 39396 7700 39406
rect 7644 39302 7700 39340
rect 5628 36484 5684 36494
rect 5292 36482 5684 36484
rect 5292 36430 5630 36482
rect 5682 36430 5684 36482
rect 5292 36428 5684 36430
rect 5292 35922 5348 36428
rect 5628 36418 5684 36428
rect 5292 35870 5294 35922
rect 5346 35870 5348 35922
rect 5292 35858 5348 35870
rect 5740 35812 5796 36764
rect 5852 36596 5908 36606
rect 5852 36502 5908 36540
rect 5964 36484 6020 36494
rect 5964 36390 6020 36428
rect 5516 35756 5796 35812
rect 6300 36370 6356 36382
rect 6300 36318 6302 36370
rect 6354 36318 6356 36370
rect 5516 35140 5572 35756
rect 5628 35586 5684 35598
rect 5628 35534 5630 35586
rect 5682 35534 5684 35586
rect 5628 35252 5684 35534
rect 5964 35476 6020 35486
rect 5628 35196 5908 35252
rect 5516 35084 5684 35140
rect 5516 34916 5572 34926
rect 5516 34822 5572 34860
rect 5180 34636 5460 34692
rect 4956 33294 4958 33346
rect 5010 33294 5012 33346
rect 4956 33282 5012 33294
rect 5292 33572 5348 33582
rect 5068 33012 5124 33022
rect 5124 32956 5236 33012
rect 5068 32946 5124 32956
rect 4060 31166 4062 31218
rect 4114 31166 4116 31218
rect 4060 31154 4116 31166
rect 4284 31612 4900 31668
rect 3724 30994 3780 31006
rect 3724 30942 3726 30994
rect 3778 30942 3780 30994
rect 3724 30212 3780 30942
rect 3724 30146 3780 30156
rect 4060 30100 4116 30110
rect 3836 30098 4116 30100
rect 3836 30046 4062 30098
rect 4114 30046 4116 30098
rect 3836 30044 4116 30046
rect 3836 29650 3892 30044
rect 4060 30034 4116 30044
rect 3836 29598 3838 29650
rect 3890 29598 3892 29650
rect 3836 29586 3892 29598
rect 4172 29652 4228 29662
rect 4172 29558 4228 29596
rect 3836 29428 3892 29438
rect 4284 29428 4340 31612
rect 4620 30882 4676 30894
rect 4620 30830 4622 30882
rect 4674 30830 4676 30882
rect 4620 30772 4676 30830
rect 4620 30716 5012 30772
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4956 30324 5012 30716
rect 4956 30268 5124 30324
rect 4844 30212 4900 30222
rect 4844 30210 5012 30212
rect 4844 30158 4846 30210
rect 4898 30158 5012 30210
rect 4844 30156 5012 30158
rect 4844 30146 4900 30156
rect 4844 29652 4900 29662
rect 4844 29538 4900 29596
rect 4844 29486 4846 29538
rect 4898 29486 4900 29538
rect 4396 29428 4452 29438
rect 4284 29426 4452 29428
rect 4284 29374 4398 29426
rect 4450 29374 4452 29426
rect 4284 29372 4452 29374
rect 3836 29334 3892 29372
rect 4396 29316 4452 29372
rect 4396 29250 4452 29260
rect 3612 29204 3668 29214
rect 3612 29202 4340 29204
rect 3612 29150 3614 29202
rect 3666 29150 4340 29202
rect 3612 29148 4340 29150
rect 3612 29138 3668 29148
rect 4284 28868 4340 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4620 28868 4676 28878
rect 4284 28866 4676 28868
rect 4284 28814 4622 28866
rect 4674 28814 4676 28866
rect 4284 28812 4676 28814
rect 4620 28802 4676 28812
rect 4284 28644 4340 28654
rect 4284 28550 4340 28588
rect 4844 28532 4900 29486
rect 4956 28756 5012 30156
rect 4956 28690 5012 28700
rect 5068 29428 5124 30268
rect 5180 29764 5236 32956
rect 5292 32786 5348 33516
rect 5404 33012 5460 34636
rect 5404 32946 5460 32956
rect 5628 32788 5684 35084
rect 5740 34690 5796 34702
rect 5740 34638 5742 34690
rect 5794 34638 5796 34690
rect 5740 34242 5796 34638
rect 5740 34190 5742 34242
rect 5794 34190 5796 34242
rect 5740 34178 5796 34190
rect 5852 34132 5908 35196
rect 5964 34914 6020 35420
rect 6300 35140 6356 36318
rect 5964 34862 5966 34914
rect 6018 34862 6020 34914
rect 5964 34850 6020 34862
rect 6188 35084 6300 35140
rect 6188 34914 6244 35084
rect 6300 35074 6356 35084
rect 6188 34862 6190 34914
rect 6242 34862 6244 34914
rect 6188 34850 6244 34862
rect 6412 34132 6468 38780
rect 7196 38836 7252 38846
rect 7196 38668 7252 38780
rect 7196 38612 7700 38668
rect 7532 37826 7588 37838
rect 7532 37774 7534 37826
rect 7586 37774 7588 37826
rect 7532 37716 7588 37774
rect 7532 37650 7588 37660
rect 6636 37604 6692 37614
rect 6524 37154 6580 37166
rect 6524 37102 6526 37154
rect 6578 37102 6580 37154
rect 6524 37044 6580 37102
rect 6636 37044 6692 37548
rect 7532 37492 7588 37502
rect 7532 37398 7588 37436
rect 6748 37380 6804 37390
rect 6748 37286 6804 37324
rect 6972 37268 7028 37278
rect 6972 37174 7028 37212
rect 7196 37268 7252 37278
rect 6524 36988 6804 37044
rect 6636 36708 6692 36718
rect 6524 36484 6580 36494
rect 6524 36390 6580 36428
rect 6636 35924 6692 36652
rect 6748 36372 6804 36988
rect 6748 36278 6804 36316
rect 6860 36370 6916 36382
rect 6860 36318 6862 36370
rect 6914 36318 6916 36370
rect 6860 36148 6916 36318
rect 7196 36260 7252 37212
rect 7420 37266 7476 37278
rect 7420 37214 7422 37266
rect 7474 37214 7476 37266
rect 7308 36932 7364 36942
rect 7308 36482 7364 36876
rect 7308 36430 7310 36482
rect 7362 36430 7364 36482
rect 7308 36418 7364 36430
rect 7420 36484 7476 37214
rect 7420 36428 7588 36484
rect 7420 36260 7476 36270
rect 7196 36258 7476 36260
rect 7196 36206 7422 36258
rect 7474 36206 7476 36258
rect 7196 36204 7476 36206
rect 7420 36194 7476 36204
rect 6860 36082 6916 36092
rect 7084 36036 7140 36046
rect 6636 35858 6692 35868
rect 6748 35924 6804 35934
rect 7084 35924 7140 35980
rect 6748 35922 7140 35924
rect 6748 35870 6750 35922
rect 6802 35870 7086 35922
rect 7138 35870 7140 35922
rect 6748 35868 7140 35870
rect 6748 35588 6804 35868
rect 7084 35858 7140 35868
rect 7196 35924 7252 35934
rect 7196 35810 7252 35868
rect 7420 35924 7476 35934
rect 7532 35924 7588 36428
rect 7644 36482 7700 38612
rect 7756 37828 7812 37838
rect 7756 37734 7812 37772
rect 7644 36430 7646 36482
rect 7698 36430 7700 36482
rect 7644 36418 7700 36430
rect 7756 37266 7812 37278
rect 7756 37214 7758 37266
rect 7810 37214 7812 37266
rect 7756 36482 7812 37214
rect 7756 36430 7758 36482
rect 7810 36430 7812 36482
rect 7756 36418 7812 36430
rect 7420 35922 7588 35924
rect 7420 35870 7422 35922
rect 7474 35870 7588 35922
rect 7420 35868 7588 35870
rect 7756 35924 7812 35934
rect 7420 35858 7476 35868
rect 7196 35758 7198 35810
rect 7250 35758 7252 35810
rect 7196 35746 7252 35758
rect 7644 35810 7700 35822
rect 7644 35758 7646 35810
rect 7698 35758 7700 35810
rect 6748 35522 6804 35532
rect 7084 35476 7140 35486
rect 7084 35382 7140 35420
rect 7644 35252 7700 35758
rect 7756 35810 7812 35868
rect 7756 35758 7758 35810
rect 7810 35758 7812 35810
rect 7756 35746 7812 35758
rect 7644 35186 7700 35196
rect 7420 34916 7476 34926
rect 7196 34914 7476 34916
rect 7196 34862 7422 34914
rect 7474 34862 7476 34914
rect 7196 34860 7476 34862
rect 6860 34804 6916 34814
rect 6748 34802 6916 34804
rect 6748 34750 6862 34802
rect 6914 34750 6916 34802
rect 6748 34748 6916 34750
rect 6524 34132 6580 34142
rect 6748 34132 6804 34748
rect 6860 34738 6916 34748
rect 7084 34804 7140 34814
rect 7084 34710 7140 34748
rect 7196 34580 7252 34860
rect 7420 34850 7476 34860
rect 6972 34524 7252 34580
rect 7308 34690 7364 34702
rect 7308 34638 7310 34690
rect 7362 34638 7364 34690
rect 6972 34356 7028 34524
rect 6972 34300 7140 34356
rect 6972 34132 7028 34142
rect 5852 34130 6692 34132
rect 5852 34078 6526 34130
rect 6578 34078 6692 34130
rect 5852 34076 6692 34078
rect 6524 34066 6580 34076
rect 6636 34020 6692 34076
rect 6748 34066 6804 34076
rect 6860 34130 7028 34132
rect 6860 34078 6974 34130
rect 7026 34078 7028 34130
rect 6860 34076 7028 34078
rect 6636 33954 6692 33964
rect 6748 33908 6804 33918
rect 6748 33814 6804 33852
rect 6860 33684 6916 34076
rect 6972 34066 7028 34076
rect 6412 33628 6916 33684
rect 6972 33796 7028 33806
rect 5292 32734 5294 32786
rect 5346 32734 5348 32786
rect 5292 32722 5348 32734
rect 5404 32732 5684 32788
rect 6076 33572 6132 33582
rect 5404 31220 5460 32732
rect 5516 32562 5572 32574
rect 5516 32510 5518 32562
rect 5570 32510 5572 32562
rect 5516 31444 5572 32510
rect 6076 32562 6132 33516
rect 6412 32786 6468 33628
rect 6748 33460 6804 33470
rect 6972 33460 7028 33740
rect 6748 33458 7028 33460
rect 6748 33406 6750 33458
rect 6802 33406 7028 33458
rect 6748 33404 7028 33406
rect 6748 33394 6804 33404
rect 6412 32734 6414 32786
rect 6466 32734 6468 32786
rect 6412 32722 6468 32734
rect 7084 33124 7140 34300
rect 7308 34244 7364 34638
rect 6188 32676 6244 32686
rect 6188 32582 6244 32620
rect 6076 32510 6078 32562
rect 6130 32510 6132 32562
rect 6076 32004 6132 32510
rect 6076 31938 6132 31948
rect 6636 32564 6692 32574
rect 7084 32564 7140 33068
rect 6636 32562 7140 32564
rect 6636 32510 6638 32562
rect 6690 32510 7140 32562
rect 6636 32508 7140 32510
rect 7196 34188 7364 34244
rect 7644 34242 7700 34254
rect 7644 34190 7646 34242
rect 7698 34190 7700 34242
rect 7196 32562 7252 34188
rect 7420 34130 7476 34142
rect 7420 34078 7422 34130
rect 7474 34078 7476 34130
rect 7308 34020 7364 34030
rect 7308 33458 7364 33964
rect 7308 33406 7310 33458
rect 7362 33406 7364 33458
rect 7308 33394 7364 33406
rect 7196 32510 7198 32562
rect 7250 32510 7252 32562
rect 5516 31378 5572 31388
rect 5964 31780 6020 31790
rect 6524 31780 6580 31790
rect 5964 31778 6580 31780
rect 5964 31726 5966 31778
rect 6018 31726 6526 31778
rect 6578 31726 6580 31778
rect 5964 31724 6580 31726
rect 5964 31332 6020 31724
rect 6524 31714 6580 31724
rect 6188 31556 6244 31566
rect 6636 31556 6692 32508
rect 7196 32498 7252 32510
rect 7308 33012 7364 33022
rect 6972 32338 7028 32350
rect 6972 32286 6974 32338
rect 7026 32286 7028 32338
rect 6748 32004 6804 32014
rect 6804 31948 6916 32004
rect 6748 31938 6804 31948
rect 6188 31554 6692 31556
rect 6188 31502 6190 31554
rect 6242 31502 6692 31554
rect 6188 31500 6692 31502
rect 6188 31490 6244 31500
rect 5964 31276 6244 31332
rect 5404 31218 6132 31220
rect 5404 31166 5406 31218
rect 5458 31166 6132 31218
rect 5404 31164 6132 31166
rect 5404 31154 5460 31164
rect 5740 30212 5796 30222
rect 5740 29986 5796 30156
rect 5740 29934 5742 29986
rect 5794 29934 5796 29986
rect 5740 29922 5796 29934
rect 5180 29708 5460 29764
rect 5292 29540 5348 29550
rect 4956 28532 5012 28542
rect 4844 28530 5012 28532
rect 4844 28478 4958 28530
rect 5010 28478 5012 28530
rect 4844 28476 5012 28478
rect 4956 28466 5012 28476
rect 4732 28418 4788 28430
rect 4732 28366 4734 28418
rect 4786 28366 4788 28418
rect 4284 27860 4340 27870
rect 4284 27766 4340 27804
rect 4732 27746 4788 28366
rect 4732 27694 4734 27746
rect 4786 27694 4788 27746
rect 4732 27636 4788 27694
rect 4284 27580 4788 27636
rect 3724 27076 3780 27086
rect 3724 26178 3780 27020
rect 4172 27076 4228 27114
rect 4172 27010 4228 27020
rect 4284 26908 4340 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 3724 26126 3726 26178
rect 3778 26126 3780 26178
rect 3724 26114 3780 26126
rect 4060 26852 4340 26908
rect 3836 25394 3892 25406
rect 3836 25342 3838 25394
rect 3890 25342 3892 25394
rect 3836 25284 3892 25342
rect 3836 25218 3892 25228
rect 3836 24052 3892 24062
rect 3836 23958 3892 23996
rect 3500 23492 4004 23548
rect 3948 23380 4004 23492
rect 3724 23324 4004 23380
rect 3612 23044 3668 23054
rect 3612 22950 3668 22988
rect 3500 21700 3556 21710
rect 3388 21644 3500 21700
rect 3164 18340 3220 18350
rect 3164 18246 3220 18284
rect 3164 17780 3220 17790
rect 3052 17778 3220 17780
rect 3052 17726 3166 17778
rect 3218 17726 3220 17778
rect 3052 17724 3220 17726
rect 3164 17714 3220 17724
rect 3276 17780 3332 17790
rect 3276 17686 3332 17724
rect 2940 17108 2996 17118
rect 3388 17108 3444 21644
rect 3500 21634 3556 21644
rect 3724 19908 3780 23324
rect 3948 21364 4004 21374
rect 3836 20916 3892 20926
rect 3836 20822 3892 20860
rect 3836 19908 3892 19918
rect 3724 19852 3836 19908
rect 3836 19842 3892 19852
rect 3948 19234 4004 21308
rect 3948 19182 3950 19234
rect 4002 19182 4004 19234
rect 3948 19170 4004 19182
rect 4060 19012 4116 26852
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4620 25508 4676 25518
rect 4844 25508 4900 25518
rect 4620 25506 4844 25508
rect 4620 25454 4622 25506
rect 4674 25454 4844 25506
rect 4620 25452 4844 25454
rect 4620 25442 4676 25452
rect 4284 25396 4340 25406
rect 4284 24722 4340 25340
rect 4284 24670 4286 24722
rect 4338 24670 4340 24722
rect 4284 24658 4340 24670
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4620 23940 4676 23950
rect 4844 23940 4900 25452
rect 5068 24500 5124 29372
rect 5180 29538 5348 29540
rect 5180 29486 5294 29538
rect 5346 29486 5348 29538
rect 5180 29484 5348 29486
rect 5180 29426 5236 29484
rect 5292 29474 5348 29484
rect 5180 29374 5182 29426
rect 5234 29374 5236 29426
rect 5180 29362 5236 29374
rect 5404 29316 5460 29708
rect 5516 29538 5572 29550
rect 5516 29486 5518 29538
rect 5570 29486 5572 29538
rect 5516 29428 5572 29486
rect 5516 29372 5684 29428
rect 5292 29260 5460 29316
rect 5628 29314 5684 29372
rect 5628 29262 5630 29314
rect 5682 29262 5684 29314
rect 5180 29204 5236 29214
rect 5292 29204 5348 29260
rect 5180 29202 5348 29204
rect 5180 29150 5182 29202
rect 5234 29150 5348 29202
rect 5180 29148 5348 29150
rect 5180 29138 5236 29148
rect 5628 24836 5684 29262
rect 5852 26908 5908 31164
rect 6076 30434 6132 31164
rect 6076 30382 6078 30434
rect 6130 30382 6132 30434
rect 6076 30370 6132 30382
rect 6188 30212 6244 31276
rect 6076 30156 6244 30212
rect 6076 29540 6132 30156
rect 6300 30098 6356 30110
rect 6300 30046 6302 30098
rect 6354 30046 6356 30098
rect 6300 29988 6356 30046
rect 6748 29988 6804 29998
rect 6300 29986 6804 29988
rect 6300 29934 6750 29986
rect 6802 29934 6804 29986
rect 6300 29932 6804 29934
rect 6748 29764 6804 29932
rect 6748 29698 6804 29708
rect 5964 29538 6132 29540
rect 5964 29486 6078 29538
rect 6130 29486 6132 29538
rect 5964 29484 6132 29486
rect 5964 28980 6020 29484
rect 6076 29474 6132 29484
rect 6188 29426 6244 29438
rect 6188 29374 6190 29426
rect 6242 29374 6244 29426
rect 6076 29316 6132 29326
rect 6188 29316 6244 29374
rect 6636 29316 6692 29326
rect 6188 29314 6692 29316
rect 6188 29262 6638 29314
rect 6690 29262 6692 29314
rect 6188 29260 6692 29262
rect 6076 29202 6132 29260
rect 6076 29150 6078 29202
rect 6130 29150 6132 29202
rect 6076 29138 6132 29150
rect 6636 29204 6692 29260
rect 6636 29138 6692 29148
rect 5964 28924 6244 28980
rect 5852 26852 6132 26908
rect 5852 26516 5908 26526
rect 5852 26402 5908 26460
rect 5852 26350 5854 26402
rect 5906 26350 5908 26402
rect 5852 26338 5908 26350
rect 5852 25620 5908 25630
rect 5852 25526 5908 25564
rect 5740 25396 5796 25406
rect 5740 25302 5796 25340
rect 5628 24780 5908 24836
rect 5068 24434 5124 24444
rect 5740 24612 5796 24622
rect 5740 24162 5796 24556
rect 5740 24110 5742 24162
rect 5794 24110 5796 24162
rect 5740 24098 5796 24110
rect 4620 23938 4900 23940
rect 4620 23886 4622 23938
rect 4674 23886 4900 23938
rect 4620 23884 4900 23886
rect 4620 23874 4676 23884
rect 4284 23828 4340 23838
rect 4172 23044 4228 23054
rect 4172 21586 4228 22988
rect 4284 22370 4340 23772
rect 5628 23828 5684 23838
rect 5628 23734 5684 23772
rect 5740 23716 5796 23726
rect 5740 23266 5796 23660
rect 5740 23214 5742 23266
rect 5794 23214 5796 23266
rect 5740 23202 5796 23214
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 22318 4286 22370
rect 4338 22318 4340 22370
rect 4284 22306 4340 22318
rect 4172 21534 4174 21586
rect 4226 21534 4228 21586
rect 4172 21522 4228 21534
rect 5068 21474 5124 21486
rect 5068 21422 5070 21474
rect 5122 21422 5124 21474
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4284 20804 4340 20814
rect 4284 20018 4340 20748
rect 4620 20802 4676 20814
rect 4620 20750 4622 20802
rect 4674 20750 4676 20802
rect 4620 20580 4676 20750
rect 5068 20804 5124 21422
rect 5180 21476 5236 21486
rect 5180 21382 5236 21420
rect 5068 20738 5124 20748
rect 5068 20580 5124 20590
rect 4620 20578 5124 20580
rect 4620 20526 5070 20578
rect 5122 20526 5124 20578
rect 4620 20524 5124 20526
rect 4284 19966 4286 20018
rect 4338 19966 4340 20018
rect 4284 19954 4340 19966
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 3724 18956 4116 19012
rect 4732 19010 4788 19022
rect 4732 18958 4734 19010
rect 4786 18958 4788 19010
rect 3612 18452 3668 18462
rect 3500 18450 3668 18452
rect 3500 18398 3614 18450
rect 3666 18398 3668 18450
rect 3500 18396 3668 18398
rect 3500 17892 3556 18396
rect 3612 18386 3668 18396
rect 3724 18228 3780 18956
rect 4508 18450 4564 18462
rect 4508 18398 4510 18450
rect 4562 18398 4564 18450
rect 3500 17826 3556 17836
rect 3612 18172 3780 18228
rect 3836 18340 3892 18350
rect 3500 17108 3556 17118
rect 3388 17106 3556 17108
rect 3388 17054 3502 17106
rect 3554 17054 3556 17106
rect 3388 17052 3556 17054
rect 2604 16882 2660 16894
rect 2940 16884 2996 17052
rect 3500 17042 3556 17052
rect 3276 16996 3332 17006
rect 3332 16940 3444 16996
rect 3276 16930 3332 16940
rect 2604 16830 2606 16882
rect 2658 16830 2660 16882
rect 2604 16212 2660 16830
rect 2604 16146 2660 16156
rect 2716 16882 2996 16884
rect 2716 16830 2942 16882
rect 2994 16830 2996 16882
rect 2716 16828 2996 16830
rect 2604 15874 2660 15886
rect 2604 15822 2606 15874
rect 2658 15822 2660 15874
rect 2604 14980 2660 15822
rect 2604 14914 2660 14924
rect 2380 14812 2548 14868
rect 2268 14756 2324 14766
rect 1932 14254 1934 14306
rect 1986 14254 1988 14306
rect 1820 13748 1876 13758
rect 1820 12962 1876 13692
rect 1820 12910 1822 12962
rect 1874 12910 1876 12962
rect 1596 11554 1652 11564
rect 1708 12178 1764 12190
rect 1708 12126 1710 12178
rect 1762 12126 1764 12178
rect 1708 11732 1764 12126
rect 1708 11060 1764 11676
rect 1820 11506 1876 12910
rect 1820 11454 1822 11506
rect 1874 11454 1876 11506
rect 1820 11442 1876 11454
rect 1708 10994 1764 11004
rect 1820 10498 1876 10510
rect 1820 10446 1822 10498
rect 1874 10446 1876 10498
rect 1708 9716 1764 9726
rect 1820 9716 1876 10446
rect 1764 9660 1876 9716
rect 1708 9622 1764 9660
rect 1708 9042 1764 9054
rect 1708 8990 1710 9042
rect 1762 8990 1764 9042
rect 1708 8372 1764 8990
rect 1932 8428 1988 14254
rect 2156 14308 2212 14318
rect 2156 13074 2212 14252
rect 2268 13746 2324 14700
rect 2380 14420 2436 14812
rect 2492 14644 2548 14654
rect 2716 14644 2772 16828
rect 2940 16818 2996 16828
rect 3164 16658 3220 16670
rect 3164 16606 3166 16658
rect 3218 16606 3220 16658
rect 3164 16324 3220 16606
rect 2940 16268 3220 16324
rect 3388 16324 3444 16940
rect 3388 16268 3556 16324
rect 2940 15988 2996 16268
rect 3052 16100 3108 16110
rect 3276 16100 3332 16110
rect 3108 16044 3220 16100
rect 3052 16006 3108 16044
rect 2940 15894 2996 15932
rect 2492 14642 2772 14644
rect 2492 14590 2494 14642
rect 2546 14590 2772 14642
rect 2492 14588 2772 14590
rect 2828 15314 2884 15326
rect 2828 15262 2830 15314
rect 2882 15262 2884 15314
rect 2492 14578 2548 14588
rect 2828 14532 2884 15262
rect 3164 15316 3220 16044
rect 3276 16006 3332 16044
rect 3388 16098 3444 16110
rect 3388 16046 3390 16098
rect 3442 16046 3444 16098
rect 3388 15876 3444 16046
rect 3388 15810 3444 15820
rect 3388 15540 3444 15550
rect 3500 15540 3556 16268
rect 3388 15538 3556 15540
rect 3388 15486 3390 15538
rect 3442 15486 3556 15538
rect 3388 15484 3556 15486
rect 3388 15474 3444 15484
rect 3500 15316 3556 15326
rect 3164 15260 3444 15316
rect 3052 15092 3108 15102
rect 3052 14998 3108 15036
rect 3164 14532 3220 14542
rect 2828 14530 3332 14532
rect 2828 14478 3166 14530
rect 3218 14478 3332 14530
rect 2828 14476 3332 14478
rect 3164 14466 3220 14476
rect 2380 14364 3108 14420
rect 3052 14308 3108 14364
rect 3052 14252 3220 14308
rect 2268 13694 2270 13746
rect 2322 13694 2324 13746
rect 2268 13682 2324 13694
rect 2492 14196 2548 14206
rect 2156 13022 2158 13074
rect 2210 13022 2212 13074
rect 2156 13010 2212 13022
rect 2492 12964 2548 14140
rect 2716 13972 2772 13982
rect 2716 13878 2772 13916
rect 3164 13860 3220 14252
rect 3052 13746 3108 13758
rect 3052 13694 3054 13746
rect 3106 13694 3108 13746
rect 2380 12908 2548 12964
rect 2716 12962 2772 12974
rect 2716 12910 2718 12962
rect 2770 12910 2772 12962
rect 2268 12180 2324 12190
rect 2268 12086 2324 12124
rect 2268 11394 2324 11406
rect 2268 11342 2270 11394
rect 2322 11342 2324 11394
rect 2268 10612 2324 11342
rect 2268 10518 2324 10556
rect 2268 9940 2324 9950
rect 2268 9846 2324 9884
rect 2044 9380 2100 9390
rect 2044 9266 2100 9324
rect 2044 9214 2046 9266
rect 2098 9214 2100 9266
rect 2044 9202 2100 9214
rect 1932 8372 2100 8428
rect 1708 8306 1764 8316
rect 2044 7698 2100 8372
rect 2044 7646 2046 7698
rect 2098 7646 2100 7698
rect 2044 7634 2100 7646
rect 1708 7474 1764 7486
rect 1708 7422 1710 7474
rect 1762 7422 1764 7474
rect 1708 7028 1764 7422
rect 1708 6962 1764 6972
rect 2380 6356 2436 12908
rect 2604 12852 2660 12862
rect 2492 8930 2548 8942
rect 2492 8878 2494 8930
rect 2546 8878 2548 8930
rect 2492 8372 2548 8878
rect 2492 8306 2548 8316
rect 2492 7362 2548 7374
rect 2492 7310 2494 7362
rect 2546 7310 2548 7362
rect 2492 7028 2548 7310
rect 2492 6962 2548 6972
rect 1932 6300 2436 6356
rect 1708 5906 1764 5918
rect 1708 5854 1710 5906
rect 1762 5854 1764 5906
rect 1708 5684 1764 5854
rect 1708 5618 1764 5628
rect 1708 5122 1764 5134
rect 1708 5070 1710 5122
rect 1762 5070 1764 5122
rect 1708 4900 1764 5070
rect 1708 4340 1764 4844
rect 1708 4274 1764 4284
rect 1820 4338 1876 4350
rect 1820 4286 1822 4338
rect 1874 4286 1876 4338
rect 1820 3442 1876 4286
rect 1932 4228 1988 6300
rect 2156 6132 2212 6142
rect 2044 6076 2156 6132
rect 2044 6018 2100 6076
rect 2156 6066 2212 6076
rect 2044 5966 2046 6018
rect 2098 5966 2100 6018
rect 2044 5954 2100 5966
rect 2492 5794 2548 5806
rect 2492 5742 2494 5794
rect 2546 5742 2548 5794
rect 2492 5684 2548 5742
rect 2492 5618 2548 5628
rect 2604 5460 2660 12796
rect 2716 12404 2772 12910
rect 3052 12852 3108 13694
rect 3164 13074 3220 13804
rect 3164 13022 3166 13074
rect 3218 13022 3220 13074
rect 3164 13010 3220 13022
rect 3276 13636 3332 14476
rect 3388 14196 3444 15260
rect 3500 14642 3556 15260
rect 3500 14590 3502 14642
rect 3554 14590 3556 14642
rect 3500 14578 3556 14590
rect 3612 14420 3668 18172
rect 3836 16884 3892 18284
rect 4172 18338 4228 18350
rect 4172 18286 4174 18338
rect 4226 18286 4228 18338
rect 3836 16790 3892 16828
rect 3948 17892 4004 17902
rect 3948 16324 4004 17836
rect 4172 17892 4228 18286
rect 4508 18340 4564 18398
rect 4732 18452 4788 18958
rect 4732 18386 4788 18396
rect 4508 18274 4564 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4844 18004 4900 20524
rect 5068 20514 5124 20524
rect 5852 19796 5908 24780
rect 6076 22484 6132 26852
rect 6076 22418 6132 22428
rect 6076 21474 6132 21486
rect 6076 21422 6078 21474
rect 6130 21422 6132 21474
rect 6076 21364 6132 21422
rect 6188 21364 6244 28924
rect 6300 28754 6356 28766
rect 6300 28702 6302 28754
rect 6354 28702 6356 28754
rect 6300 28644 6356 28702
rect 6300 28578 6356 28588
rect 6636 28756 6692 28766
rect 6524 26292 6580 26302
rect 6636 26292 6692 28700
rect 6860 27524 6916 31948
rect 6972 29652 7028 32286
rect 7084 31892 7140 31902
rect 7084 31798 7140 31836
rect 7308 31778 7364 32956
rect 7420 32788 7476 34078
rect 7420 32722 7476 32732
rect 7532 33908 7588 33918
rect 7308 31726 7310 31778
rect 7362 31726 7364 31778
rect 7308 31714 7364 31726
rect 6972 29586 7028 29596
rect 7420 30996 7476 31006
rect 6860 27458 6916 27468
rect 7084 27188 7140 27198
rect 6748 27076 6804 27086
rect 6748 26982 6804 27020
rect 6860 26852 6916 26862
rect 6860 26758 6916 26796
rect 6972 26516 7028 26526
rect 6972 26422 7028 26460
rect 7084 26404 7140 27132
rect 7084 26310 7140 26348
rect 7308 26852 7364 26862
rect 6524 26290 6692 26292
rect 6524 26238 6526 26290
rect 6578 26238 6692 26290
rect 6524 26236 6692 26238
rect 7308 26290 7364 26796
rect 7308 26238 7310 26290
rect 7362 26238 7364 26290
rect 6524 25508 6580 26236
rect 7308 26226 7364 26238
rect 7084 25956 7140 25966
rect 7084 25508 7140 25900
rect 7308 25620 7364 25630
rect 7308 25526 7364 25564
rect 6524 25442 6580 25452
rect 6748 25506 7140 25508
rect 6748 25454 7086 25506
rect 7138 25454 7140 25506
rect 6748 25452 7140 25454
rect 6748 24834 6804 25452
rect 7084 25442 7140 25452
rect 6972 25284 7028 25294
rect 6972 25190 7028 25228
rect 7420 25060 7476 30940
rect 7532 30436 7588 33852
rect 7644 33684 7700 34190
rect 7644 33618 7700 33628
rect 7756 34018 7812 34030
rect 7756 33966 7758 34018
rect 7810 33966 7812 34018
rect 7756 33908 7812 33966
rect 7756 33460 7812 33852
rect 7868 33684 7924 40462
rect 7980 39394 8036 39406
rect 7980 39342 7982 39394
rect 8034 39342 8036 39394
rect 7980 38948 8036 39342
rect 7980 38882 8036 38892
rect 7980 38724 8036 38734
rect 8092 38724 8148 40684
rect 8204 40674 8260 40684
rect 8316 40628 8372 44200
rect 8540 41746 8596 41758
rect 8540 41694 8542 41746
rect 8594 41694 8596 41746
rect 8540 41186 8596 41694
rect 9436 41746 9492 44200
rect 9436 41694 9438 41746
rect 9490 41694 9492 41746
rect 9436 41298 9492 41694
rect 9436 41246 9438 41298
rect 9490 41246 9492 41298
rect 9436 41234 9492 41246
rect 8540 41134 8542 41186
rect 8594 41134 8596 41186
rect 8540 41122 8596 41134
rect 8764 40964 8820 40974
rect 8764 40962 9380 40964
rect 8764 40910 8766 40962
rect 8818 40910 9380 40962
rect 8764 40908 9380 40910
rect 8764 40898 8820 40908
rect 8316 40516 8372 40572
rect 8428 40516 8484 40526
rect 8764 40516 8820 40526
rect 8316 40514 8484 40516
rect 8316 40462 8430 40514
rect 8482 40462 8484 40514
rect 8316 40460 8484 40462
rect 8428 40450 8484 40460
rect 8540 40514 8820 40516
rect 8540 40462 8766 40514
rect 8818 40462 8820 40514
rect 8540 40460 8820 40462
rect 8204 39732 8260 39742
rect 8204 39060 8260 39676
rect 8316 39506 8372 39518
rect 8316 39454 8318 39506
rect 8370 39454 8372 39506
rect 8316 39284 8372 39454
rect 8316 39228 8484 39284
rect 8316 39060 8372 39070
rect 8204 39058 8372 39060
rect 8204 39006 8318 39058
rect 8370 39006 8372 39058
rect 8204 39004 8372 39006
rect 8316 38994 8372 39004
rect 7980 38722 8148 38724
rect 7980 38670 7982 38722
rect 8034 38670 8148 38722
rect 7980 38668 8148 38670
rect 7980 37940 8036 38668
rect 7980 37874 8036 37884
rect 8092 38500 8148 38510
rect 8092 37938 8148 38444
rect 8092 37886 8094 37938
rect 8146 37886 8148 37938
rect 7980 37716 8036 37726
rect 7980 37266 8036 37660
rect 7980 37214 7982 37266
rect 8034 37214 8036 37266
rect 7980 36820 8036 37214
rect 7980 36754 8036 36764
rect 8092 36708 8148 37886
rect 8428 38162 8484 39228
rect 8428 38110 8430 38162
rect 8482 38110 8484 38162
rect 8428 37378 8484 38110
rect 8428 37326 8430 37378
rect 8482 37326 8484 37378
rect 8316 37266 8372 37278
rect 8316 37214 8318 37266
rect 8370 37214 8372 37266
rect 8316 36932 8372 37214
rect 8428 37044 8484 37326
rect 8428 36978 8484 36988
rect 8316 36866 8372 36876
rect 8540 36932 8596 40460
rect 8764 40450 8820 40460
rect 8652 39618 8708 39630
rect 8652 39566 8654 39618
rect 8706 39566 8708 39618
rect 8652 39396 8708 39566
rect 8652 39330 8708 39340
rect 8764 38724 8820 38734
rect 8764 38630 8820 38668
rect 9324 38668 9380 40908
rect 9660 40628 9716 40638
rect 9660 40534 9716 40572
rect 10556 40404 10612 44200
rect 11676 42196 11732 44200
rect 11228 42140 11732 42196
rect 11228 41300 11284 42140
rect 11228 41206 11284 41244
rect 12124 41300 12180 41310
rect 11676 41188 11732 41198
rect 11564 41186 11732 41188
rect 11564 41134 11678 41186
rect 11730 41134 11732 41186
rect 11564 41132 11732 41134
rect 11452 41076 11508 41086
rect 11452 40982 11508 41020
rect 10556 40338 10612 40348
rect 11452 40404 11508 40414
rect 11452 40310 11508 40348
rect 11564 39730 11620 41132
rect 11676 41122 11732 41132
rect 12124 41186 12180 41244
rect 12124 41134 12126 41186
rect 12178 41134 12180 41186
rect 12124 41122 12180 41134
rect 12796 41188 12852 44200
rect 13916 41972 13972 44200
rect 13916 41916 14420 41972
rect 13132 41188 13188 41198
rect 12796 41186 13188 41188
rect 12796 41134 13134 41186
rect 13186 41134 13188 41186
rect 12796 41132 13188 41134
rect 12460 40964 12516 40974
rect 12460 40962 13076 40964
rect 12460 40910 12462 40962
rect 12514 40910 13076 40962
rect 12460 40908 13076 40910
rect 12460 40898 12516 40908
rect 11900 40740 11956 40750
rect 11676 40516 11732 40526
rect 11676 40422 11732 40460
rect 11900 40402 11956 40684
rect 12684 40514 12740 40526
rect 12684 40462 12686 40514
rect 12738 40462 12740 40514
rect 11900 40350 11902 40402
rect 11954 40350 11956 40402
rect 11900 40338 11956 40350
rect 12348 40404 12404 40414
rect 12348 40310 12404 40348
rect 11564 39678 11566 39730
rect 11618 39678 11620 39730
rect 9436 39508 9492 39518
rect 9436 39506 9716 39508
rect 9436 39454 9438 39506
rect 9490 39454 9716 39506
rect 9436 39452 9716 39454
rect 9436 39442 9492 39452
rect 9660 39058 9716 39452
rect 9660 39006 9662 39058
rect 9714 39006 9716 39058
rect 9660 38994 9716 39006
rect 9436 38836 9492 38846
rect 9436 38742 9492 38780
rect 9884 38834 9940 38846
rect 9884 38782 9886 38834
rect 9938 38782 9940 38834
rect 9324 38612 9604 38668
rect 8652 37380 8708 37390
rect 8652 37378 9156 37380
rect 8652 37326 8654 37378
rect 8706 37326 9156 37378
rect 8652 37324 9156 37326
rect 8652 37314 8708 37324
rect 9100 37268 9156 37324
rect 9436 37268 9492 37278
rect 9100 37266 9492 37268
rect 9100 37214 9438 37266
rect 9490 37214 9492 37266
rect 9100 37212 9492 37214
rect 9436 37202 9492 37212
rect 8540 36866 8596 36876
rect 8988 37154 9044 37166
rect 8988 37102 8990 37154
rect 9042 37102 9044 37154
rect 8092 36642 8148 36652
rect 8428 36820 8484 36830
rect 8092 36484 8148 36494
rect 8092 36390 8148 36428
rect 8428 36484 8484 36764
rect 8988 36820 9044 37102
rect 8428 36390 8484 36428
rect 8764 36484 8820 36494
rect 8204 36372 8260 36382
rect 7980 36258 8036 36270
rect 7980 36206 7982 36258
rect 8034 36206 8036 36258
rect 7980 35588 8036 36206
rect 7980 35522 8036 35532
rect 8204 35252 8260 36316
rect 8764 36370 8820 36428
rect 8764 36318 8766 36370
rect 8818 36318 8820 36370
rect 8764 36148 8820 36318
rect 8764 36082 8820 36092
rect 8988 35698 9044 36764
rect 8988 35646 8990 35698
rect 9042 35646 9044 35698
rect 8204 35186 8260 35196
rect 8540 35588 8596 35598
rect 8316 34018 8372 34030
rect 8316 33966 8318 34018
rect 8370 33966 8372 34018
rect 8092 33908 8148 33918
rect 8316 33908 8372 33966
rect 8148 33852 8372 33908
rect 8092 33842 8148 33852
rect 8540 33684 8596 35532
rect 7868 33628 8372 33684
rect 7756 33404 7924 33460
rect 7756 33236 7812 33246
rect 7756 33142 7812 33180
rect 7644 32564 7700 32602
rect 7644 32498 7700 32508
rect 7756 32562 7812 32574
rect 7756 32510 7758 32562
rect 7810 32510 7812 32562
rect 7756 32452 7812 32510
rect 7868 32452 7924 33404
rect 8092 33234 8148 33246
rect 8092 33182 8094 33234
rect 8146 33182 8148 33234
rect 8092 33012 8148 33182
rect 8092 32946 8148 32956
rect 8316 32674 8372 33628
rect 8316 32622 8318 32674
rect 8370 32622 8372 32674
rect 8316 32610 8372 32622
rect 8428 33628 8596 33684
rect 7980 32452 8036 32462
rect 7868 32450 8036 32452
rect 7868 32398 7982 32450
rect 8034 32398 8036 32450
rect 7868 32396 8036 32398
rect 7756 32386 7812 32396
rect 7868 31778 7924 31790
rect 7868 31726 7870 31778
rect 7922 31726 7924 31778
rect 7644 31666 7700 31678
rect 7644 31614 7646 31666
rect 7698 31614 7700 31666
rect 7644 31556 7700 31614
rect 7644 31490 7700 31500
rect 7868 30436 7924 31726
rect 7532 30380 7700 30436
rect 7532 27188 7588 27198
rect 7532 26962 7588 27132
rect 7532 26910 7534 26962
rect 7586 26910 7588 26962
rect 7532 26898 7588 26910
rect 6748 24782 6750 24834
rect 6802 24782 6804 24834
rect 6748 24770 6804 24782
rect 7084 25004 7476 25060
rect 7532 26066 7588 26078
rect 7532 26014 7534 26066
rect 7586 26014 7588 26066
rect 7532 25506 7588 26014
rect 7532 25454 7534 25506
rect 7586 25454 7588 25506
rect 6860 24610 6916 24622
rect 6860 24558 6862 24610
rect 6914 24558 6916 24610
rect 6860 24052 6916 24558
rect 6972 24612 7028 24622
rect 6972 24518 7028 24556
rect 6860 23986 6916 23996
rect 6524 23154 6580 23166
rect 6524 23102 6526 23154
rect 6578 23102 6580 23154
rect 6524 21588 6580 23102
rect 6524 21522 6580 21532
rect 6188 21308 6804 21364
rect 6076 21298 6132 21308
rect 5964 20020 6020 20030
rect 5964 20018 6132 20020
rect 5964 19966 5966 20018
rect 6018 19966 6132 20018
rect 5964 19964 6132 19966
rect 5964 19954 6020 19964
rect 5852 19740 6020 19796
rect 5740 19234 5796 19246
rect 5740 19182 5742 19234
rect 5794 19182 5796 19234
rect 5740 19124 5796 19182
rect 5740 19058 5796 19068
rect 5852 19122 5908 19134
rect 5852 19070 5854 19122
rect 5906 19070 5908 19122
rect 5516 18452 5572 18462
rect 5404 18226 5460 18238
rect 5404 18174 5406 18226
rect 5458 18174 5460 18226
rect 5404 18116 5460 18174
rect 5404 18050 5460 18060
rect 5068 18004 5124 18014
rect 4844 17948 5012 18004
rect 4172 17826 4228 17836
rect 4284 17668 4340 17678
rect 4172 17556 4228 17566
rect 4060 17108 4116 17118
rect 4172 17108 4228 17500
rect 4060 17106 4228 17108
rect 4060 17054 4062 17106
rect 4114 17054 4228 17106
rect 4060 17052 4228 17054
rect 4284 17106 4340 17612
rect 4508 17554 4564 17566
rect 4508 17502 4510 17554
rect 4562 17502 4564 17554
rect 4508 17220 4564 17502
rect 4284 17054 4286 17106
rect 4338 17054 4340 17106
rect 4060 17042 4116 17052
rect 4284 16884 4340 17054
rect 4396 17164 4508 17220
rect 4396 16996 4452 17164
rect 4508 17154 4564 17164
rect 4396 16930 4452 16940
rect 4284 16818 4340 16828
rect 4508 16882 4564 16894
rect 4508 16830 4510 16882
rect 4562 16830 4564 16882
rect 4508 16660 4564 16830
rect 4844 16882 4900 16894
rect 4844 16830 4846 16882
rect 4898 16830 4900 16882
rect 4620 16772 4676 16782
rect 4620 16678 4676 16716
rect 3948 16100 4004 16268
rect 4284 16604 4564 16660
rect 3948 15316 4004 16044
rect 3388 14130 3444 14140
rect 3500 14364 3668 14420
rect 3724 15314 4004 15316
rect 3724 15262 3950 15314
rect 4002 15262 4004 15314
rect 3724 15260 4004 15262
rect 3052 12786 3108 12796
rect 2716 12310 2772 12348
rect 3164 12066 3220 12078
rect 3164 12014 3166 12066
rect 3218 12014 3220 12066
rect 3164 11732 3220 12014
rect 3164 11666 3220 11676
rect 2940 11284 2996 11294
rect 2940 11190 2996 11228
rect 3052 11172 3108 11182
rect 2940 10724 2996 10734
rect 3052 10724 3108 11116
rect 2940 10722 3108 10724
rect 2940 10670 2942 10722
rect 2994 10670 3108 10722
rect 2940 10668 3108 10670
rect 2940 10658 2996 10668
rect 3276 6132 3332 13580
rect 3500 13188 3556 14364
rect 3612 13860 3668 13870
rect 3724 13860 3780 15260
rect 3948 15250 4004 15260
rect 4172 16212 4228 16222
rect 4172 15316 4228 16156
rect 3612 13858 3780 13860
rect 3612 13806 3614 13858
rect 3666 13806 3780 13858
rect 3612 13804 3780 13806
rect 3836 15092 3892 15102
rect 3612 13794 3668 13804
rect 3500 13122 3556 13132
rect 3836 13074 3892 15036
rect 3948 13636 4004 13646
rect 3948 13542 4004 13580
rect 4172 13634 4228 15260
rect 4284 14644 4340 16604
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4844 16324 4900 16830
rect 4844 16258 4900 16268
rect 4508 16212 4564 16222
rect 4508 16118 4564 16156
rect 4732 16100 4788 16110
rect 4732 16006 4788 16044
rect 4620 15426 4676 15438
rect 4620 15374 4622 15426
rect 4674 15374 4676 15426
rect 4620 15092 4676 15374
rect 4620 15036 4900 15092
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4284 14578 4340 14588
rect 4508 14308 4564 14318
rect 4844 14308 4900 15036
rect 4508 14306 4900 14308
rect 4508 14254 4510 14306
rect 4562 14254 4900 14306
rect 4508 14252 4900 14254
rect 4508 14196 4564 14252
rect 4508 14130 4564 14140
rect 4172 13582 4174 13634
rect 4226 13582 4228 13634
rect 4172 13570 4228 13582
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 3836 13022 3838 13074
rect 3890 13022 3892 13074
rect 3836 13010 3892 13022
rect 4284 13188 4340 13198
rect 3500 12852 3556 12862
rect 3500 12758 3556 12796
rect 4172 11956 4228 11966
rect 4172 8428 4228 11900
rect 4284 9940 4340 13132
rect 4956 12516 5012 17948
rect 5068 17668 5124 17948
rect 5516 17892 5572 18396
rect 5516 17826 5572 17836
rect 5740 18452 5796 18462
rect 5852 18452 5908 19070
rect 5740 18450 5908 18452
rect 5740 18398 5742 18450
rect 5794 18398 5908 18450
rect 5740 18396 5908 18398
rect 5068 17574 5124 17612
rect 5292 17668 5348 17678
rect 5292 17108 5348 17612
rect 5292 17042 5348 17052
rect 5740 16884 5796 18396
rect 5852 17668 5908 17678
rect 5852 17574 5908 17612
rect 5628 16098 5684 16110
rect 5628 16046 5630 16098
rect 5682 16046 5684 16098
rect 5068 15988 5124 15998
rect 5068 15894 5124 15932
rect 5628 15316 5684 16046
rect 5740 15876 5796 16828
rect 5852 17442 5908 17454
rect 5852 17390 5854 17442
rect 5906 17390 5908 17442
rect 5852 16996 5908 17390
rect 5852 16212 5908 16940
rect 5852 16146 5908 16156
rect 5740 15810 5796 15820
rect 5740 15316 5796 15326
rect 5628 15260 5740 15316
rect 5740 15250 5796 15260
rect 5628 15092 5684 15102
rect 5068 14644 5124 14654
rect 5068 14550 5124 14588
rect 5628 14530 5684 15036
rect 5964 14756 6020 19740
rect 6076 17780 6132 19964
rect 6412 19906 6468 19918
rect 6412 19854 6414 19906
rect 6466 19854 6468 19906
rect 6412 19124 6468 19854
rect 6412 19058 6468 19068
rect 6636 19234 6692 19246
rect 6636 19182 6638 19234
rect 6690 19182 6692 19234
rect 6300 18562 6356 18574
rect 6300 18510 6302 18562
rect 6354 18510 6356 18562
rect 6300 18340 6356 18510
rect 6636 18452 6692 19182
rect 6636 18386 6692 18396
rect 6356 18284 6468 18340
rect 6300 18274 6356 18284
rect 6076 16994 6132 17724
rect 6412 17554 6468 18284
rect 6412 17502 6414 17554
rect 6466 17502 6468 17554
rect 6412 17490 6468 17502
rect 6636 17668 6692 17678
rect 6076 16942 6078 16994
rect 6130 16942 6132 16994
rect 6076 16930 6132 16942
rect 6524 17108 6580 17118
rect 6300 16436 6356 16446
rect 6300 15538 6356 16380
rect 6300 15486 6302 15538
rect 6354 15486 6356 15538
rect 6300 15474 6356 15486
rect 6076 15316 6132 15326
rect 6076 15222 6132 15260
rect 6524 15148 6580 17052
rect 6636 15988 6692 17612
rect 6748 16994 6804 21308
rect 6972 19234 7028 19246
rect 6972 19182 6974 19234
rect 7026 19182 7028 19234
rect 6860 18450 6916 18462
rect 6860 18398 6862 18450
rect 6914 18398 6916 18450
rect 6860 17668 6916 18398
rect 6860 17602 6916 17612
rect 6972 17108 7028 19182
rect 6748 16942 6750 16994
rect 6802 16942 6804 16994
rect 6748 16930 6804 16942
rect 6860 17052 7028 17108
rect 6860 16996 6916 17052
rect 6860 16930 6916 16940
rect 6972 16884 7028 16894
rect 6972 16790 7028 16828
rect 6748 15988 6804 15998
rect 6636 15986 6804 15988
rect 6636 15934 6750 15986
rect 6802 15934 6804 15986
rect 6636 15932 6804 15934
rect 6636 15426 6692 15932
rect 6748 15922 6804 15932
rect 6636 15374 6638 15426
rect 6690 15374 6692 15426
rect 6636 15362 6692 15374
rect 6524 15092 6692 15148
rect 5964 14690 6020 14700
rect 5628 14478 5630 14530
rect 5682 14478 5684 14530
rect 5628 14466 5684 14478
rect 6412 14644 6468 14654
rect 6412 13746 6468 14588
rect 6636 14418 6692 15092
rect 6636 14366 6638 14418
rect 6690 14366 6692 14418
rect 6636 14354 6692 14366
rect 7084 14306 7140 25004
rect 7196 24724 7252 24734
rect 7196 24498 7252 24668
rect 7196 24446 7198 24498
rect 7250 24446 7252 24498
rect 7196 23828 7252 24446
rect 7196 23762 7252 23772
rect 7308 24722 7364 24734
rect 7308 24670 7310 24722
rect 7362 24670 7364 24722
rect 7308 21028 7364 24670
rect 7532 24724 7588 25454
rect 7644 24834 7700 30380
rect 7868 30370 7924 30380
rect 7980 30212 8036 32396
rect 8092 31892 8148 31902
rect 8092 31798 8148 31836
rect 8092 31668 8148 31678
rect 8092 30884 8148 31612
rect 8316 31666 8372 31678
rect 8316 31614 8318 31666
rect 8370 31614 8372 31666
rect 8204 31554 8260 31566
rect 8204 31502 8206 31554
rect 8258 31502 8260 31554
rect 8204 31108 8260 31502
rect 8316 31444 8372 31614
rect 8316 31378 8372 31388
rect 8428 31332 8484 33628
rect 8652 32788 8708 32798
rect 8652 32694 8708 32732
rect 8540 32562 8596 32574
rect 8540 32510 8542 32562
rect 8594 32510 8596 32562
rect 8540 31556 8596 32510
rect 8764 32562 8820 32574
rect 8764 32510 8766 32562
rect 8818 32510 8820 32562
rect 8764 32228 8820 32510
rect 8764 32162 8820 32172
rect 8876 32562 8932 32574
rect 8876 32510 8878 32562
rect 8930 32510 8932 32562
rect 8876 32004 8932 32510
rect 8876 31938 8932 31948
rect 8540 31490 8596 31500
rect 8428 31276 8596 31332
rect 8204 31042 8260 31052
rect 8316 31220 8372 31230
rect 8092 30828 8260 30884
rect 7756 30156 8036 30212
rect 8092 30324 8148 30334
rect 7756 26908 7812 30156
rect 7868 29652 7924 29662
rect 7924 29596 8036 29652
rect 7868 29586 7924 29596
rect 7868 27524 7924 27534
rect 7868 27074 7924 27468
rect 7868 27022 7870 27074
rect 7922 27022 7924 27074
rect 7868 27010 7924 27022
rect 7756 26852 7924 26908
rect 7756 26290 7812 26302
rect 7756 26238 7758 26290
rect 7810 26238 7812 26290
rect 7756 25620 7812 26238
rect 7756 25554 7812 25564
rect 7756 25394 7812 25406
rect 7756 25342 7758 25394
rect 7810 25342 7812 25394
rect 7756 24948 7812 25342
rect 7756 24882 7812 24892
rect 7644 24782 7646 24834
rect 7698 24782 7700 24834
rect 7644 24770 7700 24782
rect 7532 24658 7588 24668
rect 7868 23828 7924 26852
rect 7980 26402 8036 29596
rect 7980 26350 7982 26402
rect 8034 26350 8036 26402
rect 7980 26338 8036 26350
rect 8092 25506 8148 30268
rect 8092 25454 8094 25506
rect 8146 25454 8148 25506
rect 8092 25442 8148 25454
rect 7532 23772 7924 23828
rect 7420 21028 7476 21038
rect 7308 20972 7420 21028
rect 7420 20962 7476 20972
rect 7532 20692 7588 23772
rect 7308 19236 7364 19246
rect 7308 19142 7364 19180
rect 7196 18452 7252 18462
rect 7196 16884 7252 18396
rect 7532 18116 7588 20636
rect 7756 23492 7812 23502
rect 8204 23492 8260 30828
rect 7756 20690 7812 23436
rect 7756 20638 7758 20690
rect 7810 20638 7812 20690
rect 7756 20626 7812 20638
rect 7980 23436 8260 23492
rect 7868 19124 7924 19134
rect 7644 18676 7700 18686
rect 7644 18582 7700 18620
rect 7868 18564 7924 19068
rect 7868 18470 7924 18508
rect 7532 18050 7588 18060
rect 7196 16818 7252 16828
rect 7308 18004 7364 18014
rect 7308 16660 7364 17948
rect 7084 14254 7086 14306
rect 7138 14254 7140 14306
rect 7084 14242 7140 14254
rect 7196 16604 7364 16660
rect 7420 17668 7476 17678
rect 6412 13694 6414 13746
rect 6466 13694 6468 13746
rect 6412 13682 6468 13694
rect 7084 13748 7140 13758
rect 7196 13748 7252 16604
rect 7420 15148 7476 17612
rect 7868 17668 7924 17678
rect 7868 17574 7924 17612
rect 7308 15092 7476 15148
rect 7532 16996 7588 17006
rect 7308 13860 7364 15092
rect 7420 14644 7476 14654
rect 7420 14550 7476 14588
rect 7420 13860 7476 13870
rect 7308 13858 7476 13860
rect 7308 13806 7422 13858
rect 7474 13806 7476 13858
rect 7308 13804 7476 13806
rect 7420 13794 7476 13804
rect 7084 13746 7252 13748
rect 7084 13694 7086 13746
rect 7138 13694 7252 13746
rect 7084 13692 7252 13694
rect 7532 13746 7588 16940
rect 7644 16098 7700 16110
rect 7644 16046 7646 16098
rect 7698 16046 7700 16098
rect 7644 15092 7700 16046
rect 7644 15026 7700 15036
rect 7756 15316 7812 15326
rect 7756 13858 7812 15260
rect 7980 15148 8036 23436
rect 8316 23268 8372 31164
rect 8428 28642 8484 28654
rect 8428 28590 8430 28642
rect 8482 28590 8484 28642
rect 8428 28420 8484 28590
rect 8428 28354 8484 28364
rect 8428 23940 8484 23950
rect 8428 23378 8484 23884
rect 8428 23326 8430 23378
rect 8482 23326 8484 23378
rect 8428 23314 8484 23326
rect 8092 23212 8372 23268
rect 8092 21252 8148 23212
rect 8316 23044 8372 23054
rect 8316 22950 8372 22988
rect 8316 22148 8372 22158
rect 8204 21476 8260 21486
rect 8316 21476 8372 22092
rect 8204 21474 8372 21476
rect 8204 21422 8206 21474
rect 8258 21422 8372 21474
rect 8204 21420 8372 21422
rect 8204 21410 8260 21420
rect 8540 21252 8596 31276
rect 8988 26908 9044 35646
rect 9324 36932 9380 36942
rect 9212 31554 9268 31566
rect 9212 31502 9214 31554
rect 9266 31502 9268 31554
rect 9212 31332 9268 31502
rect 9100 28756 9156 28766
rect 9100 28642 9156 28700
rect 9100 28590 9102 28642
rect 9154 28590 9156 28642
rect 9100 28578 9156 28590
rect 9212 26908 9268 31276
rect 8092 21196 8260 21252
rect 8092 20578 8148 20590
rect 8092 20526 8094 20578
rect 8146 20526 8148 20578
rect 8092 20020 8148 20526
rect 8092 18676 8148 19964
rect 8092 18610 8148 18620
rect 8204 16212 8260 21196
rect 8540 21186 8596 21196
rect 8652 26852 9044 26908
rect 9100 26852 9268 26908
rect 9324 26908 9380 36876
rect 9436 36484 9492 36494
rect 9548 36484 9604 38612
rect 9772 37940 9828 37950
rect 9772 37490 9828 37884
rect 9772 37438 9774 37490
rect 9826 37438 9828 37490
rect 9772 37426 9828 37438
rect 9772 37266 9828 37278
rect 9772 37214 9774 37266
rect 9826 37214 9828 37266
rect 9548 36428 9716 36484
rect 9436 36390 9492 36428
rect 9548 36260 9604 36270
rect 9548 36166 9604 36204
rect 9548 35588 9604 35598
rect 9436 35532 9548 35588
rect 9436 31106 9492 35532
rect 9548 35522 9604 35532
rect 9660 35140 9716 36428
rect 9772 36482 9828 37214
rect 9884 37156 9940 38782
rect 9884 37090 9940 37100
rect 10108 38834 10164 38846
rect 10108 38782 10110 38834
rect 10162 38782 10164 38834
rect 10108 37378 10164 38782
rect 11340 38164 11396 38174
rect 11340 38050 11396 38108
rect 11340 37998 11342 38050
rect 11394 37998 11396 38050
rect 11340 37986 11396 37998
rect 10556 37940 10612 37950
rect 10556 37846 10612 37884
rect 10108 37326 10110 37378
rect 10162 37326 10164 37378
rect 9772 36430 9774 36482
rect 9826 36430 9828 36482
rect 9772 36418 9828 36430
rect 9548 35084 9716 35140
rect 9772 35252 9828 35262
rect 9548 31778 9604 35084
rect 9772 33346 9828 35196
rect 10108 35140 10164 37326
rect 10556 37380 10612 37390
rect 10556 37378 10724 37380
rect 10556 37326 10558 37378
rect 10610 37326 10724 37378
rect 10556 37324 10724 37326
rect 10556 37314 10612 37324
rect 10444 37266 10500 37278
rect 10444 37214 10446 37266
rect 10498 37214 10500 37266
rect 10444 36484 10500 37214
rect 10556 37156 10612 37166
rect 10668 37156 10724 37324
rect 11564 37268 11620 39678
rect 12236 39732 12292 39742
rect 12012 39396 12068 39406
rect 11788 39340 12012 39396
rect 11788 38164 11844 39340
rect 12012 39302 12068 39340
rect 11788 38070 11844 38108
rect 12124 38722 12180 38734
rect 12124 38670 12126 38722
rect 12178 38670 12180 38722
rect 11564 37202 11620 37212
rect 12124 37828 12180 38670
rect 11116 37156 11172 37166
rect 10668 37100 11116 37156
rect 10556 37042 10612 37100
rect 11116 37062 11172 37100
rect 12124 37044 12180 37772
rect 10556 36990 10558 37042
rect 10610 36990 10612 37042
rect 10556 36978 10612 36990
rect 11676 36988 12180 37044
rect 10444 36418 10500 36428
rect 11004 36932 11060 36942
rect 10220 36260 10276 36270
rect 10276 36204 10388 36260
rect 10220 36166 10276 36204
rect 10108 34804 10164 35084
rect 10332 35252 10388 36204
rect 10892 35588 10948 35598
rect 10220 34804 10276 34814
rect 10108 34802 10276 34804
rect 10108 34750 10222 34802
rect 10274 34750 10276 34802
rect 10108 34748 10276 34750
rect 10220 34738 10276 34748
rect 10332 33684 10388 35196
rect 10556 35586 10948 35588
rect 10556 35534 10894 35586
rect 10946 35534 10948 35586
rect 10556 35532 10948 35534
rect 9772 33294 9774 33346
rect 9826 33294 9828 33346
rect 9772 33282 9828 33294
rect 10108 33628 10388 33684
rect 10444 34916 10500 34926
rect 9660 33124 9716 33134
rect 9884 33124 9940 33134
rect 9660 33030 9716 33068
rect 9772 33122 9940 33124
rect 9772 33070 9886 33122
rect 9938 33070 9940 33122
rect 9772 33068 9940 33070
rect 9548 31726 9550 31778
rect 9602 31726 9604 31778
rect 9548 31714 9604 31726
rect 9772 31780 9828 33068
rect 9884 33058 9940 33068
rect 9996 33124 10052 33134
rect 9996 33030 10052 33068
rect 9884 32564 9940 32574
rect 9884 31890 9940 32508
rect 9884 31838 9886 31890
rect 9938 31838 9940 31890
rect 9884 31826 9940 31838
rect 9772 31714 9828 31724
rect 9996 31668 10052 31678
rect 9996 31574 10052 31612
rect 9436 31054 9438 31106
rect 9490 31054 9492 31106
rect 9436 31042 9492 31054
rect 9660 31556 9716 31566
rect 9772 31556 9828 31566
rect 9716 31554 9828 31556
rect 9716 31502 9774 31554
rect 9826 31502 9828 31554
rect 9716 31500 9828 31502
rect 9324 26852 9604 26908
rect 8652 21028 8708 26852
rect 8988 21588 9044 21598
rect 8988 21494 9044 21532
rect 8428 20972 8708 21028
rect 8316 18004 8372 18014
rect 8316 17666 8372 17948
rect 8316 17614 8318 17666
rect 8370 17614 8372 17666
rect 8316 17602 8372 17614
rect 8316 16212 8372 16222
rect 8204 16210 8372 16212
rect 8204 16158 8318 16210
rect 8370 16158 8372 16210
rect 8204 16156 8372 16158
rect 8316 16146 8372 16156
rect 8428 15202 8484 20972
rect 8540 16772 8596 16782
rect 8540 15538 8596 16716
rect 9100 16436 9156 26852
rect 9548 24834 9604 26852
rect 9660 25396 9716 31500
rect 9772 31490 9828 31500
rect 10108 31332 10164 33628
rect 10220 33234 10276 33246
rect 10220 33182 10222 33234
rect 10274 33182 10276 33234
rect 10220 32900 10276 33182
rect 10220 32834 10276 32844
rect 10332 33012 10388 33022
rect 10332 32786 10388 32956
rect 10332 32734 10334 32786
rect 10386 32734 10388 32786
rect 10332 32722 10388 32734
rect 10444 32676 10500 34860
rect 10556 34914 10612 35532
rect 10556 34862 10558 34914
rect 10610 34862 10612 34914
rect 10556 34850 10612 34862
rect 10556 34018 10612 34030
rect 10556 33966 10558 34018
rect 10610 33966 10612 34018
rect 10556 32900 10612 33966
rect 10892 33796 10948 35532
rect 11004 35026 11060 36876
rect 11004 34974 11006 35026
rect 11058 34974 11060 35026
rect 11004 34962 11060 34974
rect 11228 36708 11284 36718
rect 10892 33730 10948 33740
rect 10892 33348 10948 33358
rect 10892 33254 10948 33292
rect 11228 33346 11284 36652
rect 11340 35364 11396 35374
rect 11340 35026 11396 35308
rect 11340 34974 11342 35026
rect 11394 34974 11396 35026
rect 11340 34916 11396 34974
rect 11340 34850 11396 34860
rect 11564 35140 11620 35150
rect 11564 34914 11620 35084
rect 11564 34862 11566 34914
rect 11618 34862 11620 34914
rect 11564 34850 11620 34862
rect 11228 33294 11230 33346
rect 11282 33294 11284 33346
rect 11228 33282 11284 33294
rect 11452 34690 11508 34702
rect 11452 34638 11454 34690
rect 11506 34638 11508 34690
rect 10780 33236 10836 33246
rect 10780 33142 10836 33180
rect 10556 32834 10612 32844
rect 10668 33124 10724 33134
rect 10556 32676 10612 32686
rect 10444 32674 10612 32676
rect 10444 32622 10558 32674
rect 10610 32622 10612 32674
rect 10444 32620 10612 32622
rect 10220 32004 10276 32014
rect 10220 31778 10276 31948
rect 10556 31892 10612 32620
rect 10556 31826 10612 31836
rect 10220 31726 10222 31778
rect 10274 31726 10276 31778
rect 10220 31556 10276 31726
rect 10556 31668 10612 31678
rect 10668 31668 10724 33068
rect 11340 33122 11396 33134
rect 11340 33070 11342 33122
rect 11394 33070 11396 33122
rect 11228 32562 11284 32574
rect 11228 32510 11230 32562
rect 11282 32510 11284 32562
rect 10556 31666 10724 31668
rect 10556 31614 10558 31666
rect 10610 31614 10724 31666
rect 10556 31612 10724 31614
rect 11004 32450 11060 32462
rect 11004 32398 11006 32450
rect 11058 32398 11060 32450
rect 10556 31602 10612 31612
rect 10220 31490 10276 31500
rect 10892 31554 10948 31566
rect 10892 31502 10894 31554
rect 10946 31502 10948 31554
rect 9996 31276 10164 31332
rect 10892 31332 10948 31502
rect 9772 31108 9828 31118
rect 9772 31106 9940 31108
rect 9772 31054 9774 31106
rect 9826 31054 9940 31106
rect 9772 31052 9940 31054
rect 9772 31042 9828 31052
rect 9884 30994 9940 31052
rect 9884 30942 9886 30994
rect 9938 30942 9940 30994
rect 9884 30930 9940 30942
rect 9772 29202 9828 29214
rect 9772 29150 9774 29202
rect 9826 29150 9828 29202
rect 9772 25732 9828 29150
rect 9996 29204 10052 31276
rect 10892 31266 10948 31276
rect 10108 31108 10164 31118
rect 10108 31014 10164 31052
rect 10220 30994 10276 31006
rect 10220 30942 10222 30994
rect 10274 30942 10276 30994
rect 10220 30884 10276 30942
rect 10108 30828 10276 30884
rect 10108 30212 10164 30828
rect 10668 30772 10724 30782
rect 10108 30146 10164 30156
rect 10220 30770 10724 30772
rect 10220 30718 10670 30770
rect 10722 30718 10724 30770
rect 10220 30716 10724 30718
rect 10108 29988 10164 29998
rect 10108 29426 10164 29932
rect 10108 29374 10110 29426
rect 10162 29374 10164 29426
rect 10108 29362 10164 29374
rect 9996 29148 10164 29204
rect 9996 27860 10052 27870
rect 9996 27186 10052 27804
rect 10108 27748 10164 29148
rect 10108 27682 10164 27692
rect 9996 27134 9998 27186
rect 10050 27134 10052 27186
rect 9996 27122 10052 27134
rect 9772 25666 9828 25676
rect 9660 25340 9828 25396
rect 9548 24782 9550 24834
rect 9602 24782 9604 24834
rect 9548 24770 9604 24782
rect 9660 25172 9716 25182
rect 9660 23940 9716 25116
rect 9772 24722 9828 25340
rect 9996 24836 10052 24846
rect 9996 24742 10052 24780
rect 9772 24670 9774 24722
rect 9826 24670 9828 24722
rect 9772 24164 9828 24670
rect 10108 24722 10164 24734
rect 10108 24670 10110 24722
rect 10162 24670 10164 24722
rect 9884 24612 9940 24622
rect 9884 24518 9940 24556
rect 10108 24388 10164 24670
rect 10108 24322 10164 24332
rect 9772 24108 10052 24164
rect 9884 23940 9940 23950
rect 9660 23938 9940 23940
rect 9660 23886 9886 23938
rect 9938 23886 9940 23938
rect 9660 23884 9940 23886
rect 9772 23716 9828 23726
rect 9772 23622 9828 23660
rect 9324 22484 9380 22494
rect 9884 22484 9940 23884
rect 9996 23492 10052 24108
rect 10108 23940 10164 23950
rect 10108 23846 10164 23884
rect 10220 23604 10276 30716
rect 10668 30706 10724 30716
rect 11004 30660 11060 32398
rect 11228 32340 11284 32510
rect 11228 32274 11284 32284
rect 11340 31892 11396 33070
rect 11452 32116 11508 34638
rect 11452 32050 11508 32060
rect 11564 33346 11620 33358
rect 11564 33294 11566 33346
rect 11618 33294 11620 33346
rect 11004 30594 11060 30604
rect 11228 31836 11396 31892
rect 10332 30548 10388 30558
rect 10332 29426 10388 30492
rect 11228 30548 11284 31836
rect 11340 31668 11396 31678
rect 11340 31574 11396 31612
rect 11564 31444 11620 33294
rect 11676 32562 11732 36988
rect 11900 35700 11956 35710
rect 12124 35700 12180 35710
rect 11900 35698 12124 35700
rect 11900 35646 11902 35698
rect 11954 35646 12124 35698
rect 11900 35644 12124 35646
rect 11900 35634 11956 35644
rect 12124 35634 12180 35644
rect 11788 34914 11844 34926
rect 11788 34862 11790 34914
rect 11842 34862 11844 34914
rect 11788 32788 11844 34862
rect 12012 34692 12068 34702
rect 12012 34598 12068 34636
rect 12124 34690 12180 34702
rect 12124 34638 12126 34690
rect 12178 34638 12180 34690
rect 11900 33572 11956 33582
rect 11900 33458 11956 33516
rect 11900 33406 11902 33458
rect 11954 33406 11956 33458
rect 11900 33394 11956 33406
rect 12124 33124 12180 34638
rect 12124 33058 12180 33068
rect 11788 32732 11956 32788
rect 11676 32510 11678 32562
rect 11730 32510 11732 32562
rect 11676 32498 11732 32510
rect 11900 32340 11956 32732
rect 12236 32340 12292 39676
rect 12572 38500 12628 38510
rect 12460 38444 12572 38500
rect 12348 37268 12404 37278
rect 12348 37174 12404 37212
rect 12348 35924 12404 35934
rect 12460 35924 12516 38444
rect 12572 38434 12628 38444
rect 12348 35922 12516 35924
rect 12348 35870 12350 35922
rect 12402 35870 12516 35922
rect 12348 35868 12516 35870
rect 12572 37378 12628 37390
rect 12572 37326 12574 37378
rect 12626 37326 12628 37378
rect 12348 35858 12404 35868
rect 12572 35364 12628 37326
rect 12572 35298 12628 35308
rect 12348 33572 12404 33582
rect 12348 33458 12404 33516
rect 12348 33406 12350 33458
rect 12402 33406 12404 33458
rect 12348 33394 12404 33406
rect 12572 33124 12628 33134
rect 12572 32674 12628 33068
rect 12572 32622 12574 32674
rect 12626 32622 12628 32674
rect 12572 32610 12628 32622
rect 11900 32274 11956 32284
rect 12124 32284 12292 32340
rect 12348 32562 12404 32574
rect 12348 32510 12350 32562
rect 12402 32510 12404 32562
rect 11564 31378 11620 31388
rect 11676 32004 11732 32014
rect 11676 31332 11732 31948
rect 11676 31266 11732 31276
rect 11228 30482 11284 30492
rect 11676 30770 11732 30782
rect 11676 30718 11678 30770
rect 11730 30718 11732 30770
rect 11676 30324 11732 30718
rect 12012 30772 12068 30782
rect 12012 30678 12068 30716
rect 11788 30436 11844 30446
rect 11788 30342 11844 30380
rect 11676 30258 11732 30268
rect 11452 30212 11508 30222
rect 11116 30100 11172 30138
rect 11340 30100 11396 30110
rect 11172 30098 11396 30100
rect 11172 30046 11342 30098
rect 11394 30046 11396 30098
rect 11172 30044 11396 30046
rect 11116 30034 11172 30044
rect 11340 30034 11396 30044
rect 11452 29876 11508 30156
rect 12012 30212 12068 30222
rect 12124 30212 12180 32284
rect 12236 32116 12292 32126
rect 12236 30994 12292 32060
rect 12236 30942 12238 30994
rect 12290 30942 12292 30994
rect 12236 30930 12292 30942
rect 12348 30996 12404 32510
rect 12572 32340 12628 32350
rect 12348 30930 12404 30940
rect 12460 31444 12516 31454
rect 12236 30212 12292 30222
rect 12124 30210 12292 30212
rect 12124 30158 12238 30210
rect 12290 30158 12292 30210
rect 12124 30156 12292 30158
rect 12012 30118 12068 30156
rect 12236 30146 12292 30156
rect 11452 29810 11508 29820
rect 11564 30098 11620 30110
rect 11564 30046 11566 30098
rect 11618 30046 11620 30098
rect 10332 29374 10334 29426
rect 10386 29374 10388 29426
rect 10332 29362 10388 29374
rect 11564 29092 11620 30046
rect 11676 29988 11732 29998
rect 11676 29894 11732 29932
rect 11228 29036 11620 29092
rect 11788 29314 11844 29326
rect 11788 29262 11790 29314
rect 11842 29262 11844 29314
rect 10332 28644 10388 28654
rect 10332 28550 10388 28588
rect 10444 28644 10500 28654
rect 10892 28644 10948 28654
rect 11116 28644 11172 28654
rect 10444 28642 10948 28644
rect 10444 28590 10446 28642
rect 10498 28590 10894 28642
rect 10946 28590 10948 28642
rect 10444 28588 10948 28590
rect 10444 28578 10500 28588
rect 10892 28578 10948 28588
rect 11004 28642 11172 28644
rect 11004 28590 11118 28642
rect 11170 28590 11172 28642
rect 11004 28588 11172 28590
rect 10780 28420 10836 28430
rect 10780 28326 10836 28364
rect 10780 27972 10836 27982
rect 11004 27972 11060 28588
rect 11116 28578 11172 28588
rect 10780 27970 11060 27972
rect 10780 27918 10782 27970
rect 10834 27918 11060 27970
rect 10780 27916 11060 27918
rect 10556 27858 10612 27870
rect 10556 27806 10558 27858
rect 10610 27806 10612 27858
rect 10556 27524 10612 27806
rect 10556 27458 10612 27468
rect 10332 25732 10388 25742
rect 10388 25676 10500 25732
rect 10332 25666 10388 25676
rect 10332 23938 10388 23950
rect 10332 23886 10334 23938
rect 10386 23886 10388 23938
rect 10332 23828 10388 23886
rect 10332 23762 10388 23772
rect 10444 23716 10500 25676
rect 10556 25284 10612 25294
rect 10780 25284 10836 27916
rect 11116 27858 11172 27870
rect 11116 27806 11118 27858
rect 11170 27806 11172 27858
rect 11004 27748 11060 27758
rect 11004 26908 11060 27692
rect 11116 27188 11172 27806
rect 11116 27122 11172 27132
rect 11228 27076 11284 29036
rect 11340 28868 11396 28878
rect 11340 28532 11396 28812
rect 11788 28756 11844 29262
rect 11788 28690 11844 28700
rect 11340 28466 11396 28476
rect 11452 28642 11508 28654
rect 11452 28590 11454 28642
rect 11506 28590 11508 28642
rect 11340 27748 11396 27758
rect 11340 27654 11396 27692
rect 11452 27188 11508 28590
rect 11900 28644 11956 28654
rect 11900 28550 11956 28588
rect 12236 28532 12292 28542
rect 11676 28084 11732 28094
rect 11676 28082 12068 28084
rect 11676 28030 11678 28082
rect 11730 28030 12068 28082
rect 11676 28028 12068 28030
rect 11676 28018 11732 28028
rect 11788 27858 11844 27870
rect 11788 27806 11790 27858
rect 11842 27806 11844 27858
rect 11564 27636 11620 27646
rect 11564 27542 11620 27580
rect 11788 27412 11844 27806
rect 11788 27346 11844 27356
rect 12012 27188 12068 28028
rect 12124 27860 12180 27870
rect 12124 27766 12180 27804
rect 12236 27636 12292 28476
rect 12460 28196 12516 31388
rect 12572 30212 12628 32284
rect 12684 30996 12740 40462
rect 12908 39396 12964 39406
rect 12908 39302 12964 39340
rect 13020 38668 13076 40908
rect 13132 40626 13188 41132
rect 13468 40964 13524 40974
rect 13468 40962 13748 40964
rect 13468 40910 13470 40962
rect 13522 40910 13748 40962
rect 13468 40908 13748 40910
rect 13468 40898 13524 40908
rect 13132 40574 13134 40626
rect 13186 40574 13188 40626
rect 13132 40562 13188 40574
rect 13468 39732 13524 39742
rect 13468 39638 13524 39676
rect 13020 38612 13300 38668
rect 12908 37826 12964 37838
rect 12908 37774 12910 37826
rect 12962 37774 12964 37826
rect 12908 37716 12964 37774
rect 12908 37650 12964 37660
rect 13020 37154 13076 37166
rect 13020 37102 13022 37154
rect 13074 37102 13076 37154
rect 12796 35810 12852 35822
rect 12796 35758 12798 35810
rect 12850 35758 12852 35810
rect 12796 35700 12852 35758
rect 13020 35812 13076 37102
rect 13020 35746 13076 35756
rect 12796 35364 12852 35644
rect 13020 35588 13076 35598
rect 13020 35494 13076 35532
rect 12796 35308 13076 35364
rect 12796 34692 12852 34702
rect 12852 34636 12964 34692
rect 12796 34598 12852 34636
rect 12796 34132 12852 34142
rect 12796 34038 12852 34076
rect 12908 33796 12964 34636
rect 12908 33730 12964 33740
rect 12908 33124 12964 33134
rect 13020 33124 13076 35308
rect 13244 33796 13300 38612
rect 13356 37266 13412 37278
rect 13356 37214 13358 37266
rect 13410 37214 13412 37266
rect 13356 35698 13412 37214
rect 13356 35646 13358 35698
rect 13410 35646 13412 35698
rect 13356 34692 13412 35646
rect 13356 34626 13412 34636
rect 13468 35812 13524 35822
rect 13356 34020 13412 34030
rect 13356 33926 13412 33964
rect 13244 33740 13412 33796
rect 12908 33122 13076 33124
rect 12908 33070 12910 33122
rect 12962 33070 13076 33122
rect 12908 33068 13076 33070
rect 12908 31220 12964 33068
rect 13132 32450 13188 32462
rect 13132 32398 13134 32450
rect 13186 32398 13188 32450
rect 13132 32004 13188 32398
rect 13132 31938 13188 31948
rect 12908 31154 12964 31164
rect 12684 30940 13300 30996
rect 12572 30146 12628 30156
rect 12796 28756 12852 28766
rect 12460 28140 12628 28196
rect 12460 27972 12516 27982
rect 12460 27878 12516 27916
rect 12348 27748 12404 27758
rect 12348 27654 12404 27692
rect 12236 27570 12292 27580
rect 12124 27188 12180 27198
rect 11452 27122 11508 27132
rect 11564 27132 11788 27188
rect 12012 27186 12180 27188
rect 12012 27134 12126 27186
rect 12178 27134 12180 27186
rect 12012 27132 12180 27134
rect 11564 27076 11620 27132
rect 11228 27020 11396 27076
rect 11340 26908 11396 27020
rect 11732 27076 11788 27132
rect 12124 27122 12180 27132
rect 11732 27020 11956 27076
rect 12572 27020 12628 28140
rect 11564 27010 11620 27020
rect 11900 26908 11956 27020
rect 12348 26964 12628 27020
rect 12796 27074 12852 28700
rect 12908 28532 12964 28542
rect 12908 28082 12964 28476
rect 12908 28030 12910 28082
rect 12962 28030 12964 28082
rect 12908 27748 12964 28030
rect 12908 27682 12964 27692
rect 12908 27412 12964 27422
rect 12964 27356 13188 27412
rect 12908 27346 12964 27356
rect 12796 27022 12798 27074
rect 12850 27022 12852 27074
rect 11004 26852 11284 26908
rect 11340 26852 11844 26908
rect 11900 26852 12068 26908
rect 10556 25282 10724 25284
rect 10556 25230 10558 25282
rect 10610 25230 10724 25282
rect 10556 25228 10724 25230
rect 10556 25218 10612 25228
rect 10556 24948 10612 24958
rect 10556 24854 10612 24892
rect 10668 24836 10724 25228
rect 10780 25218 10836 25228
rect 10780 24836 10836 24846
rect 10668 24780 10780 24836
rect 10780 24770 10836 24780
rect 10892 24724 10948 24734
rect 10892 24630 10948 24668
rect 11116 24612 11172 24622
rect 11116 24518 11172 24556
rect 11116 24052 11172 24062
rect 10556 24050 11172 24052
rect 10556 23998 11118 24050
rect 11170 23998 11172 24050
rect 10556 23996 11172 23998
rect 10556 23938 10612 23996
rect 11116 23986 11172 23996
rect 10556 23886 10558 23938
rect 10610 23886 10612 23938
rect 10556 23874 10612 23886
rect 10780 23826 10836 23838
rect 10780 23774 10782 23826
rect 10834 23774 10836 23826
rect 10780 23716 10836 23774
rect 10444 23660 10836 23716
rect 10220 23548 10836 23604
rect 9996 23426 10052 23436
rect 10444 23380 10500 23390
rect 10220 23324 10444 23380
rect 10108 22708 10164 22718
rect 9380 22428 9716 22484
rect 9324 22390 9380 22428
rect 9660 22370 9716 22428
rect 9940 22428 10052 22484
rect 9884 22418 9940 22428
rect 9660 22318 9662 22370
rect 9714 22318 9716 22370
rect 9660 22306 9716 22318
rect 9884 22146 9940 22158
rect 9884 22094 9886 22146
rect 9938 22094 9940 22146
rect 9548 20020 9604 20030
rect 9548 19926 9604 19964
rect 9884 20020 9940 22094
rect 9996 21698 10052 22428
rect 10108 22370 10164 22652
rect 10220 22482 10276 23324
rect 10444 23314 10500 23324
rect 10668 23042 10724 23054
rect 10668 22990 10670 23042
rect 10722 22990 10724 23042
rect 10668 22708 10724 22990
rect 10668 22642 10724 22652
rect 10220 22430 10222 22482
rect 10274 22430 10276 22482
rect 10220 22418 10276 22430
rect 10668 22484 10724 22494
rect 10108 22318 10110 22370
rect 10162 22318 10164 22370
rect 10108 22306 10164 22318
rect 10332 22372 10388 22382
rect 10332 22278 10388 22316
rect 10668 22370 10724 22428
rect 10668 22318 10670 22370
rect 10722 22318 10724 22370
rect 10668 22306 10724 22318
rect 10556 22148 10612 22158
rect 10556 22054 10612 22092
rect 10108 21812 10164 21822
rect 10108 21810 10388 21812
rect 10108 21758 10110 21810
rect 10162 21758 10388 21810
rect 10108 21756 10388 21758
rect 10108 21746 10164 21756
rect 9996 21646 9998 21698
rect 10050 21646 10052 21698
rect 9996 21634 10052 21646
rect 10220 21476 10276 21486
rect 10220 21382 10276 21420
rect 9884 19954 9940 19964
rect 9996 21252 10052 21262
rect 9996 18788 10052 21196
rect 10332 20916 10388 21756
rect 10780 21700 10836 23548
rect 11116 22484 11172 22494
rect 11116 22390 11172 22428
rect 10892 22370 10948 22382
rect 10892 22318 10894 22370
rect 10946 22318 10948 22370
rect 10892 22036 10948 22318
rect 11228 22148 11284 26852
rect 11564 26290 11620 26302
rect 11564 26238 11566 26290
rect 11618 26238 11620 26290
rect 11340 26180 11396 26190
rect 11564 26180 11620 26238
rect 11788 26292 11844 26852
rect 11900 26292 11956 26302
rect 11788 26290 11956 26292
rect 11788 26238 11902 26290
rect 11954 26238 11956 26290
rect 11788 26236 11956 26238
rect 11340 26178 11620 26180
rect 11340 26126 11342 26178
rect 11394 26126 11620 26178
rect 11340 26124 11620 26126
rect 11340 22596 11396 26124
rect 11564 25956 11620 25966
rect 11452 23938 11508 23950
rect 11452 23886 11454 23938
rect 11506 23886 11508 23938
rect 11452 23380 11508 23886
rect 11452 23314 11508 23324
rect 11340 22530 11396 22540
rect 11340 22260 11396 22270
rect 11340 22258 11508 22260
rect 11340 22206 11342 22258
rect 11394 22206 11508 22258
rect 11340 22204 11508 22206
rect 11340 22194 11396 22204
rect 11228 22082 11284 22092
rect 10892 21970 10948 21980
rect 11340 22036 11396 22046
rect 11340 21810 11396 21980
rect 11340 21758 11342 21810
rect 11394 21758 11396 21810
rect 11340 21746 11396 21758
rect 10892 21700 10948 21710
rect 10780 21698 10948 21700
rect 10780 21646 10894 21698
rect 10946 21646 10948 21698
rect 10780 21644 10948 21646
rect 10892 21634 10948 21644
rect 10668 21586 10724 21598
rect 10668 21534 10670 21586
rect 10722 21534 10724 21586
rect 10444 21364 10500 21374
rect 10444 21362 10612 21364
rect 10444 21310 10446 21362
rect 10498 21310 10612 21362
rect 10444 21308 10612 21310
rect 10444 21298 10500 21308
rect 10556 21252 10612 21308
rect 10556 21186 10612 21196
rect 10332 20850 10388 20860
rect 10108 20692 10164 20702
rect 10108 20598 10164 20636
rect 10444 20244 10500 20254
rect 10668 20244 10724 21534
rect 11228 21474 11284 21486
rect 11228 21422 11230 21474
rect 11282 21422 11284 21474
rect 11228 21364 11284 21422
rect 11228 21298 11284 21308
rect 10780 20692 10836 20702
rect 10836 20636 11060 20692
rect 10780 20626 10836 20636
rect 10444 20242 10724 20244
rect 10444 20190 10446 20242
rect 10498 20190 10724 20242
rect 10444 20188 10724 20190
rect 10444 20178 10500 20188
rect 10108 20020 10164 20030
rect 10108 19926 10164 19964
rect 11004 20020 11060 20636
rect 11452 20580 11508 22204
rect 11452 20514 11508 20524
rect 11564 20244 11620 25900
rect 11900 25508 11956 26236
rect 12012 25956 12068 26852
rect 12124 26404 12180 26414
rect 12124 26290 12180 26348
rect 12124 26238 12126 26290
rect 12178 26238 12180 26290
rect 12124 26226 12180 26238
rect 12348 26290 12404 26964
rect 12796 26908 12852 27022
rect 12796 26852 12964 26908
rect 12348 26238 12350 26290
rect 12402 26238 12404 26290
rect 12348 26226 12404 26238
rect 12572 26290 12628 26302
rect 12572 26238 12574 26290
rect 12626 26238 12628 26290
rect 12012 25890 12068 25900
rect 12460 26178 12516 26190
rect 12460 26126 12462 26178
rect 12514 26126 12516 26178
rect 12460 25732 12516 26126
rect 12572 26180 12628 26238
rect 12572 26114 12628 26124
rect 12348 25676 12516 25732
rect 12572 25956 12628 25966
rect 11900 25452 12068 25508
rect 11900 25284 11956 25294
rect 11788 25282 11956 25284
rect 11788 25230 11902 25282
rect 11954 25230 11956 25282
rect 11788 25228 11956 25230
rect 11676 24612 11732 24622
rect 11676 24050 11732 24556
rect 11676 23998 11678 24050
rect 11730 23998 11732 24050
rect 11676 23986 11732 23998
rect 11788 23716 11844 25228
rect 11900 25218 11956 25228
rect 12012 24948 12068 25452
rect 12348 25506 12404 25676
rect 12572 25620 12628 25900
rect 12348 25454 12350 25506
rect 12402 25454 12404 25506
rect 12348 25442 12404 25454
rect 12460 25564 12628 25620
rect 12460 25506 12516 25564
rect 12460 25454 12462 25506
rect 12514 25454 12516 25506
rect 12460 25442 12516 25454
rect 12572 25394 12628 25406
rect 12572 25342 12574 25394
rect 12626 25342 12628 25394
rect 12572 25060 12628 25342
rect 12572 24994 12628 25004
rect 12796 25172 12852 25182
rect 12684 24948 12740 24958
rect 12012 24892 12404 24948
rect 12236 24722 12292 24734
rect 12236 24670 12238 24722
rect 12290 24670 12292 24722
rect 11900 24612 11956 24622
rect 12236 24612 12292 24670
rect 12348 24724 12404 24892
rect 12684 24854 12740 24892
rect 12796 24946 12852 25116
rect 12796 24894 12798 24946
rect 12850 24894 12852 24946
rect 12796 24882 12852 24894
rect 12460 24724 12516 24734
rect 12348 24722 12516 24724
rect 12348 24670 12462 24722
rect 12514 24670 12516 24722
rect 12348 24668 12516 24670
rect 11900 24610 12292 24612
rect 11900 24558 11902 24610
rect 11954 24558 12292 24610
rect 11900 24556 12292 24558
rect 11900 24546 11956 24556
rect 11676 23660 11844 23716
rect 11676 22370 11732 23660
rect 12236 23156 12292 24556
rect 12236 23090 12292 23100
rect 12012 23044 12068 23054
rect 12012 22484 12068 22988
rect 11676 22318 11678 22370
rect 11730 22318 11732 22370
rect 11676 22306 11732 22318
rect 11788 22428 12012 22484
rect 11788 21810 11844 22428
rect 12012 22390 12068 22428
rect 11788 21758 11790 21810
rect 11842 21758 11844 21810
rect 11788 21252 11844 21758
rect 11788 21186 11844 21196
rect 11564 20178 11620 20188
rect 11788 21028 11844 21038
rect 11676 20020 11732 20030
rect 11004 20018 11284 20020
rect 11004 19966 11006 20018
rect 11058 19966 11284 20018
rect 11004 19964 11284 19966
rect 11004 19954 11060 19964
rect 10780 19794 10836 19806
rect 10780 19742 10782 19794
rect 10834 19742 10836 19794
rect 10108 19236 10164 19246
rect 10108 19234 10276 19236
rect 10108 19182 10110 19234
rect 10162 19182 10276 19234
rect 10108 19180 10276 19182
rect 10108 19170 10164 19180
rect 9772 18732 10164 18788
rect 9660 18676 9716 18686
rect 9548 18450 9604 18462
rect 9548 18398 9550 18450
rect 9602 18398 9604 18450
rect 9548 18228 9604 18398
rect 9548 18162 9604 18172
rect 9100 16370 9156 16380
rect 9548 18004 9604 18014
rect 8764 15988 8820 15998
rect 8540 15486 8542 15538
rect 8594 15486 8596 15538
rect 8540 15474 8596 15486
rect 8652 15986 8820 15988
rect 8652 15934 8766 15986
rect 8818 15934 8820 15986
rect 8652 15932 8820 15934
rect 8428 15150 8430 15202
rect 8482 15150 8484 15202
rect 7980 15092 8148 15148
rect 8428 15138 8484 15150
rect 7756 13806 7758 13858
rect 7810 13806 7812 13858
rect 7756 13794 7812 13806
rect 7532 13694 7534 13746
rect 7586 13694 7588 13746
rect 7084 13682 7140 13692
rect 7532 13682 7588 13694
rect 4396 12460 5012 12516
rect 5740 13412 5796 13422
rect 4396 12402 4452 12460
rect 4396 12350 4398 12402
rect 4450 12350 4452 12402
rect 4396 12338 4452 12350
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4844 11396 4900 12460
rect 5404 12404 5460 12414
rect 5740 12404 5796 13356
rect 5852 13076 5908 13086
rect 6636 13076 6692 13086
rect 7084 13076 7140 13086
rect 5908 13020 6244 13076
rect 5852 12982 5908 13020
rect 5404 12402 5796 12404
rect 5404 12350 5406 12402
rect 5458 12350 5742 12402
rect 5794 12350 5796 12402
rect 5404 12348 5796 12350
rect 5404 12338 5460 12348
rect 5740 12338 5796 12348
rect 5852 12852 5908 12862
rect 5852 12290 5908 12796
rect 5852 12238 5854 12290
rect 5906 12238 5908 12290
rect 5516 12178 5572 12190
rect 5516 12126 5518 12178
rect 5570 12126 5572 12178
rect 4956 12066 5012 12078
rect 4956 12014 4958 12066
rect 5010 12014 5012 12066
rect 4956 11844 5012 12014
rect 5516 11956 5572 12126
rect 5516 11890 5572 11900
rect 5740 12068 5796 12078
rect 4956 11732 5012 11788
rect 4956 11676 5124 11732
rect 5068 11506 5124 11676
rect 5068 11454 5070 11506
rect 5122 11454 5124 11506
rect 5068 11442 5124 11454
rect 5628 11396 5684 11406
rect 4844 10612 4900 11340
rect 5516 11394 5684 11396
rect 5516 11342 5630 11394
rect 5682 11342 5684 11394
rect 5516 11340 5684 11342
rect 5516 10834 5572 11340
rect 5628 11330 5684 11340
rect 5740 10836 5796 12012
rect 5852 11844 5908 12238
rect 6188 12290 6244 13020
rect 6692 13020 6804 13076
rect 6636 12982 6692 13020
rect 6300 12404 6356 12414
rect 6300 12310 6356 12348
rect 6188 12238 6190 12290
rect 6242 12238 6244 12290
rect 6188 12068 6244 12238
rect 6188 12002 6244 12012
rect 6076 11956 6132 11966
rect 5852 11732 6020 11788
rect 5852 11172 5908 11182
rect 5852 11078 5908 11116
rect 5516 10782 5518 10834
rect 5570 10782 5572 10834
rect 5516 10770 5572 10782
rect 5628 10834 5796 10836
rect 5628 10782 5742 10834
rect 5794 10782 5796 10834
rect 5628 10780 5796 10782
rect 5628 10612 5684 10780
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4844 10164 4900 10556
rect 5068 10556 5684 10612
rect 5068 10498 5124 10556
rect 5068 10446 5070 10498
rect 5122 10446 5124 10498
rect 5068 10434 5124 10446
rect 4844 10108 5124 10164
rect 4284 9874 4340 9884
rect 5068 9938 5124 10108
rect 5068 9886 5070 9938
rect 5122 9886 5124 9938
rect 5068 9874 5124 9886
rect 5740 9940 5796 10780
rect 5852 10724 5908 10734
rect 5852 10630 5908 10668
rect 5852 9940 5908 9950
rect 5740 9938 5908 9940
rect 5740 9886 5854 9938
rect 5906 9886 5908 9938
rect 5740 9884 5908 9886
rect 5852 9874 5908 9884
rect 5964 9604 6020 11732
rect 6076 11394 6132 11900
rect 6300 11956 6356 11966
rect 6300 11954 6468 11956
rect 6300 11902 6302 11954
rect 6354 11902 6468 11954
rect 6300 11900 6468 11902
rect 6300 11890 6356 11900
rect 6076 11342 6078 11394
rect 6130 11342 6132 11394
rect 6076 11330 6132 11342
rect 6188 11284 6244 11294
rect 6188 10836 6244 11228
rect 6300 11282 6356 11294
rect 6300 11230 6302 11282
rect 6354 11230 6356 11282
rect 6300 11172 6356 11230
rect 6300 11106 6356 11116
rect 6300 10836 6356 10846
rect 6188 10834 6356 10836
rect 6188 10782 6302 10834
rect 6354 10782 6356 10834
rect 6188 10780 6356 10782
rect 6300 10770 6356 10780
rect 6188 10610 6244 10622
rect 6188 10558 6190 10610
rect 6242 10558 6244 10610
rect 6188 9826 6244 10558
rect 6412 9940 6468 11900
rect 6748 11506 6804 13020
rect 7140 13020 7252 13076
rect 7084 13010 7140 13020
rect 7084 12740 7140 12750
rect 6748 11454 6750 11506
rect 6802 11454 6804 11506
rect 6636 11396 6692 11406
rect 6524 10612 6580 10622
rect 6524 10518 6580 10556
rect 6188 9774 6190 9826
rect 6242 9774 6244 9826
rect 6188 9762 6244 9774
rect 6300 9884 6468 9940
rect 6524 10388 6580 10398
rect 5964 9268 6020 9548
rect 6076 9268 6132 9278
rect 5964 9266 6132 9268
rect 5964 9214 6078 9266
rect 6130 9214 6132 9266
rect 5964 9212 6132 9214
rect 6076 9202 6132 9212
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 6300 8428 6356 9884
rect 6524 9826 6580 10332
rect 6524 9774 6526 9826
rect 6578 9774 6580 9826
rect 6524 9762 6580 9774
rect 6412 9604 6468 9614
rect 6412 9510 6468 9548
rect 4172 8372 4900 8428
rect 6300 8372 6468 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 3276 6066 3332 6076
rect 2044 5404 2660 5460
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 2044 5010 2100 5404
rect 2044 4958 2046 5010
rect 2098 4958 2100 5010
rect 2044 4946 2100 4958
rect 2492 5122 2548 5134
rect 2492 5070 2494 5122
rect 2546 5070 2548 5122
rect 2492 4900 2548 5070
rect 2492 4834 2548 4844
rect 2156 4228 2212 4238
rect 1932 4226 2212 4228
rect 1932 4174 2158 4226
rect 2210 4174 2212 4226
rect 1932 4172 2212 4174
rect 2156 4162 2212 4172
rect 4172 4116 4228 4126
rect 4172 4114 4340 4116
rect 4172 4062 4174 4114
rect 4226 4062 4340 4114
rect 4172 4060 4340 4062
rect 4172 4050 4228 4060
rect 1820 3390 1822 3442
rect 1874 3390 1876 3442
rect 1820 2996 1876 3390
rect 1820 2930 1876 2940
rect 2716 3666 2772 3678
rect 2716 3614 2718 3666
rect 2770 3614 2772 3666
rect 2716 800 2772 3614
rect 4284 980 4340 4060
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4844 3554 4900 8372
rect 6076 4340 6132 4350
rect 6076 4246 6132 4284
rect 6412 4338 6468 8372
rect 6636 6692 6692 11340
rect 6748 10836 6804 11454
rect 6972 12684 7084 12740
rect 6972 12180 7028 12684
rect 7084 12646 7140 12684
rect 7084 12404 7140 12414
rect 7196 12404 7252 13020
rect 7084 12402 7252 12404
rect 7084 12350 7086 12402
rect 7138 12350 7252 12402
rect 7084 12348 7252 12350
rect 7756 12404 7812 12414
rect 7084 12338 7140 12348
rect 7756 12310 7812 12348
rect 6972 11396 7028 12124
rect 7196 12178 7252 12190
rect 7196 12126 7198 12178
rect 7250 12126 7252 12178
rect 7084 11956 7140 11966
rect 7196 11956 7252 12126
rect 7420 11956 7476 11966
rect 7196 11900 7420 11956
rect 7084 11862 7140 11900
rect 7196 11620 7252 11630
rect 7084 11396 7140 11406
rect 6972 11394 7140 11396
rect 6972 11342 7086 11394
rect 7138 11342 7140 11394
rect 6972 11340 7140 11342
rect 7084 11330 7140 11340
rect 6748 10770 6804 10780
rect 6860 11172 6916 11182
rect 6748 10612 6804 10622
rect 6860 10612 6916 11116
rect 7196 10948 7252 11564
rect 7196 10834 7252 10892
rect 7196 10782 7198 10834
rect 7250 10782 7252 10834
rect 7196 10770 7252 10782
rect 7308 10722 7364 11900
rect 7420 11890 7476 11900
rect 8092 11732 8148 15092
rect 8652 14644 8708 15932
rect 8764 15922 8820 15932
rect 8764 15202 8820 15214
rect 8764 15150 8766 15202
rect 8818 15150 8820 15202
rect 8764 14756 8820 15150
rect 8764 14690 8820 14700
rect 8652 14578 8708 14588
rect 9548 13412 9604 17948
rect 9660 17778 9716 18620
rect 9660 17726 9662 17778
rect 9714 17726 9716 17778
rect 9660 17714 9716 17726
rect 9660 17108 9716 17118
rect 9660 16770 9716 17052
rect 9660 16718 9662 16770
rect 9714 16718 9716 16770
rect 9660 16706 9716 16718
rect 9772 16660 9828 18732
rect 9996 18564 10052 18574
rect 9996 17556 10052 18508
rect 10108 18450 10164 18732
rect 10108 18398 10110 18450
rect 10162 18398 10164 18450
rect 10108 18386 10164 18398
rect 10220 18228 10276 19180
rect 10556 19234 10612 19246
rect 10556 19182 10558 19234
rect 10610 19182 10612 19234
rect 10556 19012 10612 19182
rect 10556 18946 10612 18956
rect 10220 18162 10276 18172
rect 10108 17556 10164 17566
rect 9996 17554 10164 17556
rect 9996 17502 10110 17554
rect 10162 17502 10164 17554
rect 9996 17500 10164 17502
rect 9884 16884 9940 16894
rect 9884 16790 9940 16828
rect 10108 16882 10164 17500
rect 10108 16830 10110 16882
rect 10162 16830 10164 16882
rect 10108 16818 10164 16830
rect 10556 16660 10612 16670
rect 9772 16604 9940 16660
rect 9772 15316 9828 15326
rect 9772 15222 9828 15260
rect 9884 15092 9940 16604
rect 10556 16566 10612 16604
rect 10780 16212 10836 19742
rect 11228 19236 11284 19964
rect 10892 19234 11284 19236
rect 10892 19182 11230 19234
rect 11282 19182 11284 19234
rect 10892 19180 11284 19182
rect 10892 18674 10948 19180
rect 11228 19170 11284 19180
rect 11564 19234 11620 19246
rect 11564 19182 11566 19234
rect 11618 19182 11620 19234
rect 11564 19124 11620 19182
rect 11564 19058 11620 19068
rect 10892 18622 10894 18674
rect 10946 18622 10948 18674
rect 10892 18610 10948 18622
rect 11564 18900 11620 18910
rect 11452 18564 11508 18574
rect 11452 18470 11508 18508
rect 11452 17666 11508 17678
rect 11452 17614 11454 17666
rect 11506 17614 11508 17666
rect 10780 16146 10836 16156
rect 10892 16548 10948 16558
rect 10892 16098 10948 16492
rect 10892 16046 10894 16098
rect 10946 16046 10948 16098
rect 10892 16034 10948 16046
rect 11116 16324 11172 16334
rect 11116 15986 11172 16268
rect 11116 15934 11118 15986
rect 11170 15934 11172 15986
rect 11116 15540 11172 15934
rect 11228 16212 11284 16222
rect 11228 15540 11284 16156
rect 11452 15988 11508 17614
rect 11564 17556 11620 18844
rect 11676 18450 11732 19964
rect 11676 18398 11678 18450
rect 11730 18398 11732 18450
rect 11676 18386 11732 18398
rect 11676 17556 11732 17566
rect 11564 17554 11732 17556
rect 11564 17502 11678 17554
rect 11730 17502 11732 17554
rect 11564 17500 11732 17502
rect 11676 17490 11732 17500
rect 11788 17108 11844 20972
rect 12012 20244 12068 20254
rect 12012 20150 12068 20188
rect 12348 19796 12404 19806
rect 12236 19346 12292 19358
rect 12236 19294 12238 19346
rect 12290 19294 12292 19346
rect 12236 19236 12292 19294
rect 12236 19170 12292 19180
rect 12348 19234 12404 19740
rect 12348 19182 12350 19234
rect 12402 19182 12404 19234
rect 12348 19170 12404 19182
rect 12460 18900 12516 24668
rect 12572 24724 12628 24734
rect 12572 24630 12628 24668
rect 12796 21588 12852 21598
rect 12908 21588 12964 26852
rect 13020 26180 13076 26190
rect 13020 26086 13076 26124
rect 13132 23548 13188 27356
rect 12852 21532 12964 21588
rect 13020 23492 13188 23548
rect 12796 21494 12852 21532
rect 12908 21140 12964 21150
rect 12908 20914 12964 21084
rect 12908 20862 12910 20914
rect 12962 20862 12964 20914
rect 12908 20850 12964 20862
rect 12572 20804 12628 20814
rect 12572 20018 12628 20748
rect 12572 19966 12574 20018
rect 12626 19966 12628 20018
rect 12572 19954 12628 19966
rect 12684 19460 12740 19470
rect 12684 19122 12740 19404
rect 12684 19070 12686 19122
rect 12738 19070 12740 19122
rect 12684 19058 12740 19070
rect 12460 18834 12516 18844
rect 13020 18674 13076 23492
rect 13244 20356 13300 30940
rect 13356 20804 13412 33740
rect 13468 28868 13524 35756
rect 13580 35140 13636 35150
rect 13580 35026 13636 35084
rect 13580 34974 13582 35026
rect 13634 34974 13636 35026
rect 13580 34962 13636 34974
rect 13580 32676 13636 32686
rect 13580 32450 13636 32620
rect 13580 32398 13582 32450
rect 13634 32398 13636 32450
rect 13580 32386 13636 32398
rect 13468 28812 13636 28868
rect 13468 28644 13524 28654
rect 13468 28550 13524 28588
rect 13468 27412 13524 27422
rect 13468 24948 13524 27356
rect 13580 27076 13636 28812
rect 13580 27010 13636 27020
rect 13692 26908 13748 40908
rect 13916 40626 13972 41916
rect 14364 41186 14420 41916
rect 15036 41300 15092 44200
rect 15036 41298 15316 41300
rect 15036 41246 15038 41298
rect 15090 41246 15316 41298
rect 15036 41244 15316 41246
rect 15036 41234 15092 41244
rect 14364 41134 14366 41186
rect 14418 41134 14420 41186
rect 14364 41122 14420 41134
rect 15260 41186 15316 41244
rect 15260 41134 15262 41186
rect 15314 41134 15316 41186
rect 15260 41122 15316 41134
rect 16156 41188 16212 44200
rect 17276 41300 17332 44200
rect 18396 41300 18452 44200
rect 19516 41300 19572 44200
rect 17276 41298 17780 41300
rect 17276 41246 17278 41298
rect 17330 41246 17780 41298
rect 17276 41244 17780 41246
rect 17276 41234 17332 41244
rect 16156 41186 16660 41188
rect 16156 41134 16158 41186
rect 16210 41134 16660 41186
rect 16156 41132 16660 41134
rect 16156 41122 16212 41132
rect 13916 40574 13918 40626
rect 13970 40574 13972 40626
rect 13916 40562 13972 40574
rect 14140 40962 14196 40974
rect 14140 40910 14142 40962
rect 14194 40910 14196 40962
rect 14140 38500 14196 40910
rect 15596 40962 15652 40974
rect 15596 40910 15598 40962
rect 15650 40910 15652 40962
rect 15372 40290 15428 40302
rect 15372 40238 15374 40290
rect 15426 40238 15428 40290
rect 14924 39396 14980 39406
rect 14812 38836 14868 38846
rect 14252 38724 14308 38734
rect 14252 38722 14532 38724
rect 14252 38670 14254 38722
rect 14306 38670 14532 38722
rect 14252 38668 14532 38670
rect 14252 38658 14308 38668
rect 14140 38434 14196 38444
rect 13916 38276 13972 38286
rect 13916 38274 14196 38276
rect 13916 38222 13918 38274
rect 13970 38222 14196 38274
rect 13916 38220 14196 38222
rect 13916 38210 13972 38220
rect 14028 38052 14084 38062
rect 14140 38052 14196 38220
rect 14476 38162 14532 38668
rect 14476 38110 14478 38162
rect 14530 38110 14532 38162
rect 14476 38098 14532 38110
rect 14252 38052 14308 38062
rect 14140 38050 14308 38052
rect 14140 37998 14254 38050
rect 14306 37998 14308 38050
rect 14140 37996 14308 37998
rect 14028 37958 14084 37996
rect 14252 37986 14308 37996
rect 14812 38050 14868 38780
rect 14924 38834 14980 39340
rect 15372 39396 15428 40238
rect 15596 39844 15652 40910
rect 16380 40962 16436 40974
rect 16380 40910 16382 40962
rect 16434 40910 16436 40962
rect 15652 39788 15876 39844
rect 15596 39778 15652 39788
rect 15596 39508 15652 39518
rect 15596 39506 15764 39508
rect 15596 39454 15598 39506
rect 15650 39454 15764 39506
rect 15596 39452 15764 39454
rect 15596 39442 15652 39452
rect 15372 39330 15428 39340
rect 15708 39058 15764 39452
rect 15708 39006 15710 39058
rect 15762 39006 15764 39058
rect 15708 38994 15764 39006
rect 14924 38782 14926 38834
rect 14978 38782 14980 38834
rect 14924 38770 14980 38782
rect 15484 38836 15540 38846
rect 15484 38742 15540 38780
rect 15596 38834 15652 38846
rect 15596 38782 15598 38834
rect 15650 38782 15652 38834
rect 14812 37998 14814 38050
rect 14866 37998 14868 38050
rect 14812 37986 14868 37998
rect 15260 38050 15316 38062
rect 15260 37998 15262 38050
rect 15314 37998 15316 38050
rect 14700 37938 14756 37950
rect 14700 37886 14702 37938
rect 14754 37886 14756 37938
rect 13916 37828 13972 37838
rect 13916 37734 13972 37772
rect 14140 37716 14196 37726
rect 13916 37266 13972 37278
rect 13916 37214 13918 37266
rect 13970 37214 13972 37266
rect 13916 36596 13972 37214
rect 13916 36530 13972 36540
rect 13916 36372 13972 36382
rect 13916 35698 13972 36316
rect 13916 35646 13918 35698
rect 13970 35646 13972 35698
rect 13916 35634 13972 35646
rect 13804 33122 13860 33134
rect 13804 33070 13806 33122
rect 13858 33070 13860 33122
rect 13804 32002 13860 33070
rect 14028 33122 14084 33134
rect 14028 33070 14030 33122
rect 14082 33070 14084 33122
rect 13804 31950 13806 32002
rect 13858 31950 13860 32002
rect 13804 31938 13860 31950
rect 13916 32562 13972 32574
rect 13916 32510 13918 32562
rect 13970 32510 13972 32562
rect 13916 32004 13972 32510
rect 14028 32452 14084 33070
rect 14028 32386 14084 32396
rect 14140 32004 14196 37660
rect 14364 37492 14420 37502
rect 14364 37266 14420 37436
rect 14364 37214 14366 37266
rect 14418 37214 14420 37266
rect 14364 37202 14420 37214
rect 14588 37378 14644 37390
rect 14588 37326 14590 37378
rect 14642 37326 14644 37378
rect 14588 35812 14644 37326
rect 14700 36708 14756 37886
rect 15260 37716 15316 37998
rect 15484 38052 15540 38062
rect 15484 37958 15540 37996
rect 15260 37650 15316 37660
rect 15148 37604 15204 37614
rect 15148 37492 15204 37548
rect 15260 37492 15316 37502
rect 15148 37490 15316 37492
rect 15148 37438 15262 37490
rect 15314 37438 15316 37490
rect 15148 37436 15316 37438
rect 15260 37426 15316 37436
rect 15484 37492 15540 37502
rect 15596 37492 15652 38782
rect 15820 38668 15876 39788
rect 16156 39732 16212 39742
rect 16156 38948 16212 39676
rect 16268 39618 16324 39630
rect 16268 39566 16270 39618
rect 16322 39566 16324 39618
rect 16268 39396 16324 39566
rect 16268 39330 16324 39340
rect 15484 37490 15652 37492
rect 15484 37438 15486 37490
rect 15538 37438 15652 37490
rect 15484 37436 15652 37438
rect 15708 38612 15876 38668
rect 16044 38834 16100 38846
rect 16044 38782 16046 38834
rect 16098 38782 16100 38834
rect 15484 37426 15540 37436
rect 15148 37268 15204 37278
rect 15148 37266 15540 37268
rect 15148 37214 15150 37266
rect 15202 37214 15540 37266
rect 15148 37212 15540 37214
rect 15148 37202 15204 37212
rect 15372 37044 15428 37054
rect 14700 36642 14756 36652
rect 15148 36988 15372 37044
rect 14924 36596 14980 36606
rect 14924 36502 14980 36540
rect 14476 35810 14644 35812
rect 14476 35758 14590 35810
rect 14642 35758 14644 35810
rect 14476 35756 14644 35758
rect 14364 35700 14420 35710
rect 14364 35606 14420 35644
rect 14252 33236 14308 33246
rect 14476 33236 14532 35756
rect 14588 35746 14644 35756
rect 14924 34914 14980 34926
rect 14924 34862 14926 34914
rect 14978 34862 14980 34914
rect 14588 34804 14644 34814
rect 14924 34804 14980 34862
rect 14588 34802 14980 34804
rect 14588 34750 14590 34802
rect 14642 34750 14980 34802
rect 14588 34748 14980 34750
rect 14588 34738 14644 34748
rect 14924 34468 14980 34748
rect 15036 34468 15092 34478
rect 14924 34412 15036 34468
rect 15036 34402 15092 34412
rect 14252 33234 14532 33236
rect 14252 33182 14254 33234
rect 14306 33182 14532 33234
rect 14252 33180 14532 33182
rect 14588 33684 14644 33694
rect 14252 33170 14308 33180
rect 14364 32676 14420 33180
rect 14588 32786 14644 33628
rect 14700 33460 14756 33470
rect 14700 33346 14756 33404
rect 14700 33294 14702 33346
rect 14754 33294 14756 33346
rect 14700 33282 14756 33294
rect 14588 32734 14590 32786
rect 14642 32734 14644 32786
rect 14588 32722 14644 32734
rect 14364 32582 14420 32620
rect 14924 32564 14980 32574
rect 14924 32470 14980 32508
rect 15148 32562 15204 36988
rect 15372 36978 15428 36988
rect 15484 36932 15540 37212
rect 15372 36708 15428 36718
rect 15372 36614 15428 36652
rect 15484 36482 15540 36876
rect 15484 36430 15486 36482
rect 15538 36430 15540 36482
rect 15484 36418 15540 36430
rect 15372 36260 15428 36270
rect 15372 36166 15428 36204
rect 15260 35700 15316 35710
rect 15260 35606 15316 35644
rect 15708 35028 15764 38612
rect 15820 38276 15876 38286
rect 15820 38182 15876 38220
rect 16044 38050 16100 38782
rect 16044 37998 16046 38050
rect 16098 37998 16100 38050
rect 16044 37986 16100 37998
rect 16156 37940 16212 38892
rect 16380 39060 16436 40910
rect 16604 40626 16660 41132
rect 17724 41186 17780 41244
rect 18396 41298 18900 41300
rect 18396 41246 18398 41298
rect 18450 41246 18900 41298
rect 18396 41244 18900 41246
rect 18396 41234 18452 41244
rect 17724 41134 17726 41186
rect 17778 41134 17780 41186
rect 17724 41122 17780 41134
rect 18844 41186 18900 41244
rect 19516 41298 20020 41300
rect 19516 41246 19518 41298
rect 19570 41246 20020 41298
rect 19516 41244 20020 41246
rect 19516 41234 19572 41244
rect 18844 41134 18846 41186
rect 18898 41134 18900 41186
rect 18844 41122 18900 41134
rect 19964 41186 20020 41244
rect 19964 41134 19966 41186
rect 20018 41134 20020 41186
rect 19964 41122 20020 41134
rect 20636 41188 20692 44200
rect 21756 41412 21812 44200
rect 22428 41412 22484 41422
rect 21756 41410 22484 41412
rect 21756 41358 22430 41410
rect 22482 41358 22484 41410
rect 21756 41356 22484 41358
rect 22428 41346 22484 41356
rect 20972 41188 21028 41198
rect 20636 41186 21364 41188
rect 20636 41134 20974 41186
rect 21026 41134 21364 41186
rect 20636 41132 21364 41134
rect 20972 41122 21028 41132
rect 17500 40964 17556 40974
rect 16604 40574 16606 40626
rect 16658 40574 16660 40626
rect 16604 40562 16660 40574
rect 17052 40962 17556 40964
rect 17052 40910 17502 40962
rect 17554 40910 17556 40962
rect 17052 40908 17556 40910
rect 16268 38722 16324 38734
rect 16268 38670 16270 38722
rect 16322 38670 16324 38722
rect 16268 38388 16324 38670
rect 16380 38668 16436 39004
rect 16828 39508 16884 39518
rect 16828 39058 16884 39452
rect 16828 39006 16830 39058
rect 16882 39006 16884 39058
rect 16828 38994 16884 39006
rect 16940 39396 16996 39406
rect 16492 38948 16548 38958
rect 16492 38834 16548 38892
rect 16492 38782 16494 38834
rect 16546 38782 16548 38834
rect 16492 38770 16548 38782
rect 16380 38612 16772 38668
rect 16268 38322 16324 38332
rect 16380 38164 16436 38174
rect 16380 38052 16436 38108
rect 16380 38050 16548 38052
rect 16380 37998 16382 38050
rect 16434 37998 16548 38050
rect 16380 37996 16548 37998
rect 16380 37986 16436 37996
rect 16268 37940 16324 37950
rect 16156 37938 16324 37940
rect 16156 37886 16270 37938
rect 16322 37886 16324 37938
rect 16156 37884 16324 37886
rect 16268 37874 16324 37884
rect 16268 37604 16324 37614
rect 15932 37492 15988 37502
rect 15932 37398 15988 37436
rect 16268 37490 16324 37548
rect 16268 37438 16270 37490
rect 16322 37438 16324 37490
rect 16268 37426 16324 37438
rect 15820 36484 15876 36494
rect 15820 35138 15876 36428
rect 16492 36370 16548 37996
rect 16492 36318 16494 36370
rect 16546 36318 16548 36370
rect 16492 36306 16548 36318
rect 16044 36260 16100 36270
rect 16044 36166 16100 36204
rect 15820 35086 15822 35138
rect 15874 35086 15876 35138
rect 15820 35074 15876 35086
rect 16268 35586 16324 35598
rect 16268 35534 16270 35586
rect 16322 35534 16324 35586
rect 15596 34972 15764 35028
rect 15372 34914 15428 34926
rect 15372 34862 15374 34914
rect 15426 34862 15428 34914
rect 15372 34692 15428 34862
rect 15372 34626 15428 34636
rect 15484 34804 15540 34814
rect 15260 34580 15316 34590
rect 15260 33346 15316 34524
rect 15260 33294 15262 33346
rect 15314 33294 15316 33346
rect 15260 33282 15316 33294
rect 15484 33124 15540 34748
rect 15596 33572 15652 34972
rect 15708 34804 15764 34814
rect 15708 34710 15764 34748
rect 16268 34804 16324 35534
rect 16268 34738 16324 34748
rect 15820 34692 15876 34702
rect 16492 34692 16548 34702
rect 15596 33506 15652 33516
rect 15708 34468 15764 34478
rect 15708 33684 15764 34412
rect 15148 32510 15150 32562
rect 15202 32510 15204 32562
rect 15148 32498 15204 32510
rect 15260 33068 15540 33124
rect 15708 33346 15764 33628
rect 15708 33294 15710 33346
rect 15762 33294 15764 33346
rect 14140 31948 14420 32004
rect 13916 31938 13972 31948
rect 14140 31780 14196 31790
rect 14028 31556 14084 31566
rect 13916 31500 14028 31556
rect 13804 31220 13860 31230
rect 13916 31220 13972 31500
rect 14028 31462 14084 31500
rect 14140 31220 14196 31724
rect 13860 31164 13972 31220
rect 14028 31164 14196 31220
rect 13804 31154 13860 31164
rect 14028 30772 14084 31164
rect 14140 30996 14196 31006
rect 14196 30940 14308 30996
rect 14140 30902 14196 30940
rect 14028 30716 14196 30772
rect 13916 29652 13972 29662
rect 13916 28642 13972 29596
rect 13916 28590 13918 28642
rect 13970 28590 13972 28642
rect 13916 28578 13972 28590
rect 14140 28642 14196 30716
rect 14140 28590 14142 28642
rect 14194 28590 14196 28642
rect 14140 28578 14196 28590
rect 13468 24854 13524 24892
rect 13580 26852 13748 26908
rect 14028 28530 14084 28542
rect 14028 28478 14030 28530
rect 14082 28478 14084 28530
rect 13580 26180 13636 26852
rect 13468 24724 13524 24734
rect 13468 24388 13524 24668
rect 13468 24322 13524 24332
rect 13580 24052 13636 26124
rect 13580 23986 13636 23996
rect 13692 25620 13748 25630
rect 13468 21474 13524 21486
rect 13468 21422 13470 21474
rect 13522 21422 13524 21474
rect 13468 20916 13524 21422
rect 13468 20850 13524 20860
rect 13580 21140 13636 21150
rect 13356 20692 13412 20748
rect 13468 20692 13524 20702
rect 13356 20690 13524 20692
rect 13356 20638 13470 20690
rect 13522 20638 13524 20690
rect 13356 20636 13524 20638
rect 13468 20626 13524 20636
rect 13580 20690 13636 21084
rect 13580 20638 13582 20690
rect 13634 20638 13636 20690
rect 13580 20626 13636 20638
rect 13244 20300 13524 20356
rect 13244 20130 13300 20142
rect 13244 20078 13246 20130
rect 13298 20078 13300 20130
rect 13132 20020 13188 20030
rect 13132 19926 13188 19964
rect 13244 19460 13300 20078
rect 13244 19394 13300 19404
rect 13356 20132 13412 20142
rect 13020 18622 13022 18674
rect 13074 18622 13076 18674
rect 13020 18610 13076 18622
rect 13244 18788 13300 18798
rect 11788 17042 11844 17052
rect 12348 18450 12404 18462
rect 12348 18398 12350 18450
rect 12402 18398 12404 18450
rect 11900 16210 11956 16222
rect 11900 16158 11902 16210
rect 11954 16158 11956 16210
rect 11900 16100 11956 16158
rect 11508 15932 11844 15988
rect 11452 15894 11508 15932
rect 11452 15540 11508 15550
rect 11228 15538 11508 15540
rect 11228 15486 11454 15538
rect 11506 15486 11508 15538
rect 11228 15484 11508 15486
rect 11116 15474 11172 15484
rect 11452 15474 11508 15484
rect 11676 15540 11732 15550
rect 11676 15446 11732 15484
rect 11228 15314 11284 15326
rect 11228 15262 11230 15314
rect 11282 15262 11284 15314
rect 9548 13346 9604 13356
rect 9772 15036 9940 15092
rect 9996 15202 10052 15214
rect 9996 15150 9998 15202
rect 10050 15150 10052 15202
rect 8876 12290 8932 12302
rect 8876 12238 8878 12290
rect 8930 12238 8932 12290
rect 8764 12178 8820 12190
rect 8764 12126 8766 12178
rect 8818 12126 8820 12178
rect 7532 11396 7588 11406
rect 7532 11302 7588 11340
rect 7308 10670 7310 10722
rect 7362 10670 7364 10722
rect 7308 10658 7364 10670
rect 7756 10948 7812 10958
rect 7756 10834 7812 10892
rect 7756 10782 7758 10834
rect 7810 10782 7812 10834
rect 6748 10610 6916 10612
rect 6748 10558 6750 10610
rect 6802 10558 6916 10610
rect 6748 10556 6916 10558
rect 6972 10612 7028 10622
rect 6748 9940 6804 10556
rect 6972 10518 7028 10556
rect 6972 9940 7028 9950
rect 6748 9884 6972 9940
rect 6972 9846 7028 9884
rect 7420 9940 7476 9950
rect 7420 9846 7476 9884
rect 7756 9828 7812 10782
rect 8092 9940 8148 11676
rect 8316 12068 8372 12078
rect 8316 11506 8372 12012
rect 8316 11454 8318 11506
rect 8370 11454 8372 11506
rect 8316 11442 8372 11454
rect 8764 11284 8820 12126
rect 8876 11956 8932 12238
rect 9100 12180 9156 12190
rect 9436 12180 9492 12190
rect 9100 12178 9492 12180
rect 9100 12126 9102 12178
rect 9154 12126 9438 12178
rect 9490 12126 9492 12178
rect 9100 12124 9492 12126
rect 9100 12114 9156 12124
rect 9436 12114 9492 12124
rect 9660 12068 9716 12078
rect 9660 11974 9716 12012
rect 8876 11890 8932 11900
rect 8764 10724 8820 11228
rect 8764 10658 8820 10668
rect 8092 9874 8148 9884
rect 9548 9940 9604 9950
rect 7756 9762 7812 9772
rect 9548 9042 9604 9884
rect 9548 8990 9550 9042
rect 9602 8990 9604 9042
rect 9548 8978 9604 8990
rect 9772 8428 9828 15036
rect 9996 14756 10052 15150
rect 10220 15092 10276 15102
rect 10220 14998 10276 15036
rect 11116 15092 11172 15102
rect 9996 14690 10052 14700
rect 10892 14644 10948 14654
rect 10444 14530 10500 14542
rect 10444 14478 10446 14530
rect 10498 14478 10500 14530
rect 9996 14308 10052 14318
rect 9996 13972 10052 14252
rect 9996 13906 10052 13916
rect 10444 13972 10500 14478
rect 10444 13906 10500 13916
rect 10780 13522 10836 13534
rect 10780 13470 10782 13522
rect 10834 13470 10836 13522
rect 10332 12740 10388 12750
rect 10332 12738 10500 12740
rect 10332 12686 10334 12738
rect 10386 12686 10500 12738
rect 10332 12684 10500 12686
rect 10332 12674 10388 12684
rect 10332 12404 10388 12414
rect 9884 12402 10388 12404
rect 9884 12350 10334 12402
rect 10386 12350 10388 12402
rect 9884 12348 10388 12350
rect 9884 12290 9940 12348
rect 10332 12338 10388 12348
rect 9884 12238 9886 12290
rect 9938 12238 9940 12290
rect 9884 12226 9940 12238
rect 10108 12180 10164 12190
rect 10444 12180 10500 12684
rect 10556 12404 10612 12414
rect 10556 12310 10612 12348
rect 10108 12178 10500 12180
rect 10108 12126 10110 12178
rect 10162 12126 10500 12178
rect 10108 12124 10500 12126
rect 10668 12178 10724 12190
rect 10668 12126 10670 12178
rect 10722 12126 10724 12178
rect 10108 11732 10164 12124
rect 10108 11666 10164 11676
rect 10444 11956 10500 11966
rect 10444 11506 10500 11900
rect 10668 11844 10724 12126
rect 10668 11778 10724 11788
rect 10780 11620 10836 13470
rect 10892 13524 10948 14588
rect 11004 14084 11060 14094
rect 11004 13746 11060 14028
rect 11004 13694 11006 13746
rect 11058 13694 11060 13746
rect 11004 13682 11060 13694
rect 10892 13468 11060 13524
rect 10892 13076 10948 13086
rect 10892 11956 10948 13020
rect 10892 11890 10948 11900
rect 10444 11454 10446 11506
rect 10498 11454 10500 11506
rect 10444 11442 10500 11454
rect 10556 11564 10836 11620
rect 9996 10836 10052 10846
rect 9996 9604 10052 10780
rect 9996 9538 10052 9548
rect 10556 9380 10612 11564
rect 10668 11396 10724 11406
rect 10668 10836 10724 11340
rect 10892 11284 10948 11294
rect 10892 11190 10948 11228
rect 11004 11172 11060 13468
rect 11004 11106 11060 11116
rect 11116 10948 11172 15036
rect 11228 13634 11284 15262
rect 11340 15316 11396 15326
rect 11340 15222 11396 15260
rect 11564 15314 11620 15326
rect 11564 15262 11566 15314
rect 11618 15262 11620 15314
rect 11564 15148 11620 15262
rect 11788 15204 11844 15932
rect 11900 15316 11956 16044
rect 11900 15250 11956 15260
rect 11564 15092 11732 15148
rect 11564 14308 11620 14318
rect 11228 13582 11230 13634
rect 11282 13582 11284 13634
rect 11228 13076 11284 13582
rect 11228 13010 11284 13020
rect 11340 14306 11620 14308
rect 11340 14254 11566 14306
rect 11618 14254 11620 14306
rect 11340 14252 11620 14254
rect 11228 12404 11284 12414
rect 11228 12310 11284 12348
rect 11228 11396 11284 11406
rect 11340 11396 11396 14252
rect 11564 14242 11620 14252
rect 11676 12292 11732 15092
rect 11788 14418 11844 15148
rect 12124 15092 12180 15102
rect 12012 15090 12180 15092
rect 12012 15038 12126 15090
rect 12178 15038 12180 15090
rect 12012 15036 12180 15038
rect 11788 14366 11790 14418
rect 11842 14366 11844 14418
rect 11788 14354 11844 14366
rect 11900 14418 11956 14430
rect 11900 14366 11902 14418
rect 11954 14366 11956 14418
rect 11900 14308 11956 14366
rect 11900 14242 11956 14252
rect 11900 14084 11956 14094
rect 11900 13970 11956 14028
rect 11900 13918 11902 13970
rect 11954 13918 11956 13970
rect 11900 13906 11956 13918
rect 11676 12226 11732 12236
rect 12012 11956 12068 15036
rect 12124 15026 12180 15036
rect 12348 14532 12404 18398
rect 12908 18450 12964 18462
rect 12908 18398 12910 18450
rect 12962 18398 12964 18450
rect 12572 16212 12628 16222
rect 12460 15764 12516 15774
rect 12460 15314 12516 15708
rect 12460 15262 12462 15314
rect 12514 15262 12516 15314
rect 12460 15250 12516 15262
rect 12460 14532 12516 14542
rect 12348 14476 12460 14532
rect 12460 14466 12516 14476
rect 12348 14308 12404 14318
rect 12572 14308 12628 16156
rect 12908 16100 12964 18398
rect 13020 16882 13076 16894
rect 13020 16830 13022 16882
rect 13074 16830 13076 16882
rect 13020 16660 13076 16830
rect 13020 16594 13076 16604
rect 12908 16034 12964 16044
rect 13132 15764 13188 15774
rect 13132 15538 13188 15708
rect 13132 15486 13134 15538
rect 13186 15486 13188 15538
rect 13132 15474 13188 15486
rect 12684 15204 12740 15242
rect 12684 15138 12740 15148
rect 12404 14252 12628 14308
rect 12348 14214 12404 14252
rect 11676 11900 12068 11956
rect 13132 12740 13188 12750
rect 11676 11396 11732 11900
rect 12908 11844 12964 11854
rect 11228 11394 11396 11396
rect 11228 11342 11230 11394
rect 11282 11342 11396 11394
rect 11228 11340 11396 11342
rect 11228 11330 11284 11340
rect 11116 10892 11284 10948
rect 10668 10834 11172 10836
rect 10668 10782 10670 10834
rect 10722 10782 11172 10834
rect 10668 10780 11172 10782
rect 10668 10770 10724 10780
rect 11116 10610 11172 10780
rect 11116 10558 11118 10610
rect 11170 10558 11172 10610
rect 11116 10546 11172 10558
rect 11116 9604 11172 9614
rect 10444 9324 10612 9380
rect 10668 9602 11172 9604
rect 10668 9550 11118 9602
rect 11170 9550 11172 9602
rect 10668 9548 11172 9550
rect 9996 9044 10052 9054
rect 10332 9044 10388 9054
rect 9436 8372 9828 8428
rect 9884 9042 10052 9044
rect 9884 8990 9998 9042
rect 10050 8990 10052 9042
rect 9884 8988 10052 8990
rect 9884 8372 9940 8988
rect 9996 8978 10052 8988
rect 10220 9042 10388 9044
rect 10220 8990 10334 9042
rect 10386 8990 10388 9042
rect 10220 8988 10388 8990
rect 10220 8596 10276 8988
rect 10332 8978 10388 8988
rect 9436 8148 9492 8372
rect 9884 8306 9940 8316
rect 9996 8540 10276 8596
rect 9996 8258 10052 8540
rect 10444 8428 10500 9324
rect 10556 9154 10612 9166
rect 10556 9102 10558 9154
rect 10610 9102 10612 9154
rect 10556 8820 10612 9102
rect 10668 9156 10724 9548
rect 11116 9538 11172 9548
rect 11228 9380 11284 10892
rect 11116 9324 11284 9380
rect 10668 9154 10836 9156
rect 10668 9102 10670 9154
rect 10722 9102 10836 9154
rect 10668 9100 10836 9102
rect 10668 9090 10724 9100
rect 10556 8754 10612 8764
rect 9996 8206 9998 8258
rect 10050 8206 10052 8258
rect 9996 8194 10052 8206
rect 10108 8372 10500 8428
rect 10668 8372 10724 8382
rect 9436 8082 9492 8092
rect 9772 8146 9828 8158
rect 9772 8094 9774 8146
rect 9826 8094 9828 8146
rect 7868 8036 7924 8046
rect 7084 6692 7140 6702
rect 6636 6636 7084 6692
rect 7084 6598 7140 6636
rect 7868 6690 7924 7980
rect 9772 7700 9828 8094
rect 9884 8036 9940 8046
rect 9884 7942 9940 7980
rect 9772 7634 9828 7644
rect 9996 7476 10052 7486
rect 9996 6802 10052 7420
rect 9996 6750 9998 6802
rect 10050 6750 10052 6802
rect 9996 6738 10052 6750
rect 7868 6638 7870 6690
rect 7922 6638 7924 6690
rect 7868 6626 7924 6638
rect 8092 6692 8148 6702
rect 8092 5122 8148 6636
rect 8876 6468 8932 6478
rect 8876 5234 8932 6412
rect 8876 5182 8878 5234
rect 8930 5182 8932 5234
rect 8876 5170 8932 5182
rect 8092 5070 8094 5122
rect 8146 5070 8148 5122
rect 8092 5058 8148 5070
rect 10108 4564 10164 8372
rect 10332 8146 10388 8158
rect 10332 8094 10334 8146
rect 10386 8094 10388 8146
rect 10332 8036 10388 8094
rect 10220 7700 10276 7710
rect 10220 7606 10276 7644
rect 10220 6692 10276 6702
rect 10220 6130 10276 6636
rect 10332 6690 10388 7980
rect 10668 8146 10724 8316
rect 10780 8260 10836 9100
rect 11116 8708 11172 9324
rect 11116 8642 11172 8652
rect 11228 9154 11284 9166
rect 11228 9102 11230 9154
rect 11282 9102 11284 9154
rect 11228 8428 11284 9102
rect 11340 9044 11396 11340
rect 11452 11394 11732 11396
rect 11452 11342 11678 11394
rect 11730 11342 11732 11394
rect 11452 11340 11732 11342
rect 11452 9826 11508 11340
rect 11676 11330 11732 11340
rect 11900 11732 11956 11742
rect 11900 11282 11956 11676
rect 11900 11230 11902 11282
rect 11954 11230 11956 11282
rect 11900 11218 11956 11230
rect 12012 11284 12068 11294
rect 12236 11284 12292 11294
rect 12068 11282 12292 11284
rect 12068 11230 12238 11282
rect 12290 11230 12292 11282
rect 12068 11228 12292 11230
rect 12012 11218 12068 11228
rect 12236 11218 12292 11228
rect 12348 11284 12404 11294
rect 12348 11190 12404 11228
rect 11452 9774 11454 9826
rect 11506 9774 11508 9826
rect 11452 9762 11508 9774
rect 11564 11172 11620 11182
rect 12572 11172 12628 11182
rect 11452 9044 11508 9054
rect 11340 9042 11508 9044
rect 11340 8990 11454 9042
rect 11506 8990 11508 9042
rect 11340 8988 11508 8990
rect 11452 8978 11508 8988
rect 11564 8428 11620 11116
rect 12460 11170 12628 11172
rect 12460 11118 12574 11170
rect 12626 11118 12628 11170
rect 12460 11116 12628 11118
rect 11900 10500 11956 10510
rect 11900 10498 12292 10500
rect 11900 10446 11902 10498
rect 11954 10446 12292 10498
rect 11900 10444 12292 10446
rect 11900 10434 11956 10444
rect 12236 9938 12292 10444
rect 12236 9886 12238 9938
rect 12290 9886 12292 9938
rect 12236 9874 12292 9886
rect 12124 9826 12180 9838
rect 12124 9774 12126 9826
rect 12178 9774 12180 9826
rect 11788 9716 11844 9726
rect 11788 9714 11956 9716
rect 11788 9662 11790 9714
rect 11842 9662 11956 9714
rect 11788 9660 11956 9662
rect 11788 9650 11844 9660
rect 10780 8194 10836 8204
rect 10892 8372 11396 8428
rect 10668 8094 10670 8146
rect 10722 8094 10724 8146
rect 10668 7924 10724 8094
rect 10780 7924 10836 7934
rect 10668 7868 10780 7924
rect 10780 7858 10836 7868
rect 10444 7700 10500 7710
rect 10892 7700 10948 8372
rect 11004 8036 11060 8046
rect 11228 8036 11284 8046
rect 11004 7942 11060 7980
rect 11116 8034 11284 8036
rect 11116 7982 11230 8034
rect 11282 7982 11284 8034
rect 11116 7980 11284 7982
rect 10444 7606 10500 7644
rect 10556 7644 10948 7700
rect 10556 7586 10612 7644
rect 10556 7534 10558 7586
rect 10610 7534 10612 7586
rect 10556 7522 10612 7534
rect 11004 7364 11060 7374
rect 11004 7270 11060 7308
rect 11116 7140 11172 7980
rect 11228 7970 11284 7980
rect 10332 6638 10334 6690
rect 10386 6638 10388 6690
rect 10332 6626 10388 6638
rect 10668 7084 11172 7140
rect 10668 6690 10724 7084
rect 10668 6638 10670 6690
rect 10722 6638 10724 6690
rect 10668 6626 10724 6638
rect 11340 6692 11396 8372
rect 11452 8372 11620 8428
rect 11788 9492 11844 9502
rect 11452 8034 11508 8372
rect 11564 8260 11620 8270
rect 11564 8166 11620 8204
rect 11452 7982 11454 8034
rect 11506 7982 11508 8034
rect 11452 7252 11508 7982
rect 11788 7700 11844 9436
rect 11900 8428 11956 9660
rect 12124 9604 12180 9774
rect 12460 9826 12516 11116
rect 12572 11106 12628 11116
rect 12796 10052 12852 10062
rect 12460 9774 12462 9826
rect 12514 9774 12516 9826
rect 12460 9762 12516 9774
rect 12572 10050 12852 10052
rect 12572 9998 12798 10050
rect 12850 9998 12852 10050
rect 12572 9996 12852 9998
rect 12572 9604 12628 9996
rect 12796 9986 12852 9996
rect 12684 9828 12740 9838
rect 12908 9828 12964 11788
rect 12684 9826 12964 9828
rect 12684 9774 12686 9826
rect 12738 9774 12964 9826
rect 12684 9772 12964 9774
rect 13020 9940 13076 9950
rect 12684 9762 12740 9772
rect 12124 9548 12628 9604
rect 12796 9604 12852 9614
rect 13020 9604 13076 9884
rect 12796 9602 13076 9604
rect 12796 9550 12798 9602
rect 12850 9550 13076 9602
rect 12796 9548 13076 9550
rect 12796 9538 12852 9548
rect 12012 8930 12068 8942
rect 12012 8878 12014 8930
rect 12066 8878 12068 8930
rect 12012 8820 12068 8878
rect 12012 8754 12068 8764
rect 11900 8372 12068 8428
rect 11788 7634 11844 7644
rect 12012 8036 12068 8372
rect 13020 8372 13076 8382
rect 12908 8260 12964 8270
rect 12908 8166 12964 8204
rect 12348 8148 12404 8158
rect 12348 8054 12404 8092
rect 12796 8148 12852 8158
rect 12796 8054 12852 8092
rect 12572 8036 12628 8046
rect 12012 7586 12068 7980
rect 12460 8034 12628 8036
rect 12460 7982 12574 8034
rect 12626 7982 12628 8034
rect 12460 7980 12628 7982
rect 12460 7588 12516 7980
rect 12572 7970 12628 7980
rect 12012 7534 12014 7586
rect 12066 7534 12068 7586
rect 12012 7522 12068 7534
rect 12348 7532 12516 7588
rect 12572 7644 12964 7700
rect 12348 7474 12404 7532
rect 12348 7422 12350 7474
rect 12402 7422 12404 7474
rect 12348 7410 12404 7422
rect 11452 7186 11508 7196
rect 11676 7364 11732 7374
rect 11452 6692 11508 6702
rect 11340 6636 11452 6692
rect 11452 6598 11508 6636
rect 10892 6580 10948 6590
rect 11116 6580 11172 6590
rect 10892 6578 11172 6580
rect 10892 6526 10894 6578
rect 10946 6526 11118 6578
rect 11170 6526 11172 6578
rect 10892 6524 11172 6526
rect 10892 6514 10948 6524
rect 11116 6514 11172 6524
rect 10668 6468 10724 6478
rect 11340 6468 11396 6478
rect 10668 6374 10724 6412
rect 11228 6412 11340 6468
rect 10220 6078 10222 6130
rect 10274 6078 10276 6130
rect 10220 5908 10276 6078
rect 10220 5842 10276 5852
rect 10556 5908 10612 5918
rect 10108 4498 10164 4508
rect 10220 5236 10276 5246
rect 6412 4286 6414 4338
rect 6466 4286 6468 4338
rect 6412 4274 6468 4286
rect 10108 4340 10164 4350
rect 10220 4340 10276 5180
rect 10556 4562 10612 5852
rect 10892 5908 10948 5918
rect 10892 5814 10948 5852
rect 11004 5236 11060 5246
rect 11228 5236 11284 6412
rect 11340 6374 11396 6412
rect 11676 6018 11732 7308
rect 12460 7364 12516 7374
rect 12460 7270 12516 7308
rect 11676 5966 11678 6018
rect 11730 5966 11732 6018
rect 11676 5954 11732 5966
rect 11900 6916 11956 6926
rect 11900 6690 11956 6860
rect 11900 6638 11902 6690
rect 11954 6638 11956 6690
rect 11900 6468 11956 6638
rect 12572 6692 12628 7644
rect 12908 7586 12964 7644
rect 13020 7698 13076 8316
rect 13020 7646 13022 7698
rect 13074 7646 13076 7698
rect 13020 7634 13076 7646
rect 12908 7534 12910 7586
rect 12962 7534 12964 7586
rect 12908 7522 12964 7534
rect 12684 7474 12740 7486
rect 12684 7422 12686 7474
rect 12738 7422 12740 7474
rect 12684 7252 12740 7422
rect 13020 7252 13076 7262
rect 12684 7250 13076 7252
rect 12684 7198 13022 7250
rect 13074 7198 13076 7250
rect 12684 7196 13076 7198
rect 13020 7186 13076 7196
rect 13132 6916 13188 12684
rect 12908 6860 13188 6916
rect 13244 6916 13300 18732
rect 13356 18562 13412 20076
rect 13356 18510 13358 18562
rect 13410 18510 13412 18562
rect 13356 16772 13412 18510
rect 13468 18452 13524 20300
rect 13692 19460 13748 25564
rect 13916 24836 13972 24846
rect 13916 24500 13972 24780
rect 13916 24434 13972 24444
rect 13804 20578 13860 20590
rect 13804 20526 13806 20578
rect 13858 20526 13860 20578
rect 13804 20244 13860 20526
rect 14028 20356 14084 28478
rect 14252 28420 14308 30940
rect 14364 30882 14420 31948
rect 14476 32002 14532 32014
rect 14476 31950 14478 32002
rect 14530 31950 14532 32002
rect 14476 31780 14532 31950
rect 14476 31554 14532 31724
rect 14476 31502 14478 31554
rect 14530 31502 14532 31554
rect 14476 31108 14532 31502
rect 14924 31556 14980 31566
rect 14924 31462 14980 31500
rect 14476 31042 14532 31052
rect 14364 30830 14366 30882
rect 14418 30830 14420 30882
rect 14364 29876 14420 30830
rect 15148 29988 15204 29998
rect 15260 29988 15316 33068
rect 15596 33012 15652 33022
rect 15484 32956 15596 33012
rect 15372 31780 15428 31790
rect 15372 31686 15428 31724
rect 15148 29986 15316 29988
rect 15148 29934 15150 29986
rect 15202 29934 15316 29986
rect 15148 29932 15316 29934
rect 15372 30884 15428 30894
rect 14364 29820 14644 29876
rect 14140 28364 14308 28420
rect 14140 27972 14196 28364
rect 14140 27916 14420 27972
rect 14140 26740 14196 26750
rect 14140 20692 14196 26684
rect 14252 21924 14308 21934
rect 14252 20914 14308 21868
rect 14364 21476 14420 27916
rect 14476 27524 14532 27534
rect 14476 26962 14532 27468
rect 14476 26910 14478 26962
rect 14530 26910 14532 26962
rect 14476 26898 14532 26910
rect 14476 26740 14532 26750
rect 14588 26740 14644 29820
rect 15148 29428 15204 29932
rect 15148 29362 15204 29372
rect 15372 29426 15428 30828
rect 15484 30210 15540 32956
rect 15596 32946 15652 32956
rect 15708 31780 15764 33294
rect 15820 32562 15876 34636
rect 16380 34690 16548 34692
rect 16380 34638 16494 34690
rect 16546 34638 16548 34690
rect 16380 34636 16548 34638
rect 16380 34132 16436 34636
rect 16492 34626 16548 34636
rect 15820 32510 15822 32562
rect 15874 32510 15876 32562
rect 15820 32498 15876 32510
rect 16268 33234 16324 33246
rect 16268 33182 16270 33234
rect 16322 33182 16324 33234
rect 16268 32674 16324 33182
rect 16268 32622 16270 32674
rect 16322 32622 16324 32674
rect 15708 31714 15764 31724
rect 15820 31778 15876 31790
rect 15820 31726 15822 31778
rect 15874 31726 15876 31778
rect 15484 30158 15486 30210
rect 15538 30158 15540 30210
rect 15484 30146 15540 30158
rect 15708 31444 15764 31454
rect 15708 30210 15764 31388
rect 15708 30158 15710 30210
rect 15762 30158 15764 30210
rect 15708 30146 15764 30158
rect 15820 30212 15876 31726
rect 16156 31556 16212 31566
rect 16268 31556 16324 32622
rect 16212 31500 16324 31556
rect 16156 31462 16212 31500
rect 16380 31332 16436 34076
rect 16492 33348 16548 33358
rect 16492 33254 16548 33292
rect 16716 32786 16772 38612
rect 16940 38162 16996 39340
rect 16940 38110 16942 38162
rect 16994 38110 16996 38162
rect 16940 38098 16996 38110
rect 16940 37828 16996 37838
rect 16828 36484 16884 36494
rect 16828 36390 16884 36428
rect 16940 36372 16996 37772
rect 16940 36306 16996 36316
rect 16940 34916 16996 34926
rect 16828 34860 16940 34916
rect 16828 33572 16884 34860
rect 16940 34822 16996 34860
rect 16828 33506 16884 33516
rect 16940 33458 16996 33470
rect 16940 33406 16942 33458
rect 16994 33406 16996 33458
rect 16940 33236 16996 33406
rect 16940 33170 16996 33180
rect 17052 33012 17108 40908
rect 17500 40898 17556 40908
rect 18620 40964 18676 40974
rect 19740 40964 19796 40974
rect 18620 40962 18900 40964
rect 18620 40910 18622 40962
rect 18674 40910 18900 40962
rect 18620 40908 18900 40910
rect 18620 40898 18676 40908
rect 17724 39618 17780 39630
rect 17724 39566 17726 39618
rect 17778 39566 17780 39618
rect 17388 39396 17444 39406
rect 17388 39302 17444 39340
rect 17724 39396 17780 39566
rect 18508 39508 18564 39518
rect 18284 39506 18564 39508
rect 18284 39454 18510 39506
rect 18562 39454 18564 39506
rect 18284 39452 18564 39454
rect 18172 39396 18228 39406
rect 17780 39340 17892 39396
rect 17724 39330 17780 39340
rect 17612 38722 17668 38734
rect 17612 38670 17614 38722
rect 17666 38670 17668 38722
rect 17164 38388 17220 38398
rect 17612 38388 17668 38670
rect 17220 38332 17668 38388
rect 17164 33460 17220 38332
rect 17276 38164 17332 38174
rect 17276 38050 17332 38108
rect 17276 37998 17278 38050
rect 17330 37998 17332 38050
rect 17276 37380 17332 37998
rect 17500 38164 17556 38174
rect 17388 37828 17444 37838
rect 17388 37734 17444 37772
rect 17500 37490 17556 38108
rect 17836 38050 17892 39340
rect 17836 37998 17838 38050
rect 17890 37998 17892 38050
rect 17836 37986 17892 37998
rect 18060 38834 18116 38846
rect 18060 38782 18062 38834
rect 18114 38782 18116 38834
rect 17612 37940 17668 37950
rect 17612 37846 17668 37884
rect 18060 37940 18116 38782
rect 18060 37874 18116 37884
rect 17500 37438 17502 37490
rect 17554 37438 17556 37490
rect 17388 37380 17444 37390
rect 17276 37378 17444 37380
rect 17276 37326 17390 37378
rect 17442 37326 17444 37378
rect 17276 37324 17444 37326
rect 17388 37314 17444 37324
rect 17500 37044 17556 37438
rect 18060 37380 18116 37390
rect 18060 37286 18116 37324
rect 17724 37268 17780 37278
rect 17724 37174 17780 37212
rect 17948 37266 18004 37278
rect 17948 37214 17950 37266
rect 18002 37214 18004 37266
rect 17500 36978 17556 36988
rect 17948 36932 18004 37214
rect 17948 36372 18004 36876
rect 18172 36596 18228 39340
rect 18284 39058 18340 39452
rect 18508 39442 18564 39452
rect 18284 39006 18286 39058
rect 18338 39006 18340 39058
rect 18284 38994 18340 39006
rect 18284 38834 18340 38846
rect 18284 38782 18286 38834
rect 18338 38782 18340 38834
rect 18284 37490 18340 38782
rect 18620 38836 18676 38846
rect 18620 38742 18676 38780
rect 18284 37438 18286 37490
rect 18338 37438 18340 37490
rect 18284 37426 18340 37438
rect 18620 37938 18676 37950
rect 18620 37886 18622 37938
rect 18674 37886 18676 37938
rect 18620 37490 18676 37886
rect 18620 37438 18622 37490
rect 18674 37438 18676 37490
rect 18620 37426 18676 37438
rect 18396 37268 18452 37278
rect 18732 37268 18788 37278
rect 18396 37174 18452 37212
rect 18508 37266 18788 37268
rect 18508 37214 18734 37266
rect 18786 37214 18788 37266
rect 18508 37212 18788 37214
rect 18508 37044 18564 37212
rect 18732 37202 18788 37212
rect 18284 36988 18564 37044
rect 18284 36706 18340 36988
rect 18284 36654 18286 36706
rect 18338 36654 18340 36706
rect 18284 36642 18340 36654
rect 17724 36316 17948 36372
rect 17724 35922 17780 36316
rect 17948 36306 18004 36316
rect 18060 36540 18228 36596
rect 17724 35870 17726 35922
rect 17778 35870 17780 35922
rect 17724 35858 17780 35870
rect 17948 35698 18004 35710
rect 17948 35646 17950 35698
rect 18002 35646 18004 35698
rect 17612 34804 17668 34814
rect 17388 34690 17444 34702
rect 17388 34638 17390 34690
rect 17442 34638 17444 34690
rect 17388 34130 17444 34638
rect 17388 34078 17390 34130
rect 17442 34078 17444 34130
rect 17388 33684 17444 34078
rect 17612 34692 17668 34748
rect 17948 34804 18004 35646
rect 17724 34692 17780 34702
rect 17612 34690 17780 34692
rect 17612 34638 17726 34690
rect 17778 34638 17780 34690
rect 17612 34636 17780 34638
rect 17612 34130 17668 34636
rect 17724 34626 17780 34636
rect 17948 34354 18004 34748
rect 17948 34302 17950 34354
rect 18002 34302 18004 34354
rect 17948 34290 18004 34302
rect 17612 34078 17614 34130
rect 17666 34078 17668 34130
rect 17612 34066 17668 34078
rect 17388 33618 17444 33628
rect 17164 33404 17668 33460
rect 17052 32946 17108 32956
rect 17500 33236 17556 33246
rect 16716 32734 16718 32786
rect 16770 32734 16772 32786
rect 16716 32722 16772 32734
rect 16940 32564 16996 32574
rect 16716 32452 16772 32462
rect 16156 31276 16436 31332
rect 16492 31554 16548 31566
rect 16492 31502 16494 31554
rect 16546 31502 16548 31554
rect 16492 31444 16548 31502
rect 16156 30884 16212 31276
rect 16156 30790 16212 30828
rect 16268 30772 16324 30782
rect 15820 30146 15876 30156
rect 15932 30436 15988 30446
rect 15932 30210 15988 30380
rect 16268 30322 16324 30716
rect 16268 30270 16270 30322
rect 16322 30270 16324 30322
rect 16268 30258 16324 30270
rect 15932 30158 15934 30210
rect 15986 30158 15988 30210
rect 15932 29652 15988 30158
rect 15372 29374 15374 29426
rect 15426 29374 15428 29426
rect 15148 28420 15204 28430
rect 15260 28420 15316 28430
rect 15148 28418 15260 28420
rect 15148 28366 15150 28418
rect 15202 28366 15260 28418
rect 15148 28364 15260 28366
rect 15148 28354 15204 28364
rect 15148 27860 15204 27870
rect 15148 27298 15204 27804
rect 15148 27246 15150 27298
rect 15202 27246 15204 27298
rect 15148 27234 15204 27246
rect 15260 27300 15316 28364
rect 15260 27234 15316 27244
rect 14812 27188 14868 27198
rect 14812 27074 14868 27132
rect 14812 27022 14814 27074
rect 14866 27022 14868 27074
rect 14812 27010 14868 27022
rect 14532 26684 14644 26740
rect 15372 26740 15428 29374
rect 15820 29596 15988 29652
rect 16156 30210 16212 30222
rect 16156 30158 16158 30210
rect 16210 30158 16212 30210
rect 15820 28644 15876 29596
rect 15820 28578 15876 28588
rect 15596 28420 15652 28430
rect 15596 28326 15652 28364
rect 15932 28420 15988 28430
rect 15932 28326 15988 28364
rect 16156 27860 16212 30158
rect 16380 30098 16436 30110
rect 16380 30046 16382 30098
rect 16434 30046 16436 30098
rect 16268 29988 16324 29998
rect 16268 28532 16324 29932
rect 16380 28756 16436 30046
rect 16380 28690 16436 28700
rect 16268 28466 16324 28476
rect 16268 28308 16324 28318
rect 16268 28082 16324 28252
rect 16268 28030 16270 28082
rect 16322 28030 16324 28082
rect 16268 28018 16324 28030
rect 16380 28196 16436 28206
rect 16380 27860 16436 28140
rect 16156 27804 16436 27860
rect 15596 27188 15652 27198
rect 14476 26674 14532 26684
rect 15372 26674 15428 26684
rect 15484 27132 15596 27188
rect 15484 26516 15540 27132
rect 15596 27122 15652 27132
rect 15708 27074 15764 27086
rect 15708 27022 15710 27074
rect 15762 27022 15764 27074
rect 15260 26514 15540 26516
rect 15260 26462 15486 26514
rect 15538 26462 15540 26514
rect 15260 26460 15540 26462
rect 15260 25620 15316 26460
rect 15484 26450 15540 26460
rect 15596 26962 15652 26974
rect 15596 26910 15598 26962
rect 15650 26910 15652 26962
rect 15596 26292 15652 26910
rect 15708 26964 15764 27022
rect 15932 27076 15988 27086
rect 16380 27076 16436 27804
rect 16492 27300 16548 31388
rect 16716 30210 16772 32396
rect 16940 31668 16996 32508
rect 17500 32562 17556 33180
rect 17500 32510 17502 32562
rect 17554 32510 17556 32562
rect 17500 32498 17556 32510
rect 17612 32452 17668 33404
rect 18060 32788 18116 36540
rect 18172 36372 18228 36382
rect 18172 36278 18228 36316
rect 18284 36260 18340 36270
rect 18284 36166 18340 36204
rect 18732 35028 18788 35038
rect 18732 34356 18788 34972
rect 18732 34262 18788 34300
rect 18844 33348 18900 40908
rect 19292 40962 19796 40964
rect 19292 40910 19742 40962
rect 19794 40910 19796 40962
rect 19292 40908 19796 40910
rect 19068 38836 19124 38846
rect 19068 37266 19124 38780
rect 19292 38668 19348 40908
rect 19740 40898 19796 40908
rect 20748 40962 20804 40974
rect 20748 40910 20750 40962
rect 20802 40910 20804 40962
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19628 40404 19684 40414
rect 19628 38946 19684 40348
rect 20748 40404 20804 40910
rect 21308 40626 21364 41132
rect 21308 40574 21310 40626
rect 21362 40574 21364 40626
rect 21308 40562 21364 40574
rect 21420 41186 21476 41198
rect 21420 41134 21422 41186
rect 21474 41134 21476 41186
rect 20748 40338 20804 40348
rect 21420 40068 21476 41134
rect 20412 40012 21476 40068
rect 22764 41188 22820 41198
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20412 39058 20468 40012
rect 20412 39006 20414 39058
rect 20466 39006 20468 39058
rect 20412 38994 20468 39006
rect 20636 39730 20692 39742
rect 20636 39678 20638 39730
rect 20690 39678 20692 39730
rect 19628 38894 19630 38946
rect 19682 38894 19684 38946
rect 19628 38882 19684 38894
rect 20188 38834 20244 38846
rect 20188 38782 20190 38834
rect 20242 38782 20244 38834
rect 19516 38724 19572 38734
rect 19292 38612 19460 38668
rect 19516 38630 19572 38668
rect 19068 37214 19070 37266
rect 19122 37214 19124 37266
rect 19068 36372 19124 37214
rect 19068 36306 19124 36316
rect 18844 33282 18900 33292
rect 18956 36260 19012 36270
rect 18172 32788 18228 32798
rect 18060 32786 18228 32788
rect 18060 32734 18174 32786
rect 18226 32734 18228 32786
rect 18060 32732 18228 32734
rect 18060 32564 18116 32574
rect 18060 32470 18116 32508
rect 17724 32452 17780 32462
rect 17612 32450 17780 32452
rect 17612 32398 17726 32450
rect 17778 32398 17780 32450
rect 17612 32396 17780 32398
rect 17052 31668 17108 31678
rect 16940 31666 17108 31668
rect 16940 31614 17054 31666
rect 17106 31614 17108 31666
rect 16940 31612 17108 31614
rect 17052 31556 17108 31612
rect 17052 31490 17108 31500
rect 17276 31108 17332 31118
rect 17164 31052 17276 31108
rect 16716 30158 16718 30210
rect 16770 30158 16772 30210
rect 16716 30146 16772 30158
rect 16940 30212 16996 30222
rect 16940 30118 16996 30156
rect 17052 30210 17108 30222
rect 17052 30158 17054 30210
rect 17106 30158 17108 30210
rect 17052 29988 17108 30158
rect 17052 29922 17108 29932
rect 16716 29538 16772 29550
rect 16716 29486 16718 29538
rect 16770 29486 16772 29538
rect 16604 29428 16660 29438
rect 16604 29334 16660 29372
rect 16604 28420 16660 28430
rect 16716 28420 16772 29486
rect 17052 29540 17108 29550
rect 16940 29428 16996 29438
rect 16940 29334 16996 29372
rect 17052 29204 17108 29484
rect 16940 29148 17108 29204
rect 16940 28532 16996 29148
rect 16940 28530 17108 28532
rect 16940 28478 16942 28530
rect 16994 28478 17108 28530
rect 16940 28476 17108 28478
rect 16940 28466 16996 28476
rect 16660 28364 16772 28420
rect 16604 28326 16660 28364
rect 16492 27244 16660 27300
rect 16492 27076 16548 27086
rect 16380 27074 16548 27076
rect 16380 27022 16494 27074
rect 16546 27022 16548 27074
rect 16380 27020 16548 27022
rect 15932 26982 15988 27020
rect 15708 26898 15764 26908
rect 16156 26964 16212 26974
rect 16156 26850 16212 26908
rect 16268 26962 16324 26974
rect 16268 26910 16270 26962
rect 16322 26910 16324 26962
rect 16268 26908 16324 26910
rect 16268 26852 16436 26908
rect 16156 26798 16158 26850
rect 16210 26798 16212 26850
rect 16156 26786 16212 26798
rect 16380 26740 16436 26852
rect 16492 26852 16548 27020
rect 16604 27020 16660 27244
rect 16716 27188 16772 27198
rect 16716 27094 16772 27132
rect 16604 26964 16772 27020
rect 16940 26964 16996 26974
rect 16716 26962 16996 26964
rect 16716 26910 16942 26962
rect 16994 26910 16996 26962
rect 16716 26908 16996 26910
rect 16940 26898 16996 26908
rect 17052 26908 17108 28476
rect 17164 27074 17220 31052
rect 17276 31042 17332 31052
rect 17612 30324 17668 30334
rect 17276 30322 17668 30324
rect 17276 30270 17614 30322
rect 17666 30270 17668 30322
rect 17276 30268 17668 30270
rect 17276 29428 17332 30268
rect 17612 30258 17668 30268
rect 17724 30324 17780 32396
rect 17724 30258 17780 30268
rect 18060 30322 18116 30334
rect 18060 30270 18062 30322
rect 18114 30270 18116 30322
rect 17388 30098 17444 30110
rect 17388 30046 17390 30098
rect 17442 30046 17444 30098
rect 17388 29764 17444 30046
rect 17388 29698 17444 29708
rect 17500 29986 17556 29998
rect 17500 29934 17502 29986
rect 17554 29934 17556 29986
rect 17500 29652 17556 29934
rect 18060 29988 18116 30270
rect 18060 29922 18116 29932
rect 17612 29876 17668 29886
rect 17668 29820 17780 29876
rect 17612 29810 17668 29820
rect 17500 29586 17556 29596
rect 17724 29650 17780 29820
rect 17724 29598 17726 29650
rect 17778 29598 17780 29650
rect 17724 29586 17780 29598
rect 17836 29540 17892 29550
rect 17836 29446 17892 29484
rect 18060 29540 18116 29550
rect 18060 29446 18116 29484
rect 17388 29428 17444 29438
rect 17276 29426 17444 29428
rect 17276 29374 17390 29426
rect 17442 29374 17444 29426
rect 17276 29372 17444 29374
rect 17276 28196 17332 29372
rect 17388 29362 17444 29372
rect 17612 29426 17668 29438
rect 17612 29374 17614 29426
rect 17666 29374 17668 29426
rect 17612 29316 17668 29374
rect 17612 29250 17668 29260
rect 17948 29204 18004 29214
rect 17948 28868 18004 29148
rect 17836 28866 18004 28868
rect 17836 28814 17950 28866
rect 18002 28814 18004 28866
rect 17836 28812 18004 28814
rect 17388 28644 17444 28654
rect 17724 28644 17780 28654
rect 17444 28642 17780 28644
rect 17444 28590 17726 28642
rect 17778 28590 17780 28642
rect 17444 28588 17780 28590
rect 17388 28550 17444 28588
rect 17724 28578 17780 28588
rect 17836 28196 17892 28812
rect 17948 28802 18004 28812
rect 18172 28420 18228 32732
rect 18620 32564 18676 32574
rect 18620 32470 18676 32508
rect 18396 29988 18452 29998
rect 18396 29894 18452 29932
rect 18508 29316 18564 29326
rect 18564 29260 18676 29316
rect 18508 29222 18564 29260
rect 18508 29092 18564 29102
rect 18284 28644 18340 28654
rect 18284 28550 18340 28588
rect 18172 28364 18452 28420
rect 17276 28130 17332 28140
rect 17500 28140 17892 28196
rect 17500 28084 17556 28140
rect 17388 28082 17556 28084
rect 17388 28030 17502 28082
rect 17554 28030 17556 28082
rect 17388 28028 17556 28030
rect 17388 27076 17444 28028
rect 17500 28018 17556 28028
rect 18060 27972 18116 27982
rect 17164 27022 17166 27074
rect 17218 27022 17220 27074
rect 17164 27010 17220 27022
rect 17276 27020 17444 27076
rect 17612 27748 17668 27758
rect 17052 26852 17220 26908
rect 16492 26796 16772 26852
rect 16380 26684 16660 26740
rect 15932 26628 15988 26638
rect 15820 26404 15876 26414
rect 15820 26310 15876 26348
rect 15596 26226 15652 26236
rect 15820 26180 15876 26190
rect 15260 25564 15652 25620
rect 15596 25506 15652 25564
rect 15596 25454 15598 25506
rect 15650 25454 15652 25506
rect 15596 25442 15652 25454
rect 15708 25394 15764 25406
rect 15708 25342 15710 25394
rect 15762 25342 15764 25394
rect 15260 25284 15316 25294
rect 15708 25284 15764 25342
rect 15260 25282 15764 25284
rect 15260 25230 15262 25282
rect 15314 25230 15764 25282
rect 15260 25228 15764 25230
rect 15260 25218 15316 25228
rect 14924 25060 14980 25070
rect 15484 25060 15540 25070
rect 14980 25004 15204 25060
rect 14924 24994 14980 25004
rect 15148 24946 15204 25004
rect 15148 24894 15150 24946
rect 15202 24894 15204 24946
rect 15148 24882 15204 24894
rect 15260 24948 15316 24958
rect 15260 24854 15316 24892
rect 15484 24834 15540 25004
rect 15484 24782 15486 24834
rect 15538 24782 15540 24834
rect 15484 24770 15540 24782
rect 14812 24724 14868 24734
rect 14812 24630 14868 24668
rect 15036 24722 15092 24734
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 14588 24610 14644 24622
rect 14588 24558 14590 24610
rect 14642 24558 14644 24610
rect 14588 24500 14644 24558
rect 15036 24500 15092 24670
rect 14588 24444 15092 24500
rect 15036 23716 15092 24444
rect 15484 23828 15540 23838
rect 15260 23826 15540 23828
rect 15260 23774 15486 23826
rect 15538 23774 15540 23826
rect 15260 23772 15540 23774
rect 14812 23660 15092 23716
rect 15148 23716 15204 23726
rect 15260 23716 15316 23772
rect 15484 23762 15540 23772
rect 15148 23714 15316 23716
rect 15148 23662 15150 23714
rect 15202 23662 15316 23714
rect 15148 23660 15316 23662
rect 14476 22820 14532 22830
rect 14476 21700 14532 22764
rect 14700 22596 14756 22606
rect 14476 21634 14532 21644
rect 14588 22260 14644 22270
rect 14588 22146 14644 22204
rect 14588 22094 14590 22146
rect 14642 22094 14644 22146
rect 14588 21924 14644 22094
rect 14364 21410 14420 21420
rect 14252 20862 14254 20914
rect 14306 20862 14308 20914
rect 14252 20850 14308 20862
rect 14140 20636 14420 20692
rect 14028 20300 14196 20356
rect 13804 20178 13860 20188
rect 13916 20132 13972 20142
rect 13916 20038 13972 20076
rect 13692 19394 13748 19404
rect 13804 19796 13860 19806
rect 13580 19236 13636 19246
rect 13580 19142 13636 19180
rect 13692 19010 13748 19022
rect 13692 18958 13694 19010
rect 13746 18958 13748 19010
rect 13692 18900 13748 18958
rect 13692 18834 13748 18844
rect 13468 18386 13524 18396
rect 13692 18450 13748 18462
rect 13692 18398 13694 18450
rect 13746 18398 13748 18450
rect 13692 18228 13748 18398
rect 13804 18452 13860 19740
rect 13916 19348 13972 19358
rect 13916 19234 13972 19292
rect 14028 19348 14084 19358
rect 14140 19348 14196 20300
rect 14364 20132 14420 20636
rect 14588 20690 14644 21868
rect 14588 20638 14590 20690
rect 14642 20638 14644 20690
rect 14588 20626 14644 20638
rect 14476 20580 14532 20590
rect 14476 20486 14532 20524
rect 14028 19346 14196 19348
rect 14028 19294 14030 19346
rect 14082 19294 14196 19346
rect 14028 19292 14196 19294
rect 14252 20018 14308 20030
rect 14252 19966 14254 20018
rect 14306 19966 14308 20018
rect 14028 19282 14084 19292
rect 13916 19182 13918 19234
rect 13970 19182 13972 19234
rect 13916 19170 13972 19182
rect 14252 19122 14308 19966
rect 14252 19070 14254 19122
rect 14306 19070 14308 19122
rect 14252 19058 14308 19070
rect 14028 19010 14084 19022
rect 14028 18958 14030 19010
rect 14082 18958 14084 19010
rect 14028 18676 14084 18958
rect 14028 18610 14084 18620
rect 14252 18452 14308 18462
rect 13804 18396 14196 18452
rect 14028 18228 14084 18238
rect 13692 18226 14084 18228
rect 13692 18174 14030 18226
rect 14082 18174 14084 18226
rect 13692 18172 14084 18174
rect 14028 18162 14084 18172
rect 14140 17778 14196 18396
rect 14252 18358 14308 18396
rect 14364 18004 14420 20076
rect 14700 19796 14756 22540
rect 14812 21700 14868 23660
rect 15148 23492 15204 23660
rect 15708 23548 15764 25228
rect 15148 22820 15204 23436
rect 15148 22754 15204 22764
rect 15372 23492 15764 23548
rect 15036 22484 15092 22494
rect 15036 22372 15092 22428
rect 15036 22316 15204 22372
rect 14924 22260 14980 22270
rect 14924 22166 14980 22204
rect 15036 22146 15092 22158
rect 15036 22094 15038 22146
rect 15090 22094 15092 22146
rect 15036 22036 15092 22094
rect 14812 21634 14868 21644
rect 14924 21980 15092 22036
rect 14924 21476 14980 21980
rect 15148 21924 15204 22316
rect 14924 21410 14980 21420
rect 15036 21868 15204 21924
rect 15260 22146 15316 22158
rect 15260 22094 15262 22146
rect 15314 22094 15316 22146
rect 14812 20804 14868 20814
rect 14812 20242 14868 20748
rect 14812 20190 14814 20242
rect 14866 20190 14868 20242
rect 14812 20178 14868 20190
rect 14924 20802 14980 20814
rect 14924 20750 14926 20802
rect 14978 20750 14980 20802
rect 14924 20020 14980 20750
rect 14924 19954 14980 19964
rect 14700 19730 14756 19740
rect 14700 19460 14756 19470
rect 14476 19012 14532 19022
rect 14588 19012 14644 19022
rect 14476 19010 14644 19012
rect 14476 18958 14478 19010
rect 14530 18958 14590 19010
rect 14642 18958 14644 19010
rect 14476 18956 14644 18958
rect 14476 18946 14532 18956
rect 14364 17938 14420 17948
rect 14476 18226 14532 18238
rect 14476 18174 14478 18226
rect 14530 18174 14532 18226
rect 14140 17726 14142 17778
rect 14194 17726 14196 17778
rect 14140 17714 14196 17726
rect 13356 16678 13412 16716
rect 13580 17444 13636 17454
rect 13356 14532 13412 14542
rect 13468 14532 13524 14542
rect 13412 14530 13524 14532
rect 13412 14478 13470 14530
rect 13522 14478 13524 14530
rect 13412 14476 13524 14478
rect 13356 9492 13412 14476
rect 13468 14466 13524 14476
rect 13580 14420 13636 17388
rect 13692 17108 13748 17118
rect 13692 17014 13748 17052
rect 13804 16994 13860 17006
rect 13804 16942 13806 16994
rect 13858 16942 13860 16994
rect 13804 16212 13860 16942
rect 13692 16156 13860 16212
rect 14140 16882 14196 16894
rect 14140 16830 14142 16882
rect 14194 16830 14196 16882
rect 13692 15148 13748 16156
rect 14140 16100 14196 16830
rect 14140 16006 14196 16044
rect 13916 15986 13972 15998
rect 13916 15934 13918 15986
rect 13970 15934 13972 15986
rect 13692 15092 13860 15148
rect 13580 14354 13636 14364
rect 13692 12850 13748 12862
rect 13692 12798 13694 12850
rect 13746 12798 13748 12850
rect 13692 12740 13748 12798
rect 13692 12674 13748 12684
rect 13804 12516 13860 15092
rect 13916 14756 13972 15934
rect 13916 14700 14196 14756
rect 13916 14532 13972 14542
rect 13916 14438 13972 14476
rect 14140 13074 14196 14700
rect 14252 14418 14308 14430
rect 14252 14366 14254 14418
rect 14306 14366 14308 14418
rect 14252 13188 14308 14366
rect 14476 14308 14532 18174
rect 14588 16884 14644 18956
rect 14700 18564 14756 19404
rect 15036 19348 15092 21868
rect 15260 21252 15316 22094
rect 15260 21186 15316 21196
rect 15260 20020 15316 20030
rect 15260 19926 15316 19964
rect 15036 19254 15092 19292
rect 14700 18498 14756 18508
rect 14812 19236 14868 19246
rect 14700 18338 14756 18350
rect 14700 18286 14702 18338
rect 14754 18286 14756 18338
rect 14700 18226 14756 18286
rect 14700 18174 14702 18226
rect 14754 18174 14756 18226
rect 14700 18162 14756 18174
rect 14700 16884 14756 16894
rect 14588 16828 14700 16884
rect 14700 16818 14756 16828
rect 14700 14756 14756 14766
rect 14812 14756 14868 19180
rect 15372 19124 15428 23492
rect 15596 21476 15652 21486
rect 15596 21382 15652 21420
rect 15820 21364 15876 26124
rect 15932 21812 15988 26572
rect 16268 26516 16324 26526
rect 16268 26422 16324 26460
rect 16604 26516 16660 26684
rect 16604 26450 16660 26460
rect 16380 26404 16436 26414
rect 16380 26310 16436 26348
rect 16268 26292 16324 26302
rect 16604 26292 16660 26302
rect 16268 26178 16324 26236
rect 16268 26126 16270 26178
rect 16322 26126 16324 26178
rect 16268 26114 16324 26126
rect 16492 26290 16660 26292
rect 16492 26238 16606 26290
rect 16658 26238 16660 26290
rect 16492 26236 16660 26238
rect 16492 25508 16548 26236
rect 16604 26226 16660 26236
rect 16268 25452 16548 25508
rect 16156 24724 16212 24734
rect 16044 24722 16212 24724
rect 16044 24670 16158 24722
rect 16210 24670 16212 24722
rect 16044 24668 16212 24670
rect 16044 23938 16100 24668
rect 16156 24658 16212 24668
rect 16044 23886 16046 23938
rect 16098 23886 16100 23938
rect 16044 22148 16100 23886
rect 16268 23548 16324 25452
rect 16716 25394 16772 26796
rect 16828 26290 16884 26302
rect 16828 26238 16830 26290
rect 16882 26238 16884 26290
rect 16828 25732 16884 26238
rect 16828 25666 16884 25676
rect 16940 25844 16996 25854
rect 16716 25342 16718 25394
rect 16770 25342 16772 25394
rect 16716 25330 16772 25342
rect 16492 25284 16548 25294
rect 16492 25172 16548 25228
rect 16492 25116 16772 25172
rect 16604 24948 16660 24958
rect 16604 24854 16660 24892
rect 16380 24724 16436 24734
rect 16380 24630 16436 24668
rect 16492 24612 16548 24622
rect 16492 24518 16548 24556
rect 16492 24052 16548 24062
rect 16492 23958 16548 23996
rect 16268 23492 16436 23548
rect 16044 22082 16100 22092
rect 16380 21924 16436 23492
rect 16716 23492 16772 25116
rect 16828 24836 16884 24846
rect 16940 24836 16996 25788
rect 17052 25284 17108 25294
rect 17052 25190 17108 25228
rect 17164 24948 17220 26852
rect 17164 24882 17220 24892
rect 16828 24834 16996 24836
rect 16828 24782 16830 24834
rect 16882 24782 16996 24834
rect 16828 24780 16996 24782
rect 16828 24770 16884 24780
rect 17164 23940 17220 23950
rect 17164 23846 17220 23884
rect 16828 23828 16884 23838
rect 16828 23734 16884 23772
rect 16716 23426 16772 23436
rect 16604 23268 16660 23278
rect 15932 21746 15988 21756
rect 16044 21868 16436 21924
rect 16492 22148 16548 22158
rect 15708 21308 15876 21364
rect 15932 21588 15988 21598
rect 16044 21588 16100 21868
rect 15932 21586 16100 21588
rect 15932 21534 15934 21586
rect 15986 21534 16100 21586
rect 15932 21532 16100 21534
rect 16268 21698 16324 21710
rect 16268 21646 16270 21698
rect 16322 21646 16324 21698
rect 15708 21140 15764 21308
rect 15932 21252 15988 21532
rect 15372 19058 15428 19068
rect 15484 21084 15764 21140
rect 15820 21196 15988 21252
rect 15484 18788 15540 21084
rect 15596 20916 15652 20926
rect 15596 20242 15652 20860
rect 15708 20804 15764 20814
rect 15708 20710 15764 20748
rect 15596 20190 15598 20242
rect 15650 20190 15652 20242
rect 15596 20178 15652 20190
rect 15708 20018 15764 20030
rect 15708 19966 15710 20018
rect 15762 19966 15764 20018
rect 15708 19908 15764 19966
rect 15708 19842 15764 19852
rect 15708 19012 15764 19022
rect 15708 18918 15764 18956
rect 15372 18732 15540 18788
rect 14924 16884 14980 16894
rect 14924 16790 14980 16828
rect 15148 16882 15204 16894
rect 15148 16830 15150 16882
rect 15202 16830 15204 16882
rect 15148 16772 15204 16830
rect 14924 16548 14980 16558
rect 14924 16098 14980 16492
rect 14924 16046 14926 16098
rect 14978 16046 14980 16098
rect 14924 16034 14980 16046
rect 15148 16098 15204 16716
rect 15148 16046 15150 16098
rect 15202 16046 15204 16098
rect 15148 16034 15204 16046
rect 15372 15764 15428 18732
rect 15820 18676 15876 21196
rect 15932 21028 15988 21038
rect 15932 20802 15988 20972
rect 16268 21028 16324 21646
rect 16268 20962 16324 20972
rect 15932 20750 15934 20802
rect 15986 20750 15988 20802
rect 15932 20738 15988 20750
rect 16492 20692 16548 22092
rect 16604 20804 16660 23212
rect 17276 21588 17332 27020
rect 17500 26178 17556 26190
rect 17500 26126 17502 26178
rect 17554 26126 17556 26178
rect 17388 25956 17444 25966
rect 17388 21924 17444 25900
rect 17500 25732 17556 26126
rect 17500 25666 17556 25676
rect 17500 25282 17556 25294
rect 17500 25230 17502 25282
rect 17554 25230 17556 25282
rect 17500 24724 17556 25230
rect 17612 24948 17668 27692
rect 17724 26850 17780 26862
rect 17724 26798 17726 26850
rect 17778 26798 17780 26850
rect 17724 26516 17780 26798
rect 17724 25620 17780 26460
rect 18060 26404 18116 27916
rect 18060 26310 18116 26348
rect 17724 25554 17780 25564
rect 17612 24854 17668 24892
rect 17724 25284 17780 25294
rect 17500 24658 17556 24668
rect 17500 24052 17556 24062
rect 17500 23938 17556 23996
rect 17500 23886 17502 23938
rect 17554 23886 17556 23938
rect 17500 23874 17556 23886
rect 17612 23714 17668 23726
rect 17612 23662 17614 23714
rect 17666 23662 17668 23714
rect 17500 23492 17556 23502
rect 17500 22372 17556 23436
rect 17612 23268 17668 23662
rect 17612 23202 17668 23212
rect 17500 22316 17668 22372
rect 17388 21858 17444 21868
rect 17612 21924 17668 22316
rect 17612 21810 17668 21868
rect 17612 21758 17614 21810
rect 17666 21758 17668 21810
rect 17612 21746 17668 21758
rect 17500 21588 17556 21598
rect 17276 21586 17556 21588
rect 17276 21534 17502 21586
rect 17554 21534 17556 21586
rect 17276 21532 17556 21534
rect 16828 21476 16884 21486
rect 16828 21382 16884 21420
rect 17500 21476 17556 21532
rect 17500 21410 17556 21420
rect 17612 21364 17668 21402
rect 17612 21298 17668 21308
rect 17388 21140 17444 21150
rect 16940 20804 16996 20814
rect 16604 20802 16996 20804
rect 16604 20750 16942 20802
rect 16994 20750 16996 20802
rect 16604 20748 16996 20750
rect 16940 20738 16996 20748
rect 16156 20690 16548 20692
rect 16156 20638 16494 20690
rect 16546 20638 16548 20690
rect 16156 20636 16548 20638
rect 16044 20020 16100 20030
rect 16044 19926 16100 19964
rect 15932 19796 15988 19806
rect 15932 19794 16100 19796
rect 15932 19742 15934 19794
rect 15986 19742 16100 19794
rect 15932 19740 16100 19742
rect 15932 19730 15988 19740
rect 16044 19458 16100 19740
rect 16044 19406 16046 19458
rect 16098 19406 16100 19458
rect 16044 19394 16100 19406
rect 16044 19234 16100 19246
rect 16044 19182 16046 19234
rect 16098 19182 16100 19234
rect 16044 18788 16100 19182
rect 16044 18722 16100 18732
rect 15820 18610 15876 18620
rect 15484 18564 15540 18574
rect 16156 18564 16212 20636
rect 16492 20626 16548 20636
rect 17164 20692 17220 20702
rect 16380 20020 16436 20030
rect 15484 16210 15540 18508
rect 15932 18508 16212 18564
rect 16268 20018 16436 20020
rect 16268 19966 16382 20018
rect 16434 19966 16436 20018
rect 16268 19964 16436 19966
rect 15484 16158 15486 16210
rect 15538 16158 15540 16210
rect 15484 16146 15540 16158
rect 15708 18116 15764 18126
rect 15372 15698 15428 15708
rect 15596 15428 15652 15438
rect 15596 15334 15652 15372
rect 15036 15202 15092 15214
rect 15036 15150 15038 15202
rect 15090 15150 15092 15202
rect 14812 14700 14980 14756
rect 14700 14662 14756 14700
rect 14476 14242 14532 14252
rect 14588 14644 14644 14654
rect 14588 13970 14644 14588
rect 14812 14532 14868 14542
rect 14812 14438 14868 14476
rect 14700 14420 14756 14430
rect 14700 14326 14756 14364
rect 14588 13918 14590 13970
rect 14642 13918 14644 13970
rect 14588 13906 14644 13918
rect 14700 13300 14756 13310
rect 14252 13132 14644 13188
rect 14140 13022 14142 13074
rect 14194 13022 14196 13074
rect 13692 12460 14084 12516
rect 13692 12178 13748 12460
rect 13692 12126 13694 12178
rect 13746 12126 13748 12178
rect 13692 12114 13748 12126
rect 13916 12180 13972 12190
rect 13916 12086 13972 12124
rect 13580 11956 13636 11966
rect 13580 11954 13972 11956
rect 13580 11902 13582 11954
rect 13634 11902 13972 11954
rect 13580 11900 13972 11902
rect 13580 11890 13636 11900
rect 13692 11396 13748 11406
rect 13692 11282 13748 11340
rect 13692 11230 13694 11282
rect 13746 11230 13748 11282
rect 13692 11218 13748 11230
rect 13692 10724 13748 10734
rect 13580 9940 13636 9950
rect 13580 9846 13636 9884
rect 13356 9426 13412 9436
rect 13356 8372 13412 8382
rect 13356 7140 13412 8316
rect 13468 8260 13524 8270
rect 13468 8166 13524 8204
rect 13580 8036 13636 8046
rect 13580 7942 13636 7980
rect 13356 7074 13412 7084
rect 12684 6692 12740 6702
rect 12572 6636 12684 6692
rect 12684 6598 12740 6636
rect 12796 6580 12852 6590
rect 12796 6486 12852 6524
rect 11060 5180 11284 5236
rect 11788 5236 11844 5246
rect 11004 5142 11060 5180
rect 11788 5122 11844 5180
rect 11900 5234 11956 6412
rect 11900 5182 11902 5234
rect 11954 5182 11956 5234
rect 11900 5170 11956 5182
rect 12684 5236 12740 5246
rect 12684 5142 12740 5180
rect 11788 5070 11790 5122
rect 11842 5070 11844 5122
rect 11788 5058 11844 5070
rect 10556 4510 10558 4562
rect 10610 4510 10612 4562
rect 10556 4498 10612 4510
rect 12124 5010 12180 5022
rect 12124 4958 12126 5010
rect 12178 4958 12180 5010
rect 10108 4338 10276 4340
rect 10108 4286 10110 4338
rect 10162 4286 10276 4338
rect 10108 4284 10276 4286
rect 10108 4274 10164 4284
rect 11676 4226 11732 4238
rect 11676 4174 11678 4226
rect 11730 4174 11732 4226
rect 4844 3502 4846 3554
rect 4898 3502 4900 3554
rect 4844 3490 4900 3502
rect 6300 4116 6356 4126
rect 4284 924 4564 980
rect 4508 800 4564 924
rect 6300 800 6356 4060
rect 7420 4116 7476 4126
rect 7420 4022 7476 4060
rect 10220 3668 10276 3678
rect 9884 3666 10276 3668
rect 9884 3614 10222 3666
rect 10274 3614 10276 3666
rect 9884 3612 10276 3614
rect 8764 3556 8820 3566
rect 8764 3462 8820 3500
rect 7756 3332 7812 3342
rect 7756 3330 8148 3332
rect 7756 3278 7758 3330
rect 7810 3278 8148 3330
rect 7756 3276 8148 3278
rect 7756 3266 7812 3276
rect 8092 800 8148 3276
rect 9884 800 9940 3612
rect 10220 3602 10276 3612
rect 11676 800 11732 4174
rect 12124 3554 12180 4958
rect 12908 4338 12964 6860
rect 13244 6850 13300 6860
rect 13020 6692 13076 6702
rect 13468 6692 13524 6702
rect 13020 6690 13524 6692
rect 13020 6638 13022 6690
rect 13074 6638 13470 6690
rect 13522 6638 13524 6690
rect 13020 6636 13524 6638
rect 13020 6626 13076 6636
rect 13468 6626 13524 6636
rect 13692 6580 13748 10668
rect 13804 8034 13860 8046
rect 13804 7982 13806 8034
rect 13858 7982 13860 8034
rect 13804 6690 13860 7982
rect 13916 7476 13972 11900
rect 14028 11284 14084 12460
rect 14028 10498 14084 11228
rect 14028 10446 14030 10498
rect 14082 10446 14084 10498
rect 14028 10434 14084 10446
rect 14140 8372 14196 13022
rect 14252 12962 14308 12974
rect 14252 12910 14254 12962
rect 14306 12910 14308 12962
rect 14252 12852 14308 12910
rect 14252 12786 14308 12796
rect 14140 8306 14196 8316
rect 14476 11396 14532 11406
rect 14476 10834 14532 11340
rect 14476 10782 14478 10834
rect 14530 10782 14532 10834
rect 14364 8148 14420 8158
rect 14140 8036 14196 8046
rect 14364 8036 14420 8092
rect 14140 8034 14420 8036
rect 14140 7982 14142 8034
rect 14194 7982 14420 8034
rect 14140 7980 14420 7982
rect 14140 7970 14196 7980
rect 14140 7476 14196 7486
rect 13916 7420 14084 7476
rect 13804 6638 13806 6690
rect 13858 6638 13860 6690
rect 13804 6626 13860 6638
rect 13916 7140 13972 7150
rect 13580 6524 13692 6580
rect 13468 5236 13524 5246
rect 13580 5236 13636 6524
rect 13692 6514 13748 6524
rect 13804 6468 13860 6478
rect 13804 6374 13860 6412
rect 13804 5796 13860 5806
rect 13916 5796 13972 7084
rect 13804 5794 13972 5796
rect 13804 5742 13806 5794
rect 13858 5742 13972 5794
rect 13804 5740 13972 5742
rect 13804 5730 13860 5740
rect 13468 5234 13636 5236
rect 13468 5182 13470 5234
rect 13522 5182 13636 5234
rect 13468 5180 13636 5182
rect 13468 5170 13524 5180
rect 12908 4286 12910 4338
rect 12962 4286 12964 4338
rect 12908 4274 12964 4286
rect 12124 3502 12126 3554
rect 12178 3502 12180 3554
rect 12124 3490 12180 3502
rect 13468 4116 13524 4126
rect 13468 800 13524 4060
rect 14028 3556 14084 7420
rect 14140 6690 14196 7420
rect 14140 6638 14142 6690
rect 14194 6638 14196 6690
rect 14140 6626 14196 6638
rect 14252 6132 14308 6142
rect 14476 6132 14532 10782
rect 14252 6130 14532 6132
rect 14252 6078 14254 6130
rect 14306 6078 14532 6130
rect 14252 6076 14532 6078
rect 14252 6066 14308 6076
rect 14588 5908 14644 13132
rect 14700 12402 14756 13244
rect 14700 12350 14702 12402
rect 14754 12350 14756 12402
rect 14700 12180 14756 12350
rect 14700 12114 14756 12124
rect 14924 11732 14980 14700
rect 15036 14532 15092 15150
rect 15260 14532 15316 14542
rect 15596 14532 15652 14542
rect 15036 14530 15652 14532
rect 15036 14478 15262 14530
rect 15314 14478 15598 14530
rect 15650 14478 15652 14530
rect 15036 14476 15652 14478
rect 15260 14420 15316 14476
rect 15260 14354 15316 14364
rect 15260 13634 15316 13646
rect 15260 13582 15262 13634
rect 15314 13582 15316 13634
rect 15260 13524 15316 13582
rect 15260 13458 15316 13468
rect 15596 12964 15652 14476
rect 15596 12898 15652 12908
rect 15036 12852 15092 12862
rect 15036 12758 15092 12796
rect 15708 12516 15764 18060
rect 15932 16994 15988 18508
rect 16268 18452 16324 19964
rect 16380 19954 16436 19964
rect 16828 19908 16884 19918
rect 16828 19814 16884 19852
rect 17052 19346 17108 19358
rect 17052 19294 17054 19346
rect 17106 19294 17108 19346
rect 16380 19124 16436 19134
rect 16716 19124 16772 19134
rect 16380 19122 16772 19124
rect 16380 19070 16382 19122
rect 16434 19070 16718 19122
rect 16770 19070 16772 19122
rect 16380 19068 16772 19070
rect 16380 19058 16436 19068
rect 16268 18386 16324 18396
rect 16492 18788 16548 18798
rect 16492 18340 16548 18732
rect 16604 18340 16660 18350
rect 16492 18338 16660 18340
rect 16492 18286 16606 18338
rect 16658 18286 16660 18338
rect 16492 18284 16660 18286
rect 16156 17556 16212 17566
rect 16156 17106 16212 17500
rect 16156 17054 16158 17106
rect 16210 17054 16212 17106
rect 16156 17042 16212 17054
rect 15932 16942 15934 16994
rect 15986 16942 15988 16994
rect 15932 15986 15988 16942
rect 16268 16772 16324 16782
rect 16156 16100 16212 16110
rect 16268 16100 16324 16716
rect 16156 16098 16324 16100
rect 16156 16046 16158 16098
rect 16210 16046 16324 16098
rect 16156 16044 16324 16046
rect 16156 16034 16212 16044
rect 15932 15934 15934 15986
rect 15986 15934 15988 15986
rect 15932 15922 15988 15934
rect 16268 15764 16324 15774
rect 16268 15538 16324 15708
rect 16268 15486 16270 15538
rect 16322 15486 16324 15538
rect 16268 15474 16324 15486
rect 15932 15314 15988 15326
rect 15932 15262 15934 15314
rect 15986 15262 15988 15314
rect 15932 15148 15988 15262
rect 16492 15148 16548 18284
rect 16604 18274 16660 18284
rect 16716 18228 16772 19068
rect 16940 19012 16996 19022
rect 16940 18918 16996 18956
rect 17052 18788 17108 19294
rect 16716 18162 16772 18172
rect 16940 18732 17108 18788
rect 16940 17892 16996 18732
rect 17164 18676 17220 20636
rect 17388 19346 17444 21084
rect 17612 21140 17668 21150
rect 17500 20804 17556 20814
rect 17500 19906 17556 20748
rect 17500 19854 17502 19906
rect 17554 19854 17556 19906
rect 17500 19796 17556 19854
rect 17500 19730 17556 19740
rect 17388 19294 17390 19346
rect 17442 19294 17444 19346
rect 17388 19282 17444 19294
rect 17612 19012 17668 21084
rect 17612 18946 17668 18956
rect 16940 17826 16996 17836
rect 17052 18620 17220 18676
rect 17052 17668 17108 18620
rect 17500 18564 17556 18574
rect 17724 18564 17780 25228
rect 17948 24724 18004 24734
rect 18284 24724 18340 24734
rect 17948 24722 18340 24724
rect 17948 24670 17950 24722
rect 18002 24670 18286 24722
rect 18338 24670 18340 24722
rect 17948 24668 18340 24670
rect 17948 23940 18004 24668
rect 18284 24658 18340 24668
rect 18396 23940 18452 28364
rect 17948 23874 18004 23884
rect 18060 23884 18452 23940
rect 17836 23716 17892 23726
rect 17836 23622 17892 23660
rect 17836 21700 17892 21710
rect 17836 20804 17892 21644
rect 17836 20710 17892 20748
rect 18060 19124 18116 23884
rect 18284 23714 18340 23726
rect 18284 23662 18286 23714
rect 18338 23662 18340 23714
rect 18284 23044 18340 23662
rect 18284 22978 18340 22988
rect 18396 23380 18452 23390
rect 18172 21924 18228 21934
rect 18172 21810 18228 21868
rect 18172 21758 18174 21810
rect 18226 21758 18228 21810
rect 18172 21746 18228 21758
rect 18284 20914 18340 20926
rect 18284 20862 18286 20914
rect 18338 20862 18340 20914
rect 17500 18562 17780 18564
rect 17500 18510 17502 18562
rect 17554 18510 17780 18562
rect 17500 18508 17780 18510
rect 17836 19068 18116 19124
rect 18172 19124 18228 19134
rect 16940 17612 17108 17668
rect 17164 18452 17220 18462
rect 17164 17668 17220 18396
rect 17388 18452 17444 18462
rect 17388 18358 17444 18396
rect 17500 18116 17556 18508
rect 17836 18340 17892 19068
rect 17948 18900 18004 18910
rect 17948 18674 18004 18844
rect 17948 18622 17950 18674
rect 18002 18622 18004 18674
rect 17948 18610 18004 18622
rect 17500 18050 17556 18060
rect 17724 18284 17892 18340
rect 17948 18340 18004 18350
rect 17388 17668 17444 17678
rect 17164 17612 17388 17668
rect 16716 17556 16772 17566
rect 16604 17442 16660 17454
rect 16604 17390 16606 17442
rect 16658 17390 16660 17442
rect 16604 16548 16660 17390
rect 16716 16884 16772 17500
rect 16716 16828 16884 16884
rect 16828 16770 16884 16828
rect 16828 16718 16830 16770
rect 16882 16718 16884 16770
rect 16828 16706 16884 16718
rect 16604 16482 16660 16492
rect 16604 16212 16660 16222
rect 16604 15986 16660 16156
rect 16604 15934 16606 15986
rect 16658 15934 16660 15986
rect 16604 15922 16660 15934
rect 16828 16098 16884 16110
rect 16828 16046 16830 16098
rect 16882 16046 16884 16098
rect 16604 15316 16660 15326
rect 16828 15316 16884 16046
rect 16604 15314 16884 15316
rect 16604 15262 16606 15314
rect 16658 15262 16884 15314
rect 16604 15260 16884 15262
rect 16604 15250 16660 15260
rect 16828 15204 16884 15260
rect 15932 15092 16212 15148
rect 16492 15092 16660 15148
rect 16156 14756 16212 15092
rect 16156 14754 16548 14756
rect 16156 14702 16158 14754
rect 16210 14702 16548 14754
rect 16156 14700 16548 14702
rect 16156 14690 16212 14700
rect 15820 14532 15876 14542
rect 15820 13524 15876 14476
rect 16492 14530 16548 14700
rect 16492 14478 16494 14530
rect 16546 14478 16548 14530
rect 16492 14466 16548 14478
rect 16604 14308 16660 15092
rect 16828 14418 16884 15148
rect 16828 14366 16830 14418
rect 16882 14366 16884 14418
rect 16828 14354 16884 14366
rect 15820 13458 15876 13468
rect 16492 14252 16660 14308
rect 15708 12450 15764 12460
rect 15932 12292 15988 12302
rect 14924 11676 15316 11732
rect 15260 10724 15316 11676
rect 15260 10630 15316 10668
rect 15372 10836 15428 10846
rect 15036 10500 15092 10510
rect 15372 10500 15428 10780
rect 15596 10610 15652 10622
rect 15596 10558 15598 10610
rect 15650 10558 15652 10610
rect 15036 10498 15428 10500
rect 15036 10446 15038 10498
rect 15090 10446 15428 10498
rect 15036 10444 15428 10446
rect 15484 10500 15540 10510
rect 15036 10434 15092 10444
rect 15148 9938 15204 9950
rect 15148 9886 15150 9938
rect 15202 9886 15204 9938
rect 15148 9828 15204 9886
rect 15204 9772 15428 9828
rect 15148 9762 15204 9772
rect 14700 9602 14756 9614
rect 14700 9550 14702 9602
rect 14754 9550 14756 9602
rect 14700 9380 14756 9550
rect 14700 9314 14756 9324
rect 15372 9268 15428 9772
rect 15372 9174 15428 9212
rect 15036 8932 15092 8942
rect 15036 8148 15092 8876
rect 15036 8082 15092 8092
rect 15484 8036 15540 10444
rect 15484 7970 15540 7980
rect 15372 7700 15428 7710
rect 15372 7606 15428 7644
rect 15596 7028 15652 10558
rect 15820 10610 15876 10622
rect 15820 10558 15822 10610
rect 15874 10558 15876 10610
rect 15708 9604 15764 9614
rect 15708 9156 15764 9548
rect 15820 9380 15876 10558
rect 15932 9938 15988 12236
rect 16380 10612 16436 10622
rect 16492 10612 16548 14252
rect 16604 13634 16660 13646
rect 16604 13582 16606 13634
rect 16658 13582 16660 13634
rect 16604 13524 16660 13582
rect 16604 13458 16660 13468
rect 16940 13412 16996 17612
rect 17388 17574 17444 17612
rect 17724 17666 17780 18284
rect 17836 17892 17892 17902
rect 17836 17798 17892 17836
rect 17724 17614 17726 17666
rect 17778 17614 17780 17666
rect 16940 13346 16996 13356
rect 17052 17108 17108 17118
rect 16716 13076 16772 13086
rect 16716 12292 16772 13020
rect 17052 12964 17108 17052
rect 17724 17108 17780 17614
rect 17948 17666 18004 18284
rect 17948 17614 17950 17666
rect 18002 17614 18004 17666
rect 17948 17602 18004 17614
rect 18172 17442 18228 19068
rect 18284 17892 18340 20862
rect 18396 20690 18452 23324
rect 18396 20638 18398 20690
rect 18450 20638 18452 20690
rect 18396 20626 18452 20638
rect 18508 19796 18564 29036
rect 18620 26908 18676 29260
rect 18956 29092 19012 36204
rect 19068 35700 19124 35710
rect 19068 34020 19124 35644
rect 19404 35308 19460 38612
rect 20188 38276 20244 38782
rect 20188 38210 20244 38220
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19516 37380 19572 37390
rect 19516 37286 19572 37324
rect 20076 37380 20132 37390
rect 20132 37324 20244 37380
rect 20076 37314 20132 37324
rect 19292 35252 19460 35308
rect 19628 36148 19684 36158
rect 19180 34020 19236 34030
rect 19068 34018 19180 34020
rect 19068 33966 19070 34018
rect 19122 33966 19180 34018
rect 19068 33964 19180 33966
rect 19068 33954 19124 33964
rect 19068 33236 19124 33246
rect 19068 33142 19124 33180
rect 19068 29540 19124 29550
rect 19068 29446 19124 29484
rect 18956 29026 19012 29036
rect 19180 28868 19236 33964
rect 19292 31108 19348 35252
rect 19628 34242 19684 36092
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20188 35308 20244 37324
rect 20524 36484 20580 36494
rect 20412 36482 20580 36484
rect 20412 36430 20526 36482
rect 20578 36430 20580 36482
rect 20412 36428 20580 36430
rect 20300 36372 20356 36382
rect 20300 36278 20356 36316
rect 20188 35252 20356 35308
rect 20188 34804 20244 34814
rect 20188 34710 20244 34748
rect 20300 34580 20356 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20188 34524 20356 34580
rect 20412 34580 20468 36428
rect 20524 36418 20580 36428
rect 20636 36260 20692 39678
rect 21644 39620 21700 39630
rect 21308 39508 21364 39518
rect 20860 39506 21364 39508
rect 20860 39454 21310 39506
rect 21362 39454 21364 39506
rect 20860 39452 21364 39454
rect 20748 38164 20804 38174
rect 20748 38070 20804 38108
rect 20636 36194 20692 36204
rect 20860 36036 20916 39452
rect 21308 39442 21364 39452
rect 21644 39506 21700 39564
rect 21644 39454 21646 39506
rect 21698 39454 21700 39506
rect 21644 39442 21700 39454
rect 22428 39508 22484 39518
rect 22428 39414 22484 39452
rect 22764 39506 22820 41132
rect 22876 39844 22932 44200
rect 23996 41412 24052 44200
rect 23996 41346 24052 41356
rect 24556 41188 24612 41198
rect 24556 41094 24612 41132
rect 25116 40628 25172 44200
rect 25564 41412 25620 41422
rect 25564 41318 25620 41356
rect 26236 41412 26292 44200
rect 26236 41346 26292 41356
rect 25116 40562 25172 40572
rect 26348 40628 26404 40638
rect 26348 40534 26404 40572
rect 27356 40628 27412 44200
rect 27356 40562 27412 40572
rect 27468 41188 27524 41198
rect 24668 40516 24724 40526
rect 24668 40422 24724 40460
rect 25340 40516 25396 40526
rect 24444 40404 24500 40414
rect 24444 40402 24612 40404
rect 24444 40350 24446 40402
rect 24498 40350 24612 40402
rect 24444 40348 24612 40350
rect 24444 40338 24500 40348
rect 22876 39778 22932 39788
rect 24108 39844 24164 39854
rect 24108 39750 24164 39788
rect 23100 39620 23156 39630
rect 23100 39526 23156 39564
rect 22764 39454 22766 39506
rect 22818 39454 22820 39506
rect 22764 39442 22820 39454
rect 23884 39396 23940 39406
rect 23884 39058 23940 39340
rect 23884 39006 23886 39058
rect 23938 39006 23940 39058
rect 23884 38994 23940 39006
rect 24332 39060 24388 39070
rect 24332 38834 24388 39004
rect 24332 38782 24334 38834
rect 24386 38782 24388 38834
rect 24332 38770 24388 38782
rect 21868 38724 21924 38734
rect 20636 35980 20916 36036
rect 21196 36484 21252 36494
rect 20524 35140 20580 35150
rect 20524 34802 20580 35084
rect 20524 34750 20526 34802
rect 20578 34750 20580 34802
rect 20524 34738 20580 34750
rect 19628 34190 19630 34242
rect 19682 34190 19684 34242
rect 19628 34178 19684 34190
rect 19516 34130 19572 34142
rect 19516 34078 19518 34130
rect 19570 34078 19572 34130
rect 19516 34020 19572 34078
rect 19516 33954 19572 33964
rect 19740 33348 19796 33358
rect 19628 33346 19796 33348
rect 19628 33294 19742 33346
rect 19794 33294 19796 33346
rect 19628 33292 19796 33294
rect 19628 31892 19684 33292
rect 19740 33282 19796 33292
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 31826 19684 31836
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19292 31042 19348 31052
rect 20076 30436 20132 30446
rect 20076 30342 20132 30380
rect 20188 30324 20244 34524
rect 20412 34514 20468 34524
rect 20300 34356 20356 34366
rect 20300 34130 20356 34300
rect 20636 34354 20692 35980
rect 21196 35922 21252 36428
rect 21196 35870 21198 35922
rect 21250 35870 21252 35922
rect 21196 35858 21252 35870
rect 21532 36148 21588 36158
rect 21532 35922 21588 36092
rect 21868 35924 21924 38668
rect 24108 38724 24164 38734
rect 24108 38630 24164 38668
rect 24556 38668 24612 40348
rect 25340 40402 25396 40460
rect 25340 40350 25342 40402
rect 25394 40350 25396 40402
rect 25340 40338 25396 40350
rect 26236 39732 26292 39742
rect 26292 39676 26740 39732
rect 26236 39638 26292 39676
rect 26012 39618 26068 39630
rect 26012 39566 26014 39618
rect 26066 39566 26068 39618
rect 25788 39508 25844 39518
rect 25228 39396 25284 39406
rect 24668 39172 24724 39182
rect 24668 39058 24724 39116
rect 24668 39006 24670 39058
rect 24722 39006 24724 39058
rect 24668 38994 24724 39006
rect 25228 38834 25284 39340
rect 25788 39058 25844 39452
rect 25788 39006 25790 39058
rect 25842 39006 25844 39058
rect 25788 38994 25844 39006
rect 25228 38782 25230 38834
rect 25282 38782 25284 38834
rect 25228 38770 25284 38782
rect 25116 38724 25172 38734
rect 24556 38612 24836 38668
rect 24668 38164 24724 38174
rect 22988 38050 23044 38062
rect 22988 37998 22990 38050
rect 23042 37998 23044 38050
rect 22428 37156 22484 37166
rect 21532 35870 21534 35922
rect 21586 35870 21588 35922
rect 21532 35858 21588 35870
rect 21756 35868 21924 35924
rect 22092 36484 22148 36494
rect 20860 35812 20916 35822
rect 20860 35586 20916 35756
rect 20860 35534 20862 35586
rect 20914 35534 20916 35586
rect 20860 35476 20916 35534
rect 20860 35410 20916 35420
rect 21756 34916 21812 35868
rect 21980 35812 22036 35822
rect 21980 35718 22036 35756
rect 21868 35698 21924 35710
rect 21868 35646 21870 35698
rect 21922 35646 21924 35698
rect 21868 35140 21924 35646
rect 21980 35476 22036 35486
rect 22092 35476 22148 36428
rect 21980 35474 22148 35476
rect 21980 35422 21982 35474
rect 22034 35422 22148 35474
rect 21980 35420 22148 35422
rect 22204 36372 22260 36382
rect 21980 35410 22036 35420
rect 21868 35074 21924 35084
rect 21980 35252 22036 35262
rect 21980 35026 22036 35196
rect 21980 34974 21982 35026
rect 22034 34974 22036 35026
rect 21756 34860 21924 34916
rect 20636 34302 20638 34354
rect 20690 34302 20692 34354
rect 20636 34290 20692 34302
rect 21756 34580 21812 34590
rect 20300 34078 20302 34130
rect 20354 34078 20356 34130
rect 20300 34066 20356 34078
rect 21532 33236 21588 33246
rect 20300 32228 20356 32238
rect 20300 31780 20356 32172
rect 20300 31218 20356 31724
rect 21308 31892 21364 31902
rect 21308 31778 21364 31836
rect 21308 31726 21310 31778
rect 21362 31726 21364 31778
rect 21308 31714 21364 31726
rect 20972 31668 21028 31678
rect 20300 31166 20302 31218
rect 20354 31166 20356 31218
rect 20300 31154 20356 31166
rect 20524 31164 20804 31220
rect 20412 31108 20468 31118
rect 20524 31108 20580 31164
rect 20412 31106 20580 31108
rect 20412 31054 20414 31106
rect 20466 31054 20580 31106
rect 20412 31052 20580 31054
rect 20412 31042 20468 31052
rect 20636 30994 20692 31006
rect 20636 30942 20638 30994
rect 20690 30942 20692 30994
rect 20300 30772 20356 30782
rect 20636 30772 20692 30942
rect 20300 30770 20692 30772
rect 20300 30718 20302 30770
rect 20354 30718 20692 30770
rect 20300 30716 20692 30718
rect 20300 30706 20356 30716
rect 20188 30268 20692 30324
rect 20188 30100 20244 30110
rect 20524 30100 20580 30110
rect 20188 30098 20580 30100
rect 20188 30046 20190 30098
rect 20242 30046 20526 30098
rect 20578 30046 20580 30098
rect 20188 30044 20580 30046
rect 20188 30034 20244 30044
rect 19628 29988 19684 29998
rect 20076 29988 20132 29998
rect 19628 29986 20132 29988
rect 19628 29934 19630 29986
rect 19682 29934 20078 29986
rect 20130 29934 20132 29986
rect 19628 29932 20132 29934
rect 19628 29092 19684 29932
rect 20076 29922 20132 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20412 29428 20468 29438
rect 20412 29334 20468 29372
rect 19628 29026 19684 29036
rect 18956 28812 19236 28868
rect 18620 26852 18788 26908
rect 18620 23940 18676 23950
rect 18620 23846 18676 23884
rect 18508 19740 18676 19796
rect 18396 18450 18452 18462
rect 18396 18398 18398 18450
rect 18450 18398 18452 18450
rect 18396 18340 18452 18398
rect 18396 18274 18452 18284
rect 18508 18228 18564 18238
rect 18284 17836 18452 17892
rect 18172 17390 18174 17442
rect 18226 17390 18228 17442
rect 18172 17378 18228 17390
rect 17724 17042 17780 17052
rect 17948 16996 18004 17006
rect 17948 16902 18004 16940
rect 17612 16884 17668 16894
rect 17612 16770 17668 16828
rect 17612 16718 17614 16770
rect 17666 16718 17668 16770
rect 17276 16660 17332 16670
rect 17164 15204 17220 15214
rect 17164 14530 17220 15148
rect 17164 14478 17166 14530
rect 17218 14478 17220 14530
rect 17164 14466 17220 14478
rect 17276 14418 17332 16604
rect 17388 16436 17444 16446
rect 17388 16212 17444 16380
rect 17612 16436 17668 16718
rect 17612 16370 17668 16380
rect 18172 16882 18228 16894
rect 18172 16830 18174 16882
rect 18226 16830 18228 16882
rect 17724 16212 17780 16222
rect 17388 16210 17780 16212
rect 17388 16158 17390 16210
rect 17442 16158 17726 16210
rect 17778 16158 17780 16210
rect 17388 16156 17780 16158
rect 17388 16146 17444 16156
rect 17500 15652 17556 16156
rect 17724 16146 17780 16156
rect 17500 15538 17556 15596
rect 17948 16098 18004 16110
rect 17948 16046 17950 16098
rect 18002 16046 18004 16098
rect 17500 15486 17502 15538
rect 17554 15486 17556 15538
rect 17500 15474 17556 15486
rect 17724 15540 17780 15550
rect 17724 15446 17780 15484
rect 17948 15428 18004 16046
rect 18172 15540 18228 16830
rect 18284 15876 18340 15886
rect 18284 15782 18340 15820
rect 18284 15540 18340 15550
rect 18172 15484 18284 15540
rect 18284 15474 18340 15484
rect 18060 15428 18116 15438
rect 17948 15372 18060 15428
rect 18060 15334 18116 15372
rect 17388 15314 17444 15326
rect 17388 15262 17390 15314
rect 17442 15262 17444 15314
rect 17388 15204 17444 15262
rect 18396 15148 18452 17836
rect 18508 17666 18564 18172
rect 18508 17614 18510 17666
rect 18562 17614 18564 17666
rect 18508 16996 18564 17614
rect 18508 16930 18564 16940
rect 18508 15652 18564 15662
rect 18508 15538 18564 15596
rect 18508 15486 18510 15538
rect 18562 15486 18564 15538
rect 18508 15474 18564 15486
rect 17388 15138 17444 15148
rect 17276 14366 17278 14418
rect 17330 14366 17332 14418
rect 17276 14354 17332 14366
rect 18284 15092 18452 15148
rect 17500 14306 17556 14318
rect 17500 14254 17502 14306
rect 17554 14254 17556 14306
rect 16716 12198 16772 12236
rect 16940 12908 17108 12964
rect 17164 13188 17220 13198
rect 16828 12180 16884 12218
rect 16828 12114 16884 12124
rect 16940 10836 16996 12908
rect 17052 12740 17108 12750
rect 17164 12740 17220 13132
rect 17388 13188 17444 13198
rect 17500 13188 17556 14254
rect 17724 13860 17780 13870
rect 17724 13766 17780 13804
rect 18060 13860 18116 13870
rect 18060 13766 18116 13804
rect 17388 13186 17556 13188
rect 17388 13134 17390 13186
rect 17442 13134 17556 13186
rect 17388 13132 17556 13134
rect 17388 13122 17444 13132
rect 17052 12738 17220 12740
rect 17052 12686 17054 12738
rect 17106 12686 17220 12738
rect 17052 12684 17220 12686
rect 17052 12674 17108 12684
rect 17276 12516 17332 12526
rect 17276 11172 17332 12460
rect 17276 11106 17332 11116
rect 17388 10836 17444 10846
rect 16940 10770 16996 10780
rect 17052 10780 17388 10836
rect 16380 10610 16548 10612
rect 16380 10558 16382 10610
rect 16434 10558 16548 10610
rect 16380 10556 16548 10558
rect 16380 10546 16436 10556
rect 15932 9886 15934 9938
rect 15986 9886 15988 9938
rect 15932 9874 15988 9886
rect 15820 9314 15876 9324
rect 16156 9268 16212 9278
rect 17052 9268 17108 10780
rect 17388 10742 17444 10780
rect 17500 10612 17556 13132
rect 17612 13188 17668 13198
rect 17612 12850 17668 13132
rect 17612 12798 17614 12850
rect 17666 12798 17668 12850
rect 17612 12786 17668 12798
rect 17724 13074 17780 13086
rect 17724 13022 17726 13074
rect 17778 13022 17780 13074
rect 17612 12404 17668 12414
rect 17612 12178 17668 12348
rect 17612 12126 17614 12178
rect 17666 12126 17668 12178
rect 17612 12114 17668 12126
rect 17724 12178 17780 13022
rect 17724 12126 17726 12178
rect 17778 12126 17780 12178
rect 17724 12114 17780 12126
rect 17836 12180 17892 12190
rect 17836 12086 17892 12124
rect 18172 12178 18228 12190
rect 18172 12126 18174 12178
rect 18226 12126 18228 12178
rect 18060 12066 18116 12078
rect 18060 12014 18062 12066
rect 18114 12014 18116 12066
rect 17612 10612 17668 10622
rect 17500 10556 17612 10612
rect 17612 10518 17668 10556
rect 18060 9938 18116 12014
rect 18172 10836 18228 12126
rect 18172 10770 18228 10780
rect 18060 9886 18062 9938
rect 18114 9886 18116 9938
rect 18060 9874 18116 9886
rect 18284 9716 18340 15092
rect 18620 13746 18676 19740
rect 18732 19236 18788 26852
rect 18844 24836 18900 24846
rect 18844 24612 18900 24780
rect 18844 24518 18900 24556
rect 18844 20804 18900 20814
rect 18844 20710 18900 20748
rect 18732 18788 18788 19180
rect 18732 18722 18788 18732
rect 18956 18676 19012 28812
rect 20188 28756 20244 28766
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20188 26852 20244 28700
rect 20300 28420 20356 28430
rect 20524 28420 20580 30044
rect 20636 30098 20692 30268
rect 20636 30046 20638 30098
rect 20690 30046 20692 30098
rect 20636 29764 20692 30046
rect 20636 29698 20692 29708
rect 20748 30100 20804 31164
rect 20972 31218 21028 31612
rect 20972 31166 20974 31218
rect 21026 31166 21028 31218
rect 20972 31154 21028 31166
rect 20860 30996 20916 31006
rect 20860 30210 20916 30940
rect 20972 30994 21028 31006
rect 20972 30942 20974 30994
rect 21026 30942 21028 30994
rect 20972 30436 21028 30942
rect 21308 30994 21364 31006
rect 21308 30942 21310 30994
rect 21362 30942 21364 30994
rect 21308 30884 21364 30942
rect 21308 30818 21364 30828
rect 20972 30370 21028 30380
rect 20860 30158 20862 30210
rect 20914 30158 20916 30210
rect 20860 30146 20916 30158
rect 20748 29650 20804 30044
rect 21196 29764 21252 29774
rect 21196 29652 21252 29708
rect 20748 29598 20750 29650
rect 20802 29598 20804 29650
rect 20636 28644 20692 28654
rect 20636 28550 20692 28588
rect 20300 28418 20580 28420
rect 20300 28366 20302 28418
rect 20354 28366 20580 28418
rect 20300 28364 20580 28366
rect 20300 26908 20356 28364
rect 20748 28308 20804 29598
rect 20524 28252 20804 28308
rect 20972 29650 21252 29652
rect 20972 29598 21198 29650
rect 21250 29598 21252 29650
rect 20972 29596 21252 29598
rect 20524 27076 20580 28252
rect 20524 27010 20580 27020
rect 20636 26962 20692 26974
rect 20636 26910 20638 26962
rect 20690 26910 20692 26962
rect 20300 26852 20580 26908
rect 20188 26786 20244 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26180 19684 26190
rect 19628 25396 19684 26124
rect 20524 25508 20580 26852
rect 20636 26180 20692 26910
rect 20860 26850 20916 26862
rect 20860 26798 20862 26850
rect 20914 26798 20916 26850
rect 20860 26292 20916 26798
rect 20860 26226 20916 26236
rect 20636 26114 20692 26124
rect 20524 25414 20580 25452
rect 19628 25330 19684 25340
rect 20412 25396 20468 25406
rect 19068 25284 19124 25294
rect 19068 18900 19124 25228
rect 19852 25284 19908 25322
rect 19852 25218 19908 25228
rect 20300 25284 20356 25294
rect 20412 25284 20468 25340
rect 20636 25284 20692 25294
rect 20300 25282 20580 25284
rect 20300 25230 20302 25282
rect 20354 25230 20580 25282
rect 20300 25228 20580 25230
rect 20300 25218 20356 25228
rect 20188 25172 20244 25182
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20076 24948 20132 24958
rect 20188 24948 20244 25116
rect 19628 24946 20468 24948
rect 19628 24894 20078 24946
rect 20130 24894 20468 24946
rect 19628 24892 20468 24894
rect 19292 24834 19348 24846
rect 19292 24782 19294 24834
rect 19346 24782 19348 24834
rect 19292 23940 19348 24782
rect 19628 24834 19684 24892
rect 20076 24882 20132 24892
rect 19628 24782 19630 24834
rect 19682 24782 19684 24834
rect 19628 24770 19684 24782
rect 19292 23874 19348 23884
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23492 20244 23502
rect 20188 23378 20244 23436
rect 20188 23326 20190 23378
rect 20242 23326 20244 23378
rect 20188 23314 20244 23326
rect 19292 23268 19348 23278
rect 19180 23212 19292 23268
rect 19180 19908 19236 23212
rect 19292 23202 19348 23212
rect 20076 23268 20132 23278
rect 20076 23174 20132 23212
rect 19516 22708 19572 22718
rect 19404 22652 19516 22708
rect 19292 21812 19348 21822
rect 19292 21698 19348 21756
rect 19292 21646 19294 21698
rect 19346 21646 19348 21698
rect 19292 21634 19348 21646
rect 19292 19908 19348 19918
rect 19180 19906 19348 19908
rect 19180 19854 19294 19906
rect 19346 19854 19348 19906
rect 19180 19852 19348 19854
rect 19292 19842 19348 19852
rect 19404 18900 19460 22652
rect 19516 22642 19572 22652
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 19908 20244 19918
rect 19628 19684 19684 19694
rect 19516 19124 19572 19134
rect 19516 19030 19572 19068
rect 19404 18844 19572 18900
rect 19068 18834 19124 18844
rect 18844 18620 19012 18676
rect 18844 18228 18900 18620
rect 18956 18452 19012 18462
rect 19404 18452 19460 18462
rect 18956 18450 19460 18452
rect 18956 18398 18958 18450
rect 19010 18398 19406 18450
rect 19458 18398 19460 18450
rect 18956 18396 19460 18398
rect 18956 18386 19012 18396
rect 19404 18386 19460 18396
rect 19292 18228 19348 18238
rect 18844 18172 19012 18228
rect 18844 17668 18900 17678
rect 18844 17554 18900 17612
rect 18844 17502 18846 17554
rect 18898 17502 18900 17554
rect 18732 17108 18788 17118
rect 18732 17014 18788 17052
rect 18620 13694 18622 13746
rect 18674 13694 18676 13746
rect 16156 9174 16212 9212
rect 16828 9212 17108 9268
rect 17500 9660 18340 9716
rect 18396 13412 18452 13422
rect 15820 9156 15876 9166
rect 15708 9100 15820 9156
rect 15820 9062 15876 9100
rect 16716 9156 16772 9166
rect 16716 9062 16772 9100
rect 16268 9044 16324 9054
rect 16604 9044 16660 9054
rect 16268 9042 16660 9044
rect 16268 8990 16270 9042
rect 16322 8990 16606 9042
rect 16658 8990 16660 9042
rect 16268 8988 16660 8990
rect 16268 8978 16324 8988
rect 16156 8820 16212 8830
rect 16156 8818 16548 8820
rect 16156 8766 16158 8818
rect 16210 8766 16548 8818
rect 16156 8764 16548 8766
rect 16156 8754 16212 8764
rect 15820 8708 15876 8718
rect 15820 8370 15876 8652
rect 15820 8318 15822 8370
rect 15874 8318 15876 8370
rect 15820 8306 15876 8318
rect 16268 8372 16324 8382
rect 16268 8278 16324 8316
rect 15932 8148 15988 8158
rect 15820 7700 15876 7710
rect 15820 7606 15876 7644
rect 15932 7586 15988 8092
rect 15932 7534 15934 7586
rect 15986 7534 15988 7586
rect 15932 7522 15988 7534
rect 16156 7474 16212 7486
rect 16156 7422 16158 7474
rect 16210 7422 16212 7474
rect 15820 7252 15876 7262
rect 16156 7252 16212 7422
rect 16492 7474 16548 8764
rect 16604 8372 16660 8988
rect 16604 8306 16660 8316
rect 16716 8708 16772 8718
rect 16492 7422 16494 7474
rect 16546 7422 16548 7474
rect 16492 7410 16548 7422
rect 16604 8148 16660 8158
rect 16380 7364 16436 7374
rect 15820 7250 16212 7252
rect 15820 7198 15822 7250
rect 15874 7198 16212 7250
rect 15820 7196 16212 7198
rect 16268 7362 16436 7364
rect 16268 7310 16382 7362
rect 16434 7310 16436 7362
rect 16268 7308 16436 7310
rect 15820 7186 15876 7196
rect 15596 6972 15764 7028
rect 15148 6692 15204 6702
rect 15148 6598 15204 6636
rect 14140 5852 14644 5908
rect 15596 6468 15652 6478
rect 14140 4338 14196 5852
rect 15596 5234 15652 6412
rect 15596 5182 15598 5234
rect 15650 5182 15652 5234
rect 15596 5170 15652 5182
rect 14140 4286 14142 4338
rect 14194 4286 14196 4338
rect 14140 4274 14196 4286
rect 14700 4116 14756 4126
rect 14700 4022 14756 4060
rect 15708 3556 15764 6972
rect 16268 6916 16324 7308
rect 16380 7298 16436 7308
rect 16604 7364 16660 8092
rect 16716 8146 16772 8652
rect 16716 8094 16718 8146
rect 16770 8094 16772 8146
rect 16716 8082 16772 8094
rect 16828 8148 16884 9212
rect 16940 9044 16996 9054
rect 16940 9042 17444 9044
rect 16940 8990 16942 9042
rect 16994 8990 17444 9042
rect 16940 8988 17444 8990
rect 16940 8978 16996 8988
rect 17388 8258 17444 8988
rect 17388 8206 17390 8258
rect 17442 8206 17444 8258
rect 17388 8194 17444 8206
rect 16828 8082 16884 8092
rect 17164 8146 17220 8158
rect 17164 8094 17166 8146
rect 17218 8094 17220 8146
rect 16940 8036 16996 8046
rect 16940 7942 16996 7980
rect 17164 7588 17220 8094
rect 16828 7476 16884 7486
rect 17164 7476 17220 7532
rect 17388 7924 17444 7934
rect 17388 7586 17444 7868
rect 17388 7534 17390 7586
rect 17442 7534 17444 7586
rect 17388 7522 17444 7534
rect 16884 7420 17220 7476
rect 16828 7382 16884 7420
rect 16604 7298 16660 7308
rect 15820 6860 16324 6916
rect 15820 6802 15876 6860
rect 15820 6750 15822 6802
rect 15874 6750 15876 6802
rect 15820 6738 15876 6750
rect 17500 5906 17556 9660
rect 17836 8258 17892 8270
rect 17836 8206 17838 8258
rect 17890 8206 17892 8258
rect 17612 8034 17668 8046
rect 17612 7982 17614 8034
rect 17666 7982 17668 8034
rect 17612 7028 17668 7982
rect 17836 7812 17892 8206
rect 18396 7924 18452 13356
rect 18508 13076 18564 13086
rect 18508 12982 18564 13020
rect 18620 12628 18676 13694
rect 18732 16884 18788 16894
rect 18732 12740 18788 16828
rect 18844 15988 18900 17502
rect 18956 16212 19012 18172
rect 19292 18134 19348 18172
rect 19068 18116 19124 18126
rect 19124 18060 19236 18116
rect 19068 18050 19124 18060
rect 19180 17780 19236 18060
rect 19292 17780 19348 17790
rect 19180 17778 19348 17780
rect 19180 17726 19294 17778
rect 19346 17726 19348 17778
rect 19180 17724 19348 17726
rect 19292 17714 19348 17724
rect 18956 16210 19460 16212
rect 18956 16158 18958 16210
rect 19010 16158 19460 16210
rect 18956 16156 19460 16158
rect 18956 16146 19012 16156
rect 19292 15988 19348 15998
rect 18844 15986 19348 15988
rect 18844 15934 19294 15986
rect 19346 15934 19348 15986
rect 18844 15932 19348 15934
rect 19292 15922 19348 15932
rect 19404 15986 19460 16156
rect 19404 15934 19406 15986
rect 19458 15934 19460 15986
rect 18844 15764 18900 15774
rect 18844 13076 18900 15708
rect 19404 15148 19460 15934
rect 19068 15092 19460 15148
rect 19068 14084 19124 15092
rect 19068 13970 19124 14028
rect 19068 13918 19070 13970
rect 19122 13918 19124 13970
rect 19068 13906 19124 13918
rect 19292 13076 19348 13086
rect 18844 13074 19348 13076
rect 18844 13022 19294 13074
rect 19346 13022 19348 13074
rect 18844 13020 19348 13022
rect 18844 12962 18900 13020
rect 19292 13010 19348 13020
rect 18844 12910 18846 12962
rect 18898 12910 18900 12962
rect 18844 12898 18900 12910
rect 19180 12852 19236 12862
rect 19180 12850 19348 12852
rect 19180 12798 19182 12850
rect 19234 12798 19348 12850
rect 19180 12796 19348 12798
rect 19180 12786 19236 12796
rect 18732 12674 18788 12684
rect 18508 12572 18676 12628
rect 18508 9940 18564 12572
rect 18620 12404 18676 12414
rect 18620 12310 18676 12348
rect 18732 11394 18788 11406
rect 18732 11342 18734 11394
rect 18786 11342 18788 11394
rect 18732 11172 18788 11342
rect 19180 11172 19236 11182
rect 18732 11170 19236 11172
rect 18732 11118 19182 11170
rect 19234 11118 19236 11170
rect 18732 11116 19236 11118
rect 19180 10164 19236 11116
rect 19180 10098 19236 10108
rect 18508 8596 18564 9884
rect 18732 9826 18788 9838
rect 18732 9774 18734 9826
rect 18786 9774 18788 9826
rect 18732 9156 18788 9774
rect 19292 9156 19348 12796
rect 19404 10612 19460 10622
rect 19404 10518 19460 10556
rect 18732 9154 18900 9156
rect 18732 9102 18734 9154
rect 18786 9102 18900 9154
rect 18732 9100 18900 9102
rect 19292 9100 19460 9156
rect 18732 9090 18788 9100
rect 18508 8530 18564 8540
rect 18732 8372 18788 8382
rect 18508 8260 18564 8270
rect 18508 8166 18564 8204
rect 18732 8146 18788 8316
rect 18732 8094 18734 8146
rect 18786 8094 18788 8146
rect 18732 8082 18788 8094
rect 17836 7746 17892 7756
rect 18172 7868 18452 7924
rect 18620 8036 18676 8046
rect 18172 7700 18228 7868
rect 18172 7634 18228 7644
rect 17724 7588 17780 7598
rect 18060 7588 18116 7598
rect 17780 7586 18116 7588
rect 17780 7534 18062 7586
rect 18114 7534 18116 7586
rect 17780 7532 18116 7534
rect 17724 7494 17780 7532
rect 18060 7522 18116 7532
rect 17612 6972 18228 7028
rect 17948 6804 18004 6814
rect 17948 6710 18004 6748
rect 17500 5854 17502 5906
rect 17554 5854 17556 5906
rect 17500 5842 17556 5854
rect 17836 6692 17892 6702
rect 17052 5684 17108 5694
rect 16380 5124 16436 5134
rect 16380 5030 16436 5068
rect 15932 3556 15988 3566
rect 15708 3554 15988 3556
rect 15708 3502 15934 3554
rect 15986 3502 15988 3554
rect 15708 3500 15988 3502
rect 14028 3490 14084 3500
rect 15932 3490 15988 3500
rect 15372 3332 15428 3342
rect 15260 3330 15428 3332
rect 15260 3278 15374 3330
rect 15426 3278 15428 3330
rect 15260 3276 15428 3278
rect 15260 800 15316 3276
rect 15372 3266 15428 3276
rect 17052 800 17108 5628
rect 17500 5124 17556 5134
rect 17836 5124 17892 6636
rect 17556 5122 17892 5124
rect 17556 5070 17838 5122
rect 17890 5070 17892 5122
rect 17556 5068 17892 5070
rect 17500 4338 17556 5068
rect 17836 5058 17892 5068
rect 18172 4450 18228 6972
rect 18284 6804 18340 7868
rect 18396 7700 18452 7710
rect 18396 7474 18452 7644
rect 18620 7586 18676 7980
rect 18620 7534 18622 7586
rect 18674 7534 18676 7586
rect 18620 7522 18676 7534
rect 18396 7422 18398 7474
rect 18450 7422 18452 7474
rect 18396 7410 18452 7422
rect 18284 6738 18340 6748
rect 18508 7362 18564 7374
rect 18508 7310 18510 7362
rect 18562 7310 18564 7362
rect 18396 5684 18452 5694
rect 18396 5590 18452 5628
rect 18508 5236 18564 7310
rect 18844 6692 18900 9100
rect 19180 8596 19236 8606
rect 19068 8484 19124 8494
rect 18956 8034 19012 8046
rect 18956 7982 18958 8034
rect 19010 7982 19012 8034
rect 18956 7700 19012 7982
rect 18956 7634 19012 7644
rect 19068 7698 19124 8428
rect 19068 7646 19070 7698
rect 19122 7646 19124 7698
rect 19068 7634 19124 7646
rect 19180 8146 19236 8540
rect 19292 8372 19348 8382
rect 19292 8258 19348 8316
rect 19292 8206 19294 8258
rect 19346 8206 19348 8258
rect 19292 8194 19348 8206
rect 19180 8094 19182 8146
rect 19234 8094 19236 8146
rect 18956 7474 19012 7486
rect 18956 7422 18958 7474
rect 19010 7422 19012 7474
rect 18956 7364 19012 7422
rect 18956 7298 19012 7308
rect 19180 7028 19236 8094
rect 19292 7812 19348 7822
rect 19292 7698 19348 7756
rect 19292 7646 19294 7698
rect 19346 7646 19348 7698
rect 19292 7634 19348 7646
rect 18844 6626 18900 6636
rect 18956 6972 19236 7028
rect 18844 6468 18900 6478
rect 18956 6468 19012 6972
rect 18844 6466 19012 6468
rect 18844 6414 18846 6466
rect 18898 6414 19012 6466
rect 18844 6412 19012 6414
rect 18844 6402 18900 6412
rect 18620 5236 18676 5246
rect 18508 5234 18676 5236
rect 18508 5182 18622 5234
rect 18674 5182 18676 5234
rect 18508 5180 18676 5182
rect 18620 5170 18676 5180
rect 18172 4398 18174 4450
rect 18226 4398 18228 4450
rect 18172 4386 18228 4398
rect 17500 4286 17502 4338
rect 17554 4286 17556 4338
rect 17500 4274 17556 4286
rect 18844 3666 18900 3678
rect 18844 3614 18846 3666
rect 18898 3614 18900 3666
rect 18844 800 18900 3614
rect 19404 3556 19460 9100
rect 19516 8484 19572 18844
rect 19628 18450 19684 19628
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18398 19630 18450
rect 19682 18398 19684 18450
rect 19628 17444 19684 18398
rect 19740 17444 19796 17454
rect 19628 17442 19796 17444
rect 19628 17390 19742 17442
rect 19794 17390 19796 17442
rect 19628 17388 19796 17390
rect 19628 16884 19684 17388
rect 19740 17378 19796 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 16884 20244 19852
rect 20300 19348 20356 19358
rect 20300 19234 20356 19292
rect 20300 19182 20302 19234
rect 20354 19182 20356 19234
rect 20300 19170 20356 19182
rect 20300 18452 20356 18462
rect 20300 18338 20356 18396
rect 20300 18286 20302 18338
rect 20354 18286 20356 18338
rect 20300 17332 20356 18286
rect 20412 18004 20468 24892
rect 20524 19684 20580 25228
rect 20636 25190 20692 25228
rect 20860 25284 20916 25294
rect 20860 25190 20916 25228
rect 20748 22708 20804 22718
rect 20748 22482 20804 22652
rect 20748 22430 20750 22482
rect 20802 22430 20804 22482
rect 20748 22418 20804 22430
rect 20524 19618 20580 19628
rect 20748 19348 20804 19358
rect 20748 19254 20804 19292
rect 20748 19124 20804 19134
rect 20636 19068 20748 19124
rect 20636 18674 20692 19068
rect 20748 19058 20804 19068
rect 20972 18676 21028 29596
rect 21196 29586 21252 29596
rect 21420 27188 21476 27198
rect 21308 27076 21364 27086
rect 21308 26982 21364 27020
rect 21420 26850 21476 27132
rect 21420 26798 21422 26850
rect 21474 26798 21476 26850
rect 21420 25844 21476 26798
rect 21420 25778 21476 25788
rect 21196 25508 21252 25518
rect 21252 25452 21364 25508
rect 21196 25442 21252 25452
rect 21308 25394 21364 25452
rect 21308 25342 21310 25394
rect 21362 25342 21364 25394
rect 21308 25330 21364 25342
rect 21420 25396 21476 25406
rect 21420 25302 21476 25340
rect 21420 22708 21476 22718
rect 21420 22370 21476 22652
rect 21420 22318 21422 22370
rect 21474 22318 21476 22370
rect 21420 22306 21476 22318
rect 21308 22260 21364 22270
rect 20636 18622 20638 18674
rect 20690 18622 20692 18674
rect 20636 18340 20692 18622
rect 20636 18274 20692 18284
rect 20860 18620 21028 18676
rect 21084 22258 21364 22260
rect 21084 22206 21310 22258
rect 21362 22206 21364 22258
rect 21084 22204 21364 22206
rect 20412 17938 20468 17948
rect 20300 17276 20692 17332
rect 20412 16884 20468 16894
rect 20188 16882 20468 16884
rect 20188 16830 20414 16882
rect 20466 16830 20468 16882
rect 20188 16828 20468 16830
rect 19628 16818 19684 16828
rect 19628 15874 19684 15886
rect 19628 15822 19630 15874
rect 19682 15822 19684 15874
rect 19628 14532 19684 15822
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15540 20244 15550
rect 20188 15446 20244 15484
rect 19628 14466 19684 14476
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19740 13186 19796 13198
rect 19740 13134 19742 13186
rect 19794 13134 19796 13186
rect 19740 13074 19796 13134
rect 19740 13022 19742 13074
rect 19794 13022 19796 13074
rect 19740 13010 19796 13022
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20412 12404 20468 16828
rect 20524 15426 20580 15438
rect 20524 15374 20526 15426
rect 20578 15374 20580 15426
rect 20524 14644 20580 15374
rect 20524 14578 20580 14588
rect 20636 13188 20692 17276
rect 20860 15540 20916 18620
rect 20972 18450 21028 18462
rect 20972 18398 20974 18450
rect 21026 18398 21028 18450
rect 20972 16996 21028 18398
rect 20972 16902 21028 16940
rect 20860 15474 20916 15484
rect 21084 15148 21140 22204
rect 21308 22194 21364 22204
rect 21532 22036 21588 33180
rect 21756 30210 21812 34524
rect 21756 30158 21758 30210
rect 21810 30158 21812 30210
rect 21756 29876 21812 30158
rect 21756 29810 21812 29820
rect 21868 29764 21924 34860
rect 21980 34804 22036 34974
rect 21980 34738 22036 34748
rect 22204 32452 22260 36316
rect 22428 35924 22484 37100
rect 22652 37044 22708 37054
rect 22540 36370 22596 36382
rect 22540 36318 22542 36370
rect 22594 36318 22596 36370
rect 22540 36148 22596 36318
rect 22652 36372 22708 36988
rect 22988 36596 23044 37998
rect 23660 37940 23716 37950
rect 22988 36530 23044 36540
rect 23212 37938 23716 37940
rect 23212 37886 23662 37938
rect 23714 37886 23716 37938
rect 23212 37884 23716 37886
rect 23212 36594 23268 37884
rect 23660 37874 23716 37884
rect 23212 36542 23214 36594
rect 23266 36542 23268 36594
rect 23212 36530 23268 36542
rect 23324 36484 23380 36494
rect 23324 36390 23380 36428
rect 23660 36484 23716 36494
rect 23884 36484 23940 36494
rect 23660 36390 23716 36428
rect 23772 36482 23940 36484
rect 23772 36430 23886 36482
rect 23938 36430 23940 36482
rect 23772 36428 23940 36430
rect 22652 36278 22708 36316
rect 22876 36372 22932 36382
rect 23100 36372 23156 36382
rect 22876 36370 23156 36372
rect 22876 36318 22878 36370
rect 22930 36318 23102 36370
rect 23154 36318 23156 36370
rect 22876 36316 23156 36318
rect 22876 36306 22932 36316
rect 23100 36306 23156 36316
rect 22596 36092 23268 36148
rect 22540 36054 22596 36092
rect 22540 35924 22596 35934
rect 22428 35922 22932 35924
rect 22428 35870 22542 35922
rect 22594 35870 22932 35922
rect 22428 35868 22932 35870
rect 22540 35858 22596 35868
rect 22428 35700 22484 35710
rect 22316 35698 22484 35700
rect 22316 35646 22430 35698
rect 22482 35646 22484 35698
rect 22316 35644 22484 35646
rect 22316 35140 22372 35644
rect 22428 35634 22484 35644
rect 22764 35700 22820 35710
rect 22764 35606 22820 35644
rect 22428 35476 22484 35486
rect 22428 35364 22484 35420
rect 22428 35308 22708 35364
rect 22316 34802 22372 35084
rect 22652 34914 22708 35308
rect 22652 34862 22654 34914
rect 22706 34862 22708 34914
rect 22652 34850 22708 34862
rect 22876 35028 22932 35868
rect 22988 35810 23044 36092
rect 22988 35758 22990 35810
rect 23042 35758 23044 35810
rect 22988 35746 23044 35758
rect 23100 35924 23156 35934
rect 23100 35810 23156 35868
rect 23100 35758 23102 35810
rect 23154 35758 23156 35810
rect 22988 35028 23044 35038
rect 22876 35026 23044 35028
rect 22876 34974 22990 35026
rect 23042 34974 23044 35026
rect 22876 34972 23044 34974
rect 22316 34750 22318 34802
rect 22370 34750 22372 34802
rect 22316 34244 22372 34750
rect 22428 34804 22484 34814
rect 22428 34710 22484 34748
rect 22316 34178 22372 34188
rect 22204 32386 22260 32396
rect 22092 31668 22148 31678
rect 22092 31574 22148 31612
rect 21980 30994 22036 31006
rect 21980 30942 21982 30994
rect 22034 30942 22036 30994
rect 21980 30884 22036 30942
rect 22204 30996 22260 31006
rect 22204 30902 22260 30940
rect 22652 30994 22708 31006
rect 22652 30942 22654 30994
rect 22706 30942 22708 30994
rect 21980 29986 22036 30828
rect 22428 30882 22484 30894
rect 22428 30830 22430 30882
rect 22482 30830 22484 30882
rect 22428 30212 22484 30830
rect 22428 30146 22484 30156
rect 22652 30210 22708 30942
rect 22652 30158 22654 30210
rect 22706 30158 22708 30210
rect 22652 30146 22708 30158
rect 22316 30100 22372 30110
rect 22316 30006 22372 30044
rect 22540 30100 22596 30110
rect 21980 29934 21982 29986
rect 22034 29934 22036 29986
rect 21980 29876 22036 29934
rect 22428 29988 22484 29998
rect 22540 29988 22596 30044
rect 22428 29986 22596 29988
rect 22428 29934 22430 29986
rect 22482 29934 22596 29986
rect 22428 29932 22596 29934
rect 21980 29820 22260 29876
rect 21868 29708 22148 29764
rect 21644 27858 21700 27870
rect 21644 27806 21646 27858
rect 21698 27806 21700 27858
rect 21644 27074 21700 27806
rect 21868 27858 21924 27870
rect 21868 27806 21870 27858
rect 21922 27806 21924 27858
rect 21756 27748 21812 27758
rect 21756 27654 21812 27692
rect 21644 27022 21646 27074
rect 21698 27022 21700 27074
rect 21644 27010 21700 27022
rect 21868 26908 21924 27806
rect 21980 27076 22036 27086
rect 21980 26982 22036 27020
rect 21644 26852 21924 26908
rect 22092 26908 22148 29708
rect 22204 27970 22260 29820
rect 22428 29540 22484 29932
rect 22428 29474 22484 29484
rect 22204 27918 22206 27970
rect 22258 27918 22260 27970
rect 22204 27860 22260 27918
rect 22316 27860 22372 27870
rect 22204 27804 22316 27860
rect 22316 27794 22372 27804
rect 22652 27748 22708 27758
rect 22652 27186 22708 27692
rect 22652 27134 22654 27186
rect 22706 27134 22708 27186
rect 22652 27122 22708 27134
rect 22876 26908 22932 34972
rect 22988 34962 23044 34972
rect 23100 35028 23156 35758
rect 23212 35700 23268 36092
rect 23772 36036 23828 36428
rect 23884 36418 23940 36428
rect 24444 36484 24500 36494
rect 24500 36428 24612 36484
rect 24444 36390 24500 36428
rect 24220 36372 24276 36382
rect 23324 35980 23828 36036
rect 23884 36260 23940 36270
rect 23324 35922 23380 35980
rect 23884 35924 23940 36204
rect 24220 36258 24276 36316
rect 24220 36206 24222 36258
rect 24274 36206 24276 36258
rect 24220 36194 24276 36206
rect 24332 36370 24388 36382
rect 24332 36318 24334 36370
rect 24386 36318 24388 36370
rect 23324 35870 23326 35922
rect 23378 35870 23380 35922
rect 23324 35858 23380 35870
rect 23660 35868 23940 35924
rect 24332 35924 24388 36318
rect 23660 35810 23716 35868
rect 24332 35858 24388 35868
rect 23660 35758 23662 35810
rect 23714 35758 23716 35810
rect 23660 35746 23716 35758
rect 24556 35812 24612 36428
rect 23548 35700 23604 35710
rect 23996 35700 24052 35710
rect 23212 35698 23604 35700
rect 23212 35646 23550 35698
rect 23602 35646 23604 35698
rect 23212 35644 23604 35646
rect 23100 34962 23156 34972
rect 23436 35028 23492 35038
rect 23436 34934 23492 34972
rect 23548 34916 23604 35644
rect 23772 35698 24052 35700
rect 23772 35646 23998 35698
rect 24050 35646 24052 35698
rect 23772 35644 24052 35646
rect 23660 35476 23716 35486
rect 23772 35476 23828 35644
rect 23996 35634 24052 35644
rect 24332 35700 24388 35710
rect 24556 35700 24612 35756
rect 24332 35606 24388 35644
rect 24444 35698 24612 35700
rect 24444 35646 24558 35698
rect 24610 35646 24612 35698
rect 24444 35644 24612 35646
rect 24220 35588 24276 35598
rect 24220 35494 24276 35532
rect 23660 35474 23828 35476
rect 23660 35422 23662 35474
rect 23714 35422 23828 35474
rect 23660 35420 23828 35422
rect 24108 35476 24164 35486
rect 23660 35410 23716 35420
rect 23772 34916 23828 34926
rect 23548 34914 23828 34916
rect 23548 34862 23774 34914
rect 23826 34862 23828 34914
rect 23548 34860 23828 34862
rect 23772 34850 23828 34860
rect 24108 34914 24164 35420
rect 24332 35364 24388 35374
rect 24108 34862 24110 34914
rect 24162 34862 24164 34914
rect 24108 34850 24164 34862
rect 24220 35308 24332 35364
rect 23884 34692 23940 34702
rect 23884 34598 23940 34636
rect 24108 34356 24164 34366
rect 24220 34356 24276 35308
rect 24332 35298 24388 35308
rect 24332 34804 24388 34814
rect 24444 34804 24500 35644
rect 24556 35634 24612 35644
rect 24332 34802 24500 34804
rect 24332 34750 24334 34802
rect 24386 34750 24500 34802
rect 24332 34748 24500 34750
rect 24556 34914 24612 34926
rect 24556 34862 24558 34914
rect 24610 34862 24612 34914
rect 24332 34738 24388 34748
rect 24556 34580 24612 34862
rect 24556 34514 24612 34524
rect 24108 34354 24276 34356
rect 24108 34302 24110 34354
rect 24162 34302 24276 34354
rect 24108 34300 24276 34302
rect 24108 34290 24164 34300
rect 23772 34244 23828 34254
rect 23772 34150 23828 34188
rect 23884 34242 23940 34254
rect 23884 34190 23886 34242
rect 23938 34190 23940 34242
rect 23884 34020 23940 34190
rect 23884 33954 23940 33964
rect 24444 34020 24500 34030
rect 24444 33926 24500 33964
rect 24444 33346 24500 33358
rect 24444 33294 24446 33346
rect 24498 33294 24500 33346
rect 24444 33124 24500 33294
rect 24668 33234 24724 38108
rect 24780 34692 24836 38612
rect 25004 36260 25060 36270
rect 25004 36166 25060 36204
rect 24780 34626 24836 34636
rect 24668 33182 24670 33234
rect 24722 33182 24724 33234
rect 24668 33170 24724 33182
rect 23548 31892 23604 31902
rect 23100 31220 23156 31230
rect 23100 31106 23156 31164
rect 23100 31054 23102 31106
rect 23154 31054 23156 31106
rect 23100 31042 23156 31054
rect 23212 30772 23268 30782
rect 23436 30772 23492 30782
rect 23212 30770 23492 30772
rect 23212 30718 23214 30770
rect 23266 30718 23438 30770
rect 23490 30718 23492 30770
rect 23212 30716 23492 30718
rect 23212 30706 23268 30716
rect 22988 30100 23044 30110
rect 22988 30006 23044 30044
rect 23324 27860 23380 27870
rect 22092 26852 22260 26908
rect 21644 25506 21700 26852
rect 21756 26180 21812 26190
rect 21756 26086 21812 26124
rect 21644 25454 21646 25506
rect 21698 25454 21700 25506
rect 21644 25442 21700 25454
rect 22092 25506 22148 25518
rect 22092 25454 22094 25506
rect 22146 25454 22148 25506
rect 22092 23492 22148 25454
rect 21868 23436 22092 23492
rect 21756 23380 21812 23390
rect 21756 22258 21812 23324
rect 21756 22206 21758 22258
rect 21810 22206 21812 22258
rect 21756 22194 21812 22206
rect 21196 21980 21588 22036
rect 21196 19012 21252 21980
rect 21532 20802 21588 20814
rect 21532 20750 21534 20802
rect 21586 20750 21588 20802
rect 21308 20580 21364 20590
rect 21308 20578 21476 20580
rect 21308 20526 21310 20578
rect 21362 20526 21476 20578
rect 21308 20524 21476 20526
rect 21308 20514 21364 20524
rect 21420 20130 21476 20524
rect 21420 20078 21422 20130
rect 21474 20078 21476 20130
rect 21420 20066 21476 20078
rect 21532 19234 21588 20750
rect 21644 20802 21700 20814
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21644 20132 21700 20750
rect 21868 20802 21924 23436
rect 22092 23426 22148 23436
rect 22204 22596 22260 26852
rect 22428 26852 22932 26908
rect 22988 27076 23044 27086
rect 22316 26068 22372 26078
rect 22316 25730 22372 26012
rect 22316 25678 22318 25730
rect 22370 25678 22372 25730
rect 22316 25666 22372 25678
rect 22204 22530 22260 22540
rect 21868 20750 21870 20802
rect 21922 20750 21924 20802
rect 21868 20738 21924 20750
rect 22092 20692 22148 20702
rect 22092 20598 22148 20636
rect 21644 20066 21700 20076
rect 22204 20018 22260 20030
rect 22204 19966 22206 20018
rect 22258 19966 22260 20018
rect 21980 19572 22036 19582
rect 21756 19460 21812 19470
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 21532 19124 21588 19182
rect 21532 19058 21588 19068
rect 21644 19458 21812 19460
rect 21644 19406 21758 19458
rect 21810 19406 21812 19458
rect 21644 19404 21812 19406
rect 21196 18946 21252 18956
rect 21532 18676 21588 18686
rect 21644 18676 21700 19404
rect 21756 19394 21812 19404
rect 21532 18674 21700 18676
rect 21532 18622 21534 18674
rect 21586 18622 21700 18674
rect 21532 18620 21700 18622
rect 21868 19010 21924 19022
rect 21868 18958 21870 19010
rect 21922 18958 21924 19010
rect 21532 18610 21588 18620
rect 21420 18562 21476 18574
rect 21420 18510 21422 18562
rect 21474 18510 21476 18562
rect 21196 18452 21252 18462
rect 21420 18452 21476 18510
rect 21252 18396 21476 18452
rect 21868 18452 21924 18958
rect 21196 18386 21252 18396
rect 21868 18386 21924 18396
rect 21980 18674 22036 19516
rect 22204 19348 22260 19966
rect 22092 19124 22148 19134
rect 22092 19030 22148 19068
rect 21980 18622 21982 18674
rect 22034 18622 22036 18674
rect 21644 18228 21700 18238
rect 21980 18228 22036 18622
rect 21644 18226 22036 18228
rect 21644 18174 21646 18226
rect 21698 18174 22036 18226
rect 21644 18172 22036 18174
rect 21644 18162 21700 18172
rect 21644 18004 21700 18014
rect 21644 16884 21700 17948
rect 21868 17780 21924 17790
rect 22204 17780 22260 19292
rect 22316 19460 22372 19470
rect 22316 19234 22372 19404
rect 22428 19348 22484 26852
rect 22988 26516 23044 27020
rect 22540 26460 23156 26516
rect 22540 26290 22596 26460
rect 22540 26238 22542 26290
rect 22594 26238 22596 26290
rect 22540 26226 22596 26238
rect 22764 26292 22820 26302
rect 22764 26198 22820 26236
rect 22988 26180 23044 26190
rect 22988 26086 23044 26124
rect 23100 25618 23156 26460
rect 23100 25566 23102 25618
rect 23154 25566 23156 25618
rect 23100 25554 23156 25566
rect 23212 26290 23268 26302
rect 23212 26238 23214 26290
rect 23266 26238 23268 26290
rect 22652 25508 22708 25518
rect 22652 25414 22708 25452
rect 23212 25284 23268 26238
rect 23324 26290 23380 27804
rect 23324 26238 23326 26290
rect 23378 26238 23380 26290
rect 23324 26226 23380 26238
rect 23436 26068 23492 30716
rect 23548 30210 23604 31836
rect 24220 31890 24276 31902
rect 24220 31838 24222 31890
rect 24274 31838 24276 31890
rect 24220 31780 24276 31838
rect 24220 31714 24276 31724
rect 24108 31444 24164 31454
rect 23660 31220 23716 31230
rect 23660 31126 23716 31164
rect 23548 30158 23550 30210
rect 23602 30158 23604 30210
rect 23548 30146 23604 30158
rect 23212 25218 23268 25228
rect 23324 26012 23492 26068
rect 23996 28756 24052 28766
rect 23324 24948 23380 26012
rect 22876 24892 23380 24948
rect 23436 25284 23492 25294
rect 23436 24946 23492 25228
rect 23996 25172 24052 28700
rect 23996 25106 24052 25116
rect 23436 24894 23438 24946
rect 23490 24894 23492 24946
rect 22764 22370 22820 22382
rect 22764 22318 22766 22370
rect 22818 22318 22820 22370
rect 22764 22148 22820 22318
rect 22764 22082 22820 22092
rect 22428 19282 22484 19292
rect 22652 20692 22708 20702
rect 22652 19460 22708 20636
rect 22316 19182 22318 19234
rect 22370 19182 22372 19234
rect 22316 19170 22372 19182
rect 22652 19234 22708 19404
rect 22652 19182 22654 19234
rect 22706 19182 22708 19234
rect 22652 19170 22708 19182
rect 22764 19908 22820 19918
rect 22316 18900 22372 18910
rect 22316 18674 22372 18844
rect 22316 18622 22318 18674
rect 22370 18622 22372 18674
rect 22316 18610 22372 18622
rect 22764 18676 22820 19852
rect 22764 18610 22820 18620
rect 22876 19348 22932 24892
rect 23324 24724 23380 24734
rect 23324 24630 23380 24668
rect 22988 23380 23044 23390
rect 22988 20802 23044 23324
rect 23436 23380 23492 24894
rect 23884 25060 23940 25070
rect 23884 24946 23940 25004
rect 23884 24894 23886 24946
rect 23938 24894 23940 24946
rect 23884 24724 23940 24894
rect 23884 24658 23940 24668
rect 23436 23314 23492 23324
rect 23548 24612 23604 24622
rect 23548 23268 23604 24556
rect 23548 23202 23604 23212
rect 23436 22258 23492 22270
rect 23436 22206 23438 22258
rect 23490 22206 23492 22258
rect 23324 20916 23380 20926
rect 22988 20750 22990 20802
rect 23042 20750 23044 20802
rect 22988 20738 23044 20750
rect 23100 20804 23156 20814
rect 23100 20710 23156 20748
rect 23324 20802 23380 20860
rect 23324 20750 23326 20802
rect 23378 20750 23380 20802
rect 23324 20356 23380 20750
rect 23436 20578 23492 22206
rect 24108 21028 24164 31388
rect 24444 31444 24500 33068
rect 24668 32452 24724 32462
rect 24668 32358 24724 32396
rect 25116 31948 25172 38668
rect 25452 38610 25508 38622
rect 25452 38558 25454 38610
rect 25506 38558 25508 38610
rect 25452 38164 25508 38558
rect 25788 38164 25844 38174
rect 25452 38162 25844 38164
rect 25452 38110 25790 38162
rect 25842 38110 25844 38162
rect 25452 38108 25844 38110
rect 25788 37044 25844 38108
rect 26012 37828 26068 39566
rect 26572 39396 26628 39406
rect 26572 39302 26628 39340
rect 26684 39058 26740 39676
rect 27244 39620 27300 39630
rect 27244 39618 27412 39620
rect 27244 39566 27246 39618
rect 27298 39566 27412 39618
rect 27244 39564 27412 39566
rect 27244 39554 27300 39564
rect 26684 39006 26686 39058
rect 26738 39006 26740 39058
rect 26684 38994 26740 39006
rect 27356 39060 27412 39564
rect 27468 39506 27524 41132
rect 28364 41188 28420 41198
rect 28364 41094 28420 41132
rect 28252 40404 28308 40414
rect 27916 40402 28308 40404
rect 27916 40350 28254 40402
rect 28306 40350 28308 40402
rect 27916 40348 28308 40350
rect 27468 39454 27470 39506
rect 27522 39454 27524 39506
rect 27468 39442 27524 39454
rect 27804 39508 27860 39518
rect 27804 39414 27860 39452
rect 27356 39004 27860 39060
rect 27580 38836 27636 38846
rect 27356 38834 27636 38836
rect 27356 38782 27582 38834
rect 27634 38782 27636 38834
rect 27356 38780 27636 38782
rect 26236 38724 26292 38734
rect 26236 38630 26292 38668
rect 26236 37828 26292 37838
rect 26012 37826 26292 37828
rect 26012 37774 26238 37826
rect 26290 37774 26292 37826
rect 26012 37772 26292 37774
rect 25788 36978 25844 36988
rect 25676 36596 25732 36606
rect 25676 36484 25732 36540
rect 25564 36482 25732 36484
rect 25564 36430 25678 36482
rect 25730 36430 25732 36482
rect 25564 36428 25732 36430
rect 25228 35812 25284 35822
rect 25228 35718 25284 35756
rect 25452 35700 25508 35710
rect 25340 35698 25508 35700
rect 25340 35646 25454 35698
rect 25506 35646 25508 35698
rect 25340 35644 25508 35646
rect 25340 35364 25396 35644
rect 25452 35634 25508 35644
rect 25340 35298 25396 35308
rect 25564 35364 25620 36428
rect 25676 36418 25732 36428
rect 25788 35698 25844 35710
rect 25788 35646 25790 35698
rect 25842 35646 25844 35698
rect 25564 34914 25620 35308
rect 25676 35586 25732 35598
rect 25676 35534 25678 35586
rect 25730 35534 25732 35586
rect 25676 35140 25732 35534
rect 25788 35476 25844 35646
rect 25788 35410 25844 35420
rect 26236 35252 26292 37772
rect 26572 37044 26628 37054
rect 26460 36372 26516 36382
rect 26460 36278 26516 36316
rect 26236 35196 26516 35252
rect 25676 35084 26404 35140
rect 26348 35026 26404 35084
rect 26348 34974 26350 35026
rect 26402 34974 26404 35026
rect 26348 34962 26404 34974
rect 25564 34862 25566 34914
rect 25618 34862 25620 34914
rect 25564 34850 25620 34862
rect 25564 34692 25620 34702
rect 25564 33570 25620 34636
rect 26460 34468 26516 35196
rect 25564 33518 25566 33570
rect 25618 33518 25620 33570
rect 25564 33506 25620 33518
rect 25900 34412 26516 34468
rect 25228 33348 25284 33358
rect 25228 33254 25284 33292
rect 25004 31892 25172 31948
rect 24444 31378 24500 31388
rect 24556 31778 24612 31790
rect 24556 31726 24558 31778
rect 24610 31726 24612 31778
rect 24220 30884 24276 30894
rect 24556 30884 24612 31726
rect 24780 31780 24836 31790
rect 24780 31686 24836 31724
rect 24220 30882 24612 30884
rect 24220 30830 24222 30882
rect 24274 30830 24612 30882
rect 24220 30828 24612 30830
rect 25004 31220 25060 31892
rect 25116 31780 25172 31790
rect 25116 31686 25172 31724
rect 24220 30770 24276 30828
rect 24220 30718 24222 30770
rect 24274 30718 24276 30770
rect 24220 30706 24276 30718
rect 24332 30212 24388 30222
rect 24332 30118 24388 30156
rect 24780 27188 24836 27198
rect 24780 27094 24836 27132
rect 25004 26908 25060 31164
rect 25340 29876 25396 29886
rect 25340 28530 25396 29820
rect 25564 28756 25620 28766
rect 25564 28642 25620 28700
rect 25564 28590 25566 28642
rect 25618 28590 25620 28642
rect 25564 28578 25620 28590
rect 25340 28478 25342 28530
rect 25394 28478 25396 28530
rect 25340 28466 25396 28478
rect 25676 27412 25732 27422
rect 25452 27188 25508 27198
rect 25228 27076 25284 27086
rect 25228 26982 25284 27020
rect 25004 26852 25172 26908
rect 24892 24500 24948 24510
rect 24892 21700 24948 24444
rect 24332 21588 24388 21598
rect 24332 21494 24388 21532
rect 23996 20972 24164 21028
rect 24220 21364 24276 21374
rect 23772 20692 23828 20702
rect 23772 20598 23828 20636
rect 23436 20526 23438 20578
rect 23490 20526 23492 20578
rect 23436 20514 23492 20526
rect 23324 20300 23492 20356
rect 22988 20132 23044 20142
rect 22988 19796 23044 20076
rect 23100 20020 23156 20030
rect 23436 20020 23492 20300
rect 23100 19926 23156 19964
rect 23324 19964 23492 20020
rect 23548 20132 23604 20142
rect 23100 19796 23156 19806
rect 22988 19794 23156 19796
rect 22988 19742 23102 19794
rect 23154 19742 23156 19794
rect 22988 19740 23156 19742
rect 23100 19730 23156 19740
rect 23100 19460 23156 19470
rect 23100 19366 23156 19404
rect 22876 19234 22932 19292
rect 23324 19236 23380 19964
rect 23436 19794 23492 19806
rect 23436 19742 23438 19794
rect 23490 19742 23492 19794
rect 23436 19572 23492 19742
rect 23436 19506 23492 19516
rect 22876 19182 22878 19234
rect 22930 19182 22932 19234
rect 22764 18450 22820 18462
rect 22764 18398 22766 18450
rect 22818 18398 22820 18450
rect 22316 17780 22372 17790
rect 21924 17724 22148 17780
rect 22204 17724 22316 17780
rect 21868 17686 21924 17724
rect 22092 17108 22148 17724
rect 22316 17666 22372 17724
rect 22316 17614 22318 17666
rect 22370 17614 22372 17666
rect 22316 17602 22372 17614
rect 22204 17108 22260 17118
rect 22092 17052 22204 17108
rect 22204 17014 22260 17052
rect 21868 16996 21924 17006
rect 21644 16882 21812 16884
rect 21644 16830 21646 16882
rect 21698 16830 21812 16882
rect 21644 16828 21812 16830
rect 21644 16818 21700 16828
rect 21756 16548 21812 16828
rect 21868 16660 21924 16940
rect 22764 16996 22820 18398
rect 22764 16930 22820 16940
rect 22652 16884 22708 16894
rect 22652 16772 22708 16828
rect 22876 16772 22932 19182
rect 23100 19234 23380 19236
rect 23100 19182 23326 19234
rect 23378 19182 23380 19234
rect 23100 19180 23380 19182
rect 22988 19010 23044 19022
rect 22988 18958 22990 19010
rect 23042 18958 23044 19010
rect 22988 17778 23044 18958
rect 23100 18674 23156 19180
rect 23324 19170 23380 19180
rect 23100 18622 23102 18674
rect 23154 18622 23156 18674
rect 23100 18610 23156 18622
rect 23324 18676 23380 18686
rect 22988 17726 22990 17778
rect 23042 17726 23044 17778
rect 22988 17714 23044 17726
rect 22428 16770 22708 16772
rect 22428 16718 22654 16770
rect 22706 16718 22708 16770
rect 22428 16716 22708 16718
rect 21868 16604 22260 16660
rect 21756 16492 22148 16548
rect 21532 15540 21588 15550
rect 21588 15484 21812 15540
rect 21532 15446 21588 15484
rect 20972 15092 21140 15148
rect 21644 15314 21700 15326
rect 21644 15262 21646 15314
rect 21698 15262 21700 15314
rect 20748 13188 20804 13198
rect 20636 13132 20748 13188
rect 20748 13074 20804 13132
rect 20748 13022 20750 13074
rect 20802 13022 20804 13074
rect 20748 13010 20804 13022
rect 20412 12338 20468 12348
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19740 10724 19796 10734
rect 19740 10630 19796 10668
rect 20524 10724 20580 10734
rect 20300 10498 20356 10510
rect 20300 10446 20302 10498
rect 20354 10446 20356 10498
rect 20300 10386 20356 10446
rect 20300 10334 20302 10386
rect 20354 10334 20356 10386
rect 19740 9604 19796 9642
rect 19740 9538 19796 9548
rect 20188 9604 20244 9614
rect 20300 9604 20356 10334
rect 20188 9602 20356 9604
rect 20188 9550 20190 9602
rect 20242 9550 20356 9602
rect 20188 9548 20356 9550
rect 20524 9826 20580 10668
rect 20748 10500 20804 10510
rect 20748 10406 20804 10444
rect 20524 9774 20526 9826
rect 20578 9774 20580 9826
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 8484 20244 9548
rect 19572 8428 19684 8484
rect 19516 8418 19572 8428
rect 19516 8036 19572 8046
rect 19516 7252 19572 7980
rect 19628 7364 19684 8428
rect 20076 8428 20244 8484
rect 19852 8372 19908 8382
rect 19852 8258 19908 8316
rect 19852 8206 19854 8258
rect 19906 8206 19908 8258
rect 19852 8194 19908 8206
rect 19964 8260 20020 8270
rect 20076 8260 20132 8428
rect 20524 8372 20580 9774
rect 20972 9716 21028 15092
rect 21532 15090 21588 15102
rect 21532 15038 21534 15090
rect 21586 15038 21588 15090
rect 21196 14532 21252 14542
rect 21196 14438 21252 14476
rect 21532 14530 21588 15038
rect 21532 14478 21534 14530
rect 21586 14478 21588 14530
rect 21532 14466 21588 14478
rect 21644 14532 21700 15262
rect 21644 14466 21700 14476
rect 21420 14306 21476 14318
rect 21420 14254 21422 14306
rect 21474 14254 21476 14306
rect 21308 13860 21364 13870
rect 21420 13860 21476 14254
rect 21308 13858 21476 13860
rect 21308 13806 21310 13858
rect 21362 13806 21476 13858
rect 21308 13804 21476 13806
rect 21308 13794 21364 13804
rect 21308 13188 21364 13198
rect 21308 12962 21364 13132
rect 21308 12910 21310 12962
rect 21362 12910 21364 12962
rect 21308 12898 21364 12910
rect 21756 13074 21812 15484
rect 21868 14418 21924 14430
rect 21868 14366 21870 14418
rect 21922 14366 21924 14418
rect 21868 14196 21924 14366
rect 21868 14130 21924 14140
rect 21756 13022 21758 13074
rect 21810 13022 21812 13074
rect 21756 12292 21812 13022
rect 21756 12226 21812 12236
rect 20972 9650 21028 9660
rect 21196 10948 21252 10958
rect 21196 10498 21252 10892
rect 21644 10722 21700 10734
rect 21644 10670 21646 10722
rect 21698 10670 21700 10722
rect 21196 10446 21198 10498
rect 21250 10446 21252 10498
rect 20636 9604 20692 9614
rect 20636 9510 20692 9548
rect 20860 9602 20916 9614
rect 20860 9550 20862 9602
rect 20914 9550 20916 9602
rect 20748 9492 20804 9502
rect 20748 9044 20804 9436
rect 20860 9380 20916 9550
rect 21196 9492 21252 10446
rect 21532 10610 21588 10622
rect 21532 10558 21534 10610
rect 21586 10558 21588 10610
rect 21308 10388 21364 10398
rect 21532 10388 21588 10558
rect 21644 10500 21700 10670
rect 21868 10612 21924 10622
rect 21868 10518 21924 10556
rect 21644 10434 21700 10444
rect 21308 10386 21588 10388
rect 21308 10334 21310 10386
rect 21362 10334 21588 10386
rect 21308 10332 21588 10334
rect 21308 10322 21364 10332
rect 21196 9426 21252 9436
rect 21420 9716 21476 9726
rect 20860 9314 20916 9324
rect 21308 9380 21364 9390
rect 21196 9044 21252 9054
rect 20748 8988 20916 9044
rect 20748 8708 20804 8988
rect 20748 8642 20804 8652
rect 20524 8306 20580 8316
rect 20020 8204 20132 8260
rect 20188 8260 20244 8270
rect 19964 8194 20020 8204
rect 20188 8166 20244 8204
rect 20412 8146 20468 8158
rect 20412 8094 20414 8146
rect 20466 8094 20468 8146
rect 19964 8036 20020 8074
rect 19964 7970 20020 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20300 7700 20356 7710
rect 20412 7700 20468 8094
rect 20748 8148 20804 8158
rect 20748 8054 20804 8092
rect 20356 7644 20468 7700
rect 20300 7606 20356 7644
rect 19964 7588 20020 7598
rect 19964 7494 20020 7532
rect 20636 7588 20692 7598
rect 20636 7494 20692 7532
rect 19628 7308 20020 7364
rect 19516 6804 19572 7196
rect 19628 6804 19684 6814
rect 19516 6802 19684 6804
rect 19516 6750 19630 6802
rect 19682 6750 19684 6802
rect 19516 6748 19684 6750
rect 19628 6738 19684 6748
rect 19964 6804 20020 7308
rect 19964 6802 20356 6804
rect 19964 6750 19966 6802
rect 20018 6750 20356 6802
rect 19964 6748 20356 6750
rect 19964 6738 20020 6748
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20300 4226 20356 6748
rect 20748 5236 20804 5246
rect 20860 5236 20916 8988
rect 20972 8708 21028 8718
rect 20972 5684 21028 8652
rect 21196 7700 21252 8988
rect 21308 8258 21364 9324
rect 21420 8932 21476 9660
rect 21532 9604 21588 10332
rect 21980 10276 22036 16492
rect 22092 16210 22148 16492
rect 22092 16158 22094 16210
rect 22146 16158 22148 16210
rect 22092 16146 22148 16158
rect 22092 15426 22148 15438
rect 22092 15374 22094 15426
rect 22146 15374 22148 15426
rect 22092 14196 22148 15374
rect 22204 15316 22260 16604
rect 22316 15316 22372 15326
rect 22204 15314 22372 15316
rect 22204 15262 22318 15314
rect 22370 15262 22372 15314
rect 22204 15260 22372 15262
rect 22316 15250 22372 15260
rect 22092 14130 22148 14140
rect 22092 13748 22148 13758
rect 22092 13654 22148 13692
rect 22428 13524 22484 16716
rect 22652 16706 22708 16716
rect 22764 16716 22932 16772
rect 22652 14868 22708 14878
rect 22540 14532 22596 14542
rect 22540 14438 22596 14476
rect 22652 14308 22708 14812
rect 22540 14306 22708 14308
rect 22540 14254 22654 14306
rect 22706 14254 22708 14306
rect 22540 14252 22708 14254
rect 22540 13860 22596 14252
rect 22652 14242 22708 14252
rect 22540 13766 22596 13804
rect 22092 13468 22484 13524
rect 22652 13748 22708 13758
rect 22092 11172 22148 13468
rect 22652 12962 22708 13692
rect 22652 12910 22654 12962
rect 22706 12910 22708 12962
rect 22652 12898 22708 12910
rect 22764 12068 22820 16716
rect 22876 15540 22932 15550
rect 22876 15446 22932 15484
rect 23324 14868 23380 18620
rect 23548 18564 23604 20076
rect 23884 20130 23940 20142
rect 23884 20078 23886 20130
rect 23938 20078 23940 20130
rect 23884 19908 23940 20078
rect 23884 19842 23940 19852
rect 23772 19794 23828 19806
rect 23772 19742 23774 19794
rect 23826 19742 23828 19794
rect 23772 19460 23828 19742
rect 23772 19394 23828 19404
rect 23884 19236 23940 19246
rect 23884 19142 23940 19180
rect 23772 19124 23828 19134
rect 23772 19030 23828 19068
rect 23548 18450 23604 18508
rect 23548 18398 23550 18450
rect 23602 18398 23604 18450
rect 23548 18386 23604 18398
rect 23996 15148 24052 20972
rect 24108 20804 24164 20814
rect 24220 20804 24276 21308
rect 24108 20802 24276 20804
rect 24108 20750 24110 20802
rect 24162 20750 24276 20802
rect 24108 20748 24276 20750
rect 24556 20804 24612 20814
rect 24108 20738 24164 20748
rect 24556 20710 24612 20748
rect 24444 20692 24500 20702
rect 24220 20690 24500 20692
rect 24220 20638 24446 20690
rect 24498 20638 24500 20690
rect 24220 20636 24500 20638
rect 24108 20132 24164 20142
rect 24220 20132 24276 20636
rect 24444 20626 24500 20636
rect 24108 20130 24276 20132
rect 24108 20078 24110 20130
rect 24162 20078 24276 20130
rect 24108 20076 24276 20078
rect 24668 20578 24724 20590
rect 24668 20526 24670 20578
rect 24722 20526 24724 20578
rect 24108 19572 24164 20076
rect 24556 19908 24612 19918
rect 24668 19908 24724 20526
rect 24556 19906 24724 19908
rect 24556 19854 24558 19906
rect 24610 19854 24724 19906
rect 24556 19852 24724 19854
rect 24556 19684 24612 19852
rect 24556 19618 24612 19628
rect 24108 19506 24164 19516
rect 24332 19348 24388 19358
rect 24332 19254 24388 19292
rect 24780 19236 24836 19246
rect 24780 19142 24836 19180
rect 24892 15148 24948 21644
rect 25116 17778 25172 26852
rect 25452 26290 25508 27132
rect 25676 27186 25732 27356
rect 25676 27134 25678 27186
rect 25730 27134 25732 27186
rect 25676 27122 25732 27134
rect 25452 26238 25454 26290
rect 25506 26238 25508 26290
rect 25452 26226 25508 26238
rect 25564 26852 25620 26862
rect 25228 26178 25284 26190
rect 25228 26126 25230 26178
rect 25282 26126 25284 26178
rect 25228 25284 25284 26126
rect 25228 25218 25284 25228
rect 25564 25396 25620 26796
rect 25788 26516 25844 26526
rect 25788 26422 25844 26460
rect 25452 25060 25508 25070
rect 25452 22484 25508 25004
rect 25564 24610 25620 25340
rect 25900 25060 25956 34412
rect 26348 34020 26404 34030
rect 26124 33124 26180 33134
rect 26124 33030 26180 33068
rect 26236 29428 26292 29438
rect 26236 29334 26292 29372
rect 26348 28868 26404 33964
rect 26572 33572 26628 36988
rect 26908 34916 26964 34926
rect 26908 34356 26964 34860
rect 26908 34262 26964 34300
rect 26460 33516 26628 33572
rect 27356 33570 27412 38780
rect 27580 38770 27636 38780
rect 27804 36820 27860 39004
rect 27916 39058 27972 40348
rect 28252 40338 28308 40348
rect 28364 40404 28420 40414
rect 28140 39508 28196 39518
rect 28364 39508 28420 40348
rect 28476 39844 28532 44200
rect 29372 41412 29428 41422
rect 29372 41318 29428 41356
rect 29596 41412 29652 44200
rect 29596 41346 29652 41356
rect 29708 40852 29764 40862
rect 29260 40628 29316 40638
rect 29260 40534 29316 40572
rect 29484 40068 29540 40078
rect 28476 39778 28532 39788
rect 29372 39844 29428 39854
rect 29372 39750 29428 39788
rect 28140 39506 28420 39508
rect 28140 39454 28142 39506
rect 28194 39454 28420 39506
rect 28140 39452 28420 39454
rect 28140 39442 28196 39452
rect 27916 39006 27918 39058
rect 27970 39006 27972 39058
rect 27916 38994 27972 39006
rect 28700 39394 28756 39406
rect 28700 39342 28702 39394
rect 28754 39342 28756 39394
rect 28700 39060 28756 39342
rect 28700 39004 29092 39060
rect 29036 38948 29092 39004
rect 29148 38948 29204 38958
rect 29036 38946 29204 38948
rect 29036 38894 29150 38946
rect 29202 38894 29204 38946
rect 29036 38892 29204 38894
rect 28924 38834 28980 38846
rect 28924 38782 28926 38834
rect 28978 38782 28980 38834
rect 28364 38724 28420 38734
rect 28924 38724 28980 38782
rect 28364 38722 28980 38724
rect 28364 38670 28366 38722
rect 28418 38670 28980 38722
rect 28364 38668 28980 38670
rect 27804 36764 28308 36820
rect 27356 33518 27358 33570
rect 27410 33518 27412 33570
rect 26460 30322 26516 33516
rect 27356 33506 27412 33518
rect 27916 34356 27972 34366
rect 26572 33348 26628 33358
rect 26572 33254 26628 33292
rect 27692 33346 27748 33358
rect 27692 33294 27694 33346
rect 27746 33294 27748 33346
rect 27692 32900 27748 33294
rect 27916 33236 27972 34300
rect 28252 34354 28308 36764
rect 28252 34302 28254 34354
rect 28306 34302 28308 34354
rect 28252 34290 28308 34302
rect 28364 34132 28420 38668
rect 28700 37940 28756 37950
rect 28700 37846 28756 37884
rect 28700 37492 28756 37502
rect 28588 36594 28644 36606
rect 28588 36542 28590 36594
rect 28642 36542 28644 36594
rect 28588 35924 28644 36542
rect 28588 35858 28644 35868
rect 27692 32834 27748 32844
rect 27804 33234 27972 33236
rect 27804 33182 27918 33234
rect 27970 33182 27972 33234
rect 27804 33180 27972 33182
rect 26684 32562 26740 32574
rect 26684 32510 26686 32562
rect 26738 32510 26740 32562
rect 26684 32452 26740 32510
rect 26684 31948 26740 32396
rect 27244 32450 27300 32462
rect 27244 32398 27246 32450
rect 27298 32398 27300 32450
rect 26684 31892 27076 31948
rect 26460 30270 26462 30322
rect 26514 30270 26516 30322
rect 26460 30212 26516 30270
rect 26460 30146 26516 30156
rect 26572 30100 26628 30110
rect 26572 29650 26628 30044
rect 26796 29986 26852 29998
rect 26796 29934 26798 29986
rect 26850 29934 26852 29986
rect 26796 29876 26852 29934
rect 26796 29810 26852 29820
rect 26572 29598 26574 29650
rect 26626 29598 26628 29650
rect 26572 29586 26628 29598
rect 26572 28868 26628 28878
rect 26348 28812 26572 28868
rect 26012 28644 26068 28654
rect 26012 28550 26068 28588
rect 26348 28644 26404 28654
rect 26348 28530 26404 28588
rect 26348 28478 26350 28530
rect 26402 28478 26404 28530
rect 26348 28466 26404 28478
rect 25900 24994 25956 25004
rect 25564 24558 25566 24610
rect 25618 24558 25620 24610
rect 25564 24546 25620 24558
rect 25564 22484 25620 22494
rect 25452 22482 25620 22484
rect 25452 22430 25566 22482
rect 25618 22430 25620 22482
rect 25452 22428 25620 22430
rect 25564 22418 25620 22428
rect 25900 22260 25956 22270
rect 25452 22148 25508 22158
rect 25340 21700 25396 21710
rect 25340 21588 25396 21644
rect 25228 21586 25396 21588
rect 25228 21534 25342 21586
rect 25394 21534 25396 21586
rect 25228 21532 25396 21534
rect 25228 20914 25284 21532
rect 25340 21522 25396 21532
rect 25228 20862 25230 20914
rect 25282 20862 25284 20914
rect 25228 20850 25284 20862
rect 25116 17726 25118 17778
rect 25170 17726 25172 17778
rect 25116 17556 25172 17726
rect 25340 19908 25396 19918
rect 25452 19908 25508 22092
rect 25900 21698 25956 22204
rect 26012 22148 26068 22158
rect 26012 22054 26068 22092
rect 25900 21646 25902 21698
rect 25954 21646 25956 21698
rect 25900 21634 25956 21646
rect 25676 21588 25732 21598
rect 25676 20914 25732 21532
rect 25676 20862 25678 20914
rect 25730 20862 25732 20914
rect 25676 20580 25732 20862
rect 25676 20514 25732 20524
rect 25788 21362 25844 21374
rect 25788 21310 25790 21362
rect 25842 21310 25844 21362
rect 25340 19906 25508 19908
rect 25340 19854 25342 19906
rect 25394 19854 25508 19906
rect 25340 19852 25508 19854
rect 25340 18450 25396 19852
rect 25340 18398 25342 18450
rect 25394 18398 25396 18450
rect 25340 17780 25396 18398
rect 25564 17780 25620 17790
rect 25340 17724 25564 17780
rect 25564 17686 25620 17724
rect 25116 17490 25172 17500
rect 25676 15426 25732 15438
rect 25676 15374 25678 15426
rect 25730 15374 25732 15426
rect 25564 15316 25620 15326
rect 23996 15092 24164 15148
rect 23324 14802 23380 14812
rect 24108 14868 24164 15092
rect 24780 15092 24948 15148
rect 25340 15202 25396 15214
rect 25340 15150 25342 15202
rect 25394 15150 25396 15202
rect 24108 14812 24724 14868
rect 22988 14588 23380 14644
rect 22876 14532 22932 14542
rect 22988 14532 23044 14588
rect 22876 14530 23044 14532
rect 22876 14478 22878 14530
rect 22930 14478 23044 14530
rect 22876 14476 23044 14478
rect 23324 14530 23380 14588
rect 23324 14478 23326 14530
rect 23378 14478 23380 14530
rect 22876 14466 22932 14476
rect 23324 14466 23380 14478
rect 23100 14418 23156 14430
rect 23100 14366 23102 14418
rect 23154 14366 23156 14418
rect 22092 11106 22148 11116
rect 22204 12012 22820 12068
rect 22876 14308 22932 14318
rect 22092 10948 22148 10958
rect 22092 10722 22148 10892
rect 22204 10836 22260 12012
rect 22876 11396 22932 14252
rect 23100 14196 23156 14366
rect 23660 14420 23716 14430
rect 23884 14420 23940 14430
rect 23660 14418 23940 14420
rect 23660 14366 23662 14418
rect 23714 14366 23886 14418
rect 23938 14366 23940 14418
rect 23660 14364 23940 14366
rect 23660 14354 23716 14364
rect 23884 14354 23940 14364
rect 23436 14306 23492 14318
rect 23436 14254 23438 14306
rect 23490 14254 23492 14306
rect 23212 14196 23268 14206
rect 23100 14140 23212 14196
rect 23212 14130 23268 14140
rect 23324 13076 23380 13086
rect 23436 13076 23492 14254
rect 24108 14306 24164 14812
rect 24108 14254 24110 14306
rect 24162 14254 24164 14306
rect 24108 13300 24164 14254
rect 24220 14644 24276 14654
rect 24220 14530 24276 14588
rect 24668 14642 24724 14812
rect 24668 14590 24670 14642
rect 24722 14590 24724 14642
rect 24668 14578 24724 14590
rect 24220 14478 24222 14530
rect 24274 14478 24276 14530
rect 24220 14084 24276 14478
rect 24220 14018 24276 14028
rect 24108 13234 24164 13244
rect 23324 13074 23492 13076
rect 23324 13022 23326 13074
rect 23378 13022 23492 13074
rect 23324 13020 23492 13022
rect 23324 13010 23380 13020
rect 22428 11340 22932 11396
rect 22204 10742 22260 10780
rect 22316 11282 22372 11294
rect 22316 11230 22318 11282
rect 22370 11230 22372 11282
rect 22092 10670 22094 10722
rect 22146 10670 22148 10722
rect 22092 10658 22148 10670
rect 22316 10724 22372 11230
rect 22428 11282 22484 11340
rect 22428 11230 22430 11282
rect 22482 11230 22484 11282
rect 22428 11218 22484 11230
rect 22876 11284 22932 11340
rect 24108 12404 24164 12414
rect 22988 11284 23044 11294
rect 22876 11282 23268 11284
rect 22876 11230 22990 11282
rect 23042 11230 23268 11282
rect 22876 11228 23268 11230
rect 22988 11218 23044 11228
rect 22652 11172 22708 11182
rect 22652 11170 22820 11172
rect 22652 11118 22654 11170
rect 22706 11118 22820 11170
rect 22652 11116 22820 11118
rect 22652 11106 22708 11116
rect 22316 10658 22372 10668
rect 22204 10388 22260 10398
rect 21980 10210 22036 10220
rect 22092 10386 22260 10388
rect 22092 10334 22206 10386
rect 22258 10334 22260 10386
rect 22092 10332 22260 10334
rect 22092 10052 22148 10332
rect 22204 10322 22260 10332
rect 21980 9996 22148 10052
rect 22652 10052 22708 10062
rect 22764 10052 22820 11116
rect 22876 10610 22932 10622
rect 22876 10558 22878 10610
rect 22930 10558 22932 10610
rect 22876 10164 22932 10558
rect 23100 10612 23156 10622
rect 23100 10518 23156 10556
rect 22988 10500 23044 10510
rect 22988 10406 23044 10444
rect 22876 10108 23156 10164
rect 22764 9996 23044 10052
rect 21868 9716 21924 9754
rect 21756 9658 21812 9670
rect 21756 9606 21758 9658
rect 21810 9606 21812 9658
rect 21868 9650 21924 9660
rect 21756 9604 21812 9606
rect 21532 9548 21812 9604
rect 21420 8866 21476 8876
rect 21980 8708 22036 9996
rect 22204 9884 22596 9940
rect 22092 9828 22148 9838
rect 22204 9828 22260 9884
rect 22092 9826 22260 9828
rect 22092 9774 22094 9826
rect 22146 9774 22260 9826
rect 22092 9772 22260 9774
rect 22540 9826 22596 9884
rect 22540 9774 22542 9826
rect 22594 9774 22596 9826
rect 22092 9762 22148 9772
rect 22540 9762 22596 9774
rect 22316 9716 22372 9726
rect 22316 9714 22484 9716
rect 22316 9662 22318 9714
rect 22370 9662 22484 9714
rect 22316 9660 22484 9662
rect 22316 9650 22372 9660
rect 22316 9492 22372 9502
rect 21980 8642 22036 8652
rect 22092 9436 22316 9492
rect 21308 8206 21310 8258
rect 21362 8206 21364 8258
rect 21308 8194 21364 8206
rect 21644 8372 21700 8382
rect 21532 8034 21588 8046
rect 21532 7982 21534 8034
rect 21586 7982 21588 8034
rect 21420 7700 21476 7710
rect 21196 7644 21420 7700
rect 21420 7606 21476 7644
rect 21532 7476 21588 7982
rect 21644 7642 21700 8316
rect 21756 8260 21812 8270
rect 21756 8166 21812 8204
rect 21868 8258 21924 8270
rect 21868 8206 21870 8258
rect 21922 8206 21924 8258
rect 21868 8148 21924 8206
rect 21868 8082 21924 8092
rect 21644 7590 21646 7642
rect 21698 7590 21700 7642
rect 21756 7700 21812 7710
rect 21756 7606 21812 7644
rect 21980 7700 22036 7710
rect 22092 7700 22148 9436
rect 22316 9426 22372 9436
rect 22428 9156 22484 9660
rect 22204 9100 22428 9156
rect 22204 8148 22260 9100
rect 22428 9062 22484 9100
rect 22652 9268 22708 9996
rect 22764 9716 22820 9726
rect 22764 9622 22820 9660
rect 22876 9714 22932 9726
rect 22876 9662 22878 9714
rect 22930 9662 22932 9714
rect 22652 9042 22708 9212
rect 22652 8990 22654 9042
rect 22706 8990 22708 9042
rect 22652 8978 22708 8990
rect 22876 8820 22932 9662
rect 22988 9154 23044 9996
rect 23100 9492 23156 10108
rect 23212 9828 23268 11228
rect 23996 10836 24052 10846
rect 23996 10742 24052 10780
rect 23436 10610 23492 10622
rect 23436 10558 23438 10610
rect 23490 10558 23492 10610
rect 23212 9762 23268 9772
rect 23324 10052 23380 10062
rect 23324 9826 23380 9996
rect 23324 9774 23326 9826
rect 23378 9774 23380 9826
rect 23324 9762 23380 9774
rect 23100 9426 23156 9436
rect 22988 9102 22990 9154
rect 23042 9102 23044 9154
rect 22988 9090 23044 9102
rect 23436 9156 23492 10558
rect 23996 9716 24052 9726
rect 23996 9622 24052 9660
rect 23996 9268 24052 9278
rect 24108 9268 24164 12348
rect 24052 9212 24164 9268
rect 24220 10836 24276 10846
rect 23996 9174 24052 9212
rect 23212 9042 23268 9054
rect 23212 8990 23214 9042
rect 23266 8990 23268 9042
rect 23100 8932 23156 8942
rect 23100 8838 23156 8876
rect 22652 8764 22932 8820
rect 22988 8820 23044 8830
rect 22316 8372 22372 8382
rect 22316 8258 22372 8316
rect 22316 8206 22318 8258
rect 22370 8206 22372 8258
rect 22316 8194 22372 8206
rect 22540 8372 22596 8382
rect 22204 8082 22260 8092
rect 22428 8148 22484 8158
rect 22540 8148 22596 8316
rect 22652 8258 22708 8764
rect 22988 8372 23044 8764
rect 22652 8206 22654 8258
rect 22706 8206 22708 8258
rect 22652 8194 22708 8206
rect 22764 8316 23044 8372
rect 22428 8146 22596 8148
rect 22428 8094 22430 8146
rect 22482 8094 22596 8146
rect 22428 8092 22596 8094
rect 22428 8082 22484 8092
rect 21980 7698 22148 7700
rect 21980 7646 21982 7698
rect 22034 7646 22148 7698
rect 21980 7644 22148 7646
rect 22652 7700 22708 7710
rect 22764 7700 22820 8316
rect 22652 7698 22820 7700
rect 22652 7646 22654 7698
rect 22706 7646 22820 7698
rect 22652 7644 22820 7646
rect 22876 8146 22932 8158
rect 22876 8094 22878 8146
rect 22930 8094 22932 8146
rect 22876 8036 22932 8094
rect 22988 8146 23044 8316
rect 23212 8258 23268 8990
rect 23436 9042 23492 9100
rect 23436 8990 23438 9042
rect 23490 8990 23492 9042
rect 23436 8978 23492 8990
rect 23548 8372 23604 8382
rect 23548 8278 23604 8316
rect 23212 8206 23214 8258
rect 23266 8206 23268 8258
rect 23212 8194 23268 8206
rect 22988 8094 22990 8146
rect 23042 8094 23044 8146
rect 22988 8082 23044 8094
rect 22876 7700 22932 7980
rect 22988 7700 23044 7710
rect 22876 7698 23044 7700
rect 22876 7646 22990 7698
rect 23042 7646 23044 7698
rect 22876 7644 23044 7646
rect 21980 7634 22036 7644
rect 22652 7634 22708 7644
rect 22988 7634 23044 7644
rect 21644 7578 21700 7590
rect 21532 7420 21812 7476
rect 21308 6692 21364 6702
rect 21756 6692 21812 7420
rect 21756 6636 22148 6692
rect 21308 5906 21364 6636
rect 22092 6018 22148 6636
rect 22092 5966 22094 6018
rect 22146 5966 22148 6018
rect 22092 5954 22148 5966
rect 21308 5854 21310 5906
rect 21362 5854 21364 5906
rect 21308 5842 21364 5854
rect 20972 5628 21476 5684
rect 20748 5234 20916 5236
rect 20748 5182 20750 5234
rect 20802 5182 20916 5234
rect 20748 5180 20916 5182
rect 20748 5170 20804 5180
rect 20300 4174 20302 4226
rect 20354 4174 20356 4226
rect 20300 4162 20356 4174
rect 21084 4114 21140 4126
rect 21084 4062 21086 4114
rect 21138 4062 21140 4114
rect 19740 3556 19796 3566
rect 19404 3554 19796 3556
rect 19404 3502 19742 3554
rect 19794 3502 19796 3554
rect 19404 3500 19796 3502
rect 19740 3490 19796 3500
rect 21084 3388 21140 4062
rect 21420 3554 21476 5628
rect 24220 5236 24276 10780
rect 24780 10052 24836 15092
rect 25340 14980 25396 15150
rect 25228 14644 25284 14654
rect 25340 14644 25396 14924
rect 25228 14642 25396 14644
rect 25228 14590 25230 14642
rect 25282 14590 25396 14642
rect 25228 14588 25396 14590
rect 25228 14578 25284 14588
rect 25452 13300 25508 13310
rect 25452 13074 25508 13244
rect 25452 13022 25454 13074
rect 25506 13022 25508 13074
rect 25452 13010 25508 13022
rect 25564 11844 25620 15260
rect 25676 14532 25732 15374
rect 25788 15204 25844 21310
rect 26012 18452 26068 18462
rect 26012 18358 26068 18396
rect 26348 16100 26404 16110
rect 25900 15876 25956 15886
rect 25900 15314 25956 15820
rect 25900 15262 25902 15314
rect 25954 15262 25956 15314
rect 25900 15250 25956 15262
rect 26348 15538 26404 16044
rect 26348 15486 26350 15538
rect 26402 15486 26404 15538
rect 25788 15138 25844 15148
rect 26348 14980 26404 15486
rect 26572 15316 26628 28812
rect 26908 28756 26964 28766
rect 26908 28662 26964 28700
rect 26908 27748 26964 27758
rect 27020 27748 27076 31892
rect 27244 31892 27300 32398
rect 27804 32004 27860 33180
rect 27916 33170 27972 33180
rect 28140 34076 28420 34132
rect 28476 35026 28532 35038
rect 28476 34974 28478 35026
rect 28530 34974 28532 35026
rect 28476 34692 28532 34974
rect 28140 32004 28196 34076
rect 28476 33234 28532 34636
rect 28700 34580 28756 37436
rect 29148 37044 29204 38892
rect 29260 38050 29316 38062
rect 29260 37998 29262 38050
rect 29314 37998 29316 38050
rect 29260 37940 29316 37998
rect 29260 37874 29316 37884
rect 29484 37938 29540 40012
rect 29708 38834 29764 40796
rect 30716 40516 30772 44200
rect 30716 40450 30772 40460
rect 31500 40514 31556 40526
rect 31500 40462 31502 40514
rect 31554 40462 31556 40514
rect 31164 40404 31220 40414
rect 31164 40402 31444 40404
rect 31164 40350 31166 40402
rect 31218 40350 31444 40402
rect 31164 40348 31444 40350
rect 31164 40338 31220 40348
rect 31276 39620 31332 39630
rect 30828 39618 31332 39620
rect 30828 39566 31278 39618
rect 31330 39566 31332 39618
rect 30828 39564 31332 39566
rect 30828 39058 30884 39564
rect 31276 39554 31332 39564
rect 30828 39006 30830 39058
rect 30882 39006 30884 39058
rect 30828 38994 30884 39006
rect 29708 38782 29710 38834
rect 29762 38782 29764 38834
rect 29708 38770 29764 38782
rect 30044 38836 30100 38846
rect 30044 38742 30100 38780
rect 30604 38836 30660 38846
rect 31164 38836 31220 38846
rect 30604 38834 30884 38836
rect 30604 38782 30606 38834
rect 30658 38782 30884 38834
rect 30604 38780 30884 38782
rect 30604 38770 30660 38780
rect 29484 37886 29486 37938
rect 29538 37886 29540 37938
rect 29484 37874 29540 37886
rect 29148 36978 29204 36988
rect 29148 35924 29204 35934
rect 28700 34514 28756 34524
rect 28812 35698 28868 35710
rect 28812 35646 28814 35698
rect 28866 35646 28868 35698
rect 28812 35364 28868 35646
rect 28588 33906 28644 33918
rect 28588 33854 28590 33906
rect 28642 33854 28644 33906
rect 28588 33460 28644 33854
rect 28588 33394 28644 33404
rect 28476 33182 28478 33234
rect 28530 33182 28532 33234
rect 28476 33170 28532 33182
rect 27804 31938 27860 31948
rect 27916 31948 28196 32004
rect 28252 32004 28308 32014
rect 28812 31948 28868 35308
rect 29148 34356 29204 35868
rect 29596 35588 29652 35598
rect 29596 35494 29652 35532
rect 29932 34356 29988 34366
rect 29148 34354 29988 34356
rect 29148 34302 29934 34354
rect 29986 34302 29988 34354
rect 29148 34300 29988 34302
rect 28924 34242 28980 34254
rect 28924 34190 28926 34242
rect 28978 34190 28980 34242
rect 28924 33796 28980 34190
rect 29148 34242 29204 34300
rect 29932 34290 29988 34300
rect 30828 34354 30884 38780
rect 31164 38742 31220 38780
rect 30828 34302 30830 34354
rect 30882 34302 30884 34354
rect 30828 34290 30884 34302
rect 29148 34190 29150 34242
rect 29202 34190 29204 34242
rect 29148 34178 29204 34190
rect 30380 34018 30436 34030
rect 30380 33966 30382 34018
rect 30434 33966 30436 34018
rect 28924 33730 28980 33740
rect 29372 33796 29428 33806
rect 29260 33122 29316 33134
rect 29260 33070 29262 33122
rect 29314 33070 29316 33122
rect 29260 32900 29316 33070
rect 29260 32834 29316 32844
rect 27244 31826 27300 31836
rect 27692 31556 27748 31566
rect 27692 31218 27748 31500
rect 27692 31166 27694 31218
rect 27746 31166 27748 31218
rect 27692 31154 27748 31166
rect 27916 30772 27972 31948
rect 28140 31556 28196 31566
rect 28140 31218 28196 31500
rect 28140 31166 28142 31218
rect 28194 31166 28196 31218
rect 28140 31154 28196 31166
rect 28028 30994 28084 31006
rect 28028 30942 28030 30994
rect 28082 30942 28084 30994
rect 28028 30884 28084 30942
rect 28028 30828 28196 30884
rect 27916 30716 28084 30772
rect 27916 30212 27972 30222
rect 27916 30118 27972 30156
rect 27580 30098 27636 30110
rect 27580 30046 27582 30098
rect 27634 30046 27636 30098
rect 27132 29988 27188 29998
rect 27132 29986 27524 29988
rect 27132 29934 27134 29986
rect 27186 29934 27524 29986
rect 27132 29932 27524 29934
rect 27132 29922 27188 29932
rect 27132 29314 27188 29326
rect 27132 29262 27134 29314
rect 27186 29262 27188 29314
rect 27132 28420 27188 29262
rect 27356 28756 27412 28766
rect 27468 28756 27524 29932
rect 27412 28700 27524 28756
rect 27356 28690 27412 28700
rect 27244 28644 27300 28654
rect 27244 28550 27300 28588
rect 27580 28644 27636 30046
rect 27692 29986 27748 29998
rect 27692 29934 27694 29986
rect 27746 29934 27748 29986
rect 27692 29876 27748 29934
rect 27692 28868 27748 29820
rect 27692 28802 27748 28812
rect 28028 28644 28084 30716
rect 28140 30100 28196 30828
rect 28252 30212 28308 31948
rect 28700 31892 28868 31948
rect 29260 31892 29316 31902
rect 28700 31826 28756 31836
rect 29260 31778 29316 31836
rect 29260 31726 29262 31778
rect 29314 31726 29316 31778
rect 29260 31714 29316 31726
rect 28700 31668 28756 31678
rect 28700 31218 28756 31612
rect 28700 31166 28702 31218
rect 28754 31166 28756 31218
rect 28700 31154 28756 31166
rect 28364 31108 28420 31118
rect 28364 31106 28532 31108
rect 28364 31054 28366 31106
rect 28418 31054 28532 31106
rect 28364 31052 28532 31054
rect 28364 31042 28420 31052
rect 28476 30994 28532 31052
rect 28476 30942 28478 30994
rect 28530 30942 28532 30994
rect 28476 30930 28532 30942
rect 28812 30994 28868 31006
rect 28812 30942 28814 30994
rect 28866 30942 28868 30994
rect 28812 30212 28868 30942
rect 29148 30996 29204 31006
rect 29148 30994 29316 30996
rect 29148 30942 29150 30994
rect 29202 30942 29316 30994
rect 29148 30940 29316 30942
rect 29148 30930 29204 30940
rect 28252 30156 28420 30212
rect 28140 30034 28196 30044
rect 28252 29986 28308 29998
rect 28252 29934 28254 29986
rect 28306 29934 28308 29986
rect 28252 29876 28308 29934
rect 28252 29810 28308 29820
rect 28028 28588 28308 28644
rect 27580 28578 27636 28588
rect 27804 28532 27860 28542
rect 27804 28438 27860 28476
rect 27356 28420 27412 28430
rect 27132 28418 27524 28420
rect 27132 28366 27358 28418
rect 27410 28366 27524 28418
rect 27132 28364 27524 28366
rect 27356 28354 27412 28364
rect 27356 28196 27412 28206
rect 27244 27858 27300 27870
rect 27244 27806 27246 27858
rect 27298 27806 27300 27858
rect 27244 27748 27300 27806
rect 26908 27746 27300 27748
rect 26908 27694 26910 27746
rect 26962 27694 27300 27746
rect 26908 27692 27300 27694
rect 26908 27682 26964 27692
rect 27132 25732 27188 25742
rect 27020 25396 27076 25406
rect 27020 25302 27076 25340
rect 27020 24612 27076 24622
rect 26796 22370 26852 22382
rect 26796 22318 26798 22370
rect 26850 22318 26852 22370
rect 26684 21588 26740 21598
rect 26684 21364 26740 21532
rect 26684 21298 26740 21308
rect 26796 20804 26852 22318
rect 26908 22372 26964 22410
rect 26908 22306 26964 22316
rect 27020 22146 27076 24556
rect 27132 22370 27188 25676
rect 27132 22318 27134 22370
rect 27186 22318 27188 22370
rect 27132 22260 27188 22318
rect 27132 22194 27188 22204
rect 27020 22094 27022 22146
rect 27074 22094 27076 22146
rect 27020 22082 27076 22094
rect 27132 22036 27188 22046
rect 27020 21924 27076 21934
rect 27020 21810 27076 21868
rect 27020 21758 27022 21810
rect 27074 21758 27076 21810
rect 27020 21746 27076 21758
rect 27132 21028 27188 21980
rect 26796 20738 26852 20748
rect 27020 20972 27188 21028
rect 27244 21476 27300 27692
rect 27356 26402 27412 28140
rect 27356 26350 27358 26402
rect 27410 26350 27412 26402
rect 27356 26338 27412 26350
rect 27356 23044 27412 23054
rect 27468 23044 27524 28364
rect 27580 28418 27636 28430
rect 27580 28366 27582 28418
rect 27634 28366 27636 28418
rect 27580 26402 27636 28366
rect 27916 28418 27972 28430
rect 28140 28420 28196 28430
rect 27916 28366 27918 28418
rect 27970 28366 27972 28418
rect 27916 28308 27972 28366
rect 27916 27300 27972 28252
rect 27916 27234 27972 27244
rect 28028 28418 28196 28420
rect 28028 28366 28142 28418
rect 28194 28366 28196 28418
rect 28028 28364 28196 28366
rect 27804 26962 27860 26974
rect 27804 26910 27806 26962
rect 27858 26910 27860 26962
rect 27804 26514 27860 26910
rect 27804 26462 27806 26514
rect 27858 26462 27860 26514
rect 27804 26450 27860 26462
rect 27580 26350 27582 26402
rect 27634 26350 27636 26402
rect 27580 26338 27636 26350
rect 28028 26290 28084 28364
rect 28140 28354 28196 28364
rect 28252 26908 28308 28588
rect 28028 26238 28030 26290
rect 28082 26238 28084 26290
rect 28028 26226 28084 26238
rect 28140 26852 28308 26908
rect 27692 24612 27748 24622
rect 27692 24518 27748 24556
rect 27356 23042 27524 23044
rect 27356 22990 27358 23042
rect 27410 22990 27524 23042
rect 27356 22988 27524 22990
rect 27356 22978 27412 22988
rect 27356 22484 27412 22494
rect 27356 22370 27412 22428
rect 27356 22318 27358 22370
rect 27410 22318 27412 22370
rect 27356 22306 27412 22318
rect 27468 22148 27524 22988
rect 28028 23044 28084 23054
rect 28028 22950 28084 22988
rect 27692 22482 27748 22494
rect 27692 22430 27694 22482
rect 27746 22430 27748 22482
rect 27692 22372 27748 22430
rect 27804 22484 27860 22494
rect 27860 22428 27972 22484
rect 27804 22418 27860 22428
rect 27692 22306 27748 22316
rect 27804 22148 27860 22158
rect 27468 22146 27860 22148
rect 27468 22094 27806 22146
rect 27858 22094 27860 22146
rect 27468 22092 27860 22094
rect 27356 21700 27412 21710
rect 27356 21606 27412 21644
rect 27020 19236 27076 20972
rect 27132 20804 27188 20814
rect 27132 20710 27188 20748
rect 27020 19170 27076 19180
rect 27244 19348 27300 21420
rect 27468 21364 27524 21374
rect 27468 21026 27524 21308
rect 27468 20974 27470 21026
rect 27522 20974 27524 21026
rect 27468 20962 27524 20974
rect 27580 20580 27636 22092
rect 27804 22082 27860 22092
rect 27692 21812 27748 21822
rect 27916 21812 27972 22428
rect 28028 22258 28084 22270
rect 28028 22206 28030 22258
rect 28082 22206 28084 22258
rect 28028 21924 28084 22206
rect 28140 22036 28196 26852
rect 28364 23156 28420 30156
rect 28812 30146 28868 30156
rect 29260 30212 29316 30940
rect 29260 30146 29316 30156
rect 29036 30100 29092 30110
rect 29148 30100 29204 30110
rect 29092 30098 29204 30100
rect 29092 30046 29150 30098
rect 29202 30046 29204 30098
rect 29092 30044 29204 30046
rect 28924 29314 28980 29326
rect 28924 29262 28926 29314
rect 28978 29262 28980 29314
rect 28588 28418 28644 28430
rect 28588 28366 28590 28418
rect 28642 28366 28644 28418
rect 28588 28308 28644 28366
rect 28588 28242 28644 28252
rect 28924 27524 28980 29262
rect 29036 28644 29092 30044
rect 29148 30034 29204 30044
rect 29260 29986 29316 29998
rect 29260 29934 29262 29986
rect 29314 29934 29316 29986
rect 29260 29652 29316 29934
rect 29260 29586 29316 29596
rect 29036 28578 29092 28588
rect 29148 28530 29204 28542
rect 29148 28478 29150 28530
rect 29202 28478 29204 28530
rect 29148 28420 29204 28478
rect 29148 28354 29204 28364
rect 29260 28418 29316 28430
rect 29260 28366 29262 28418
rect 29314 28366 29316 28418
rect 29260 27524 29316 28366
rect 28700 27468 29316 27524
rect 29372 27524 29428 33740
rect 30380 33796 30436 33966
rect 31164 33908 31220 33918
rect 31164 33814 31220 33852
rect 30380 33730 30436 33740
rect 31388 33684 31444 40348
rect 31500 40292 31556 40462
rect 31500 40226 31556 40236
rect 31836 39844 31892 44200
rect 32956 41972 33012 44200
rect 32956 41906 33012 41916
rect 33180 41412 33236 41422
rect 33180 41318 33236 41356
rect 32172 41186 32228 41198
rect 32396 41188 32452 41198
rect 32172 41134 32174 41186
rect 32226 41134 32228 41186
rect 32172 40404 32228 41134
rect 32172 40338 32228 40348
rect 32284 41132 32396 41188
rect 31836 39778 31892 39788
rect 32060 39620 32116 39630
rect 31500 39618 32116 39620
rect 31500 39566 32062 39618
rect 32114 39566 32116 39618
rect 31500 39564 32116 39566
rect 31500 39058 31556 39564
rect 32060 39554 32116 39564
rect 31500 39006 31502 39058
rect 31554 39006 31556 39058
rect 31500 38994 31556 39006
rect 32172 39060 32228 39070
rect 32284 39060 32340 41132
rect 32396 41122 32452 41132
rect 34076 41076 34132 44200
rect 35196 41748 35252 44200
rect 36316 41860 36372 44200
rect 36988 41972 37044 41982
rect 36316 41804 36484 41860
rect 34076 41010 34132 41020
rect 35084 41692 35252 41748
rect 34076 40628 34132 40638
rect 34076 40534 34132 40572
rect 33068 40402 33124 40414
rect 33068 40350 33070 40402
rect 33122 40350 33124 40402
rect 33068 40068 33124 40350
rect 33068 40002 33124 40012
rect 33404 40404 33460 40414
rect 33068 39844 33124 39854
rect 33068 39750 33124 39788
rect 32172 39058 32340 39060
rect 32172 39006 32174 39058
rect 32226 39006 32340 39058
rect 32172 39004 32340 39006
rect 33404 39058 33460 40348
rect 33404 39006 33406 39058
rect 33458 39006 33460 39058
rect 32172 38994 32228 39004
rect 33404 38994 33460 39006
rect 34972 39506 35028 39518
rect 34972 39454 34974 39506
rect 35026 39454 35028 39506
rect 31948 38834 32004 38846
rect 31948 38782 31950 38834
rect 32002 38782 32004 38834
rect 31836 38724 31892 38734
rect 31052 33628 31444 33684
rect 31500 37828 31556 37838
rect 30156 33460 30212 33470
rect 30156 33366 30212 33404
rect 31052 31948 31108 33628
rect 31500 31948 31556 37772
rect 31724 36260 31780 36270
rect 31724 35586 31780 36204
rect 31724 35534 31726 35586
rect 31778 35534 31780 35586
rect 31724 34356 31780 35534
rect 31724 34242 31780 34300
rect 31724 34190 31726 34242
rect 31778 34190 31780 34242
rect 31724 34178 31780 34190
rect 30716 31892 31108 31948
rect 31388 31892 31556 31948
rect 29932 31668 29988 31678
rect 29932 31574 29988 31612
rect 30492 30436 30548 30446
rect 30380 30434 30548 30436
rect 30380 30382 30494 30434
rect 30546 30382 30548 30434
rect 30380 30380 30548 30382
rect 29484 30212 29540 30222
rect 29708 30212 29764 30222
rect 29484 30210 29764 30212
rect 29484 30158 29486 30210
rect 29538 30158 29710 30210
rect 29762 30158 29764 30210
rect 29484 30156 29764 30158
rect 29484 30146 29540 30156
rect 29708 30146 29764 30156
rect 30044 30210 30100 30222
rect 30044 30158 30046 30210
rect 30098 30158 30100 30210
rect 29932 30100 29988 30110
rect 29932 30006 29988 30044
rect 30044 29316 30100 30158
rect 29484 29260 30100 29316
rect 30268 30212 30324 30222
rect 29484 28642 29540 29260
rect 29484 28590 29486 28642
rect 29538 28590 29540 28642
rect 29484 28578 29540 28590
rect 29708 29092 29764 29102
rect 29372 27468 29652 27524
rect 28588 27076 28644 27086
rect 28588 26982 28644 27020
rect 28476 25060 28532 25070
rect 28700 25060 28756 27468
rect 28812 27300 28868 27310
rect 28812 26514 28868 27244
rect 29372 27300 29428 27310
rect 29372 27206 29428 27244
rect 28812 26462 28814 26514
rect 28866 26462 28868 26514
rect 28812 26450 28868 26462
rect 29148 27074 29204 27086
rect 29148 27022 29150 27074
rect 29202 27022 29204 27074
rect 29148 25732 29204 27022
rect 29148 25666 29204 25676
rect 29260 27076 29316 27086
rect 29260 26514 29316 27020
rect 29596 26908 29652 27468
rect 29708 27298 29764 29036
rect 29820 28756 29876 28766
rect 29820 28642 29876 28700
rect 30268 28756 30324 30156
rect 30268 28690 30324 28700
rect 29820 28590 29822 28642
rect 29874 28590 29876 28642
rect 29820 28578 29876 28590
rect 30156 28642 30212 28654
rect 30156 28590 30158 28642
rect 30210 28590 30212 28642
rect 29708 27246 29710 27298
rect 29762 27246 29764 27298
rect 29708 27234 29764 27246
rect 30044 28420 30100 28430
rect 30044 27074 30100 28364
rect 30156 27298 30212 28590
rect 30268 28420 30324 28430
rect 30268 28326 30324 28364
rect 30156 27246 30158 27298
rect 30210 27246 30212 27298
rect 30156 27234 30212 27246
rect 30044 27022 30046 27074
rect 30098 27022 30100 27074
rect 30044 27010 30100 27022
rect 30380 26908 30436 30380
rect 30492 30370 30548 30380
rect 30716 29092 30772 31892
rect 31052 30884 31108 30894
rect 31276 30884 31332 30894
rect 30940 30882 31332 30884
rect 30940 30830 31054 30882
rect 31106 30830 31278 30882
rect 31330 30830 31332 30882
rect 30940 30828 31332 30830
rect 30940 30434 30996 30828
rect 31052 30818 31108 30828
rect 31276 30818 31332 30828
rect 30940 30382 30942 30434
rect 30994 30382 30996 30434
rect 30940 30370 30996 30382
rect 30828 30212 30884 30222
rect 31164 30212 31220 30222
rect 30828 30210 31220 30212
rect 30828 30158 30830 30210
rect 30882 30158 31166 30210
rect 31218 30158 31220 30210
rect 30828 30156 31220 30158
rect 30828 30146 30884 30156
rect 30716 29026 30772 29036
rect 30828 28866 30884 28878
rect 30828 28814 30830 28866
rect 30882 28814 30884 28866
rect 30828 28756 30884 28814
rect 30604 28700 30884 28756
rect 30492 28644 30548 28654
rect 30604 28644 30660 28700
rect 30492 28642 30660 28644
rect 30492 28590 30494 28642
rect 30546 28590 30660 28642
rect 30492 28588 30660 28590
rect 30492 28578 30548 28588
rect 30716 28532 30772 28542
rect 30716 28438 30772 28476
rect 30828 28418 30884 28430
rect 30828 28366 30830 28418
rect 30882 28366 30884 28418
rect 30828 28196 30884 28366
rect 30716 28140 30884 28196
rect 30716 27972 30772 28140
rect 30940 27972 30996 30156
rect 31164 30146 31220 30156
rect 30716 27906 30772 27916
rect 30828 27970 30996 27972
rect 30828 27918 30942 27970
rect 30994 27918 30996 27970
rect 30828 27916 30996 27918
rect 30828 27860 30884 27916
rect 30940 27906 30996 27916
rect 30828 27076 30884 27804
rect 30828 26982 30884 27020
rect 29596 26852 29876 26908
rect 29260 26462 29262 26514
rect 29314 26462 29316 26514
rect 28476 24722 28532 25004
rect 28476 24670 28478 24722
rect 28530 24670 28532 24722
rect 28476 24658 28532 24670
rect 28588 25004 28756 25060
rect 28924 25060 28980 25070
rect 28588 23268 28644 25004
rect 28924 24948 28980 25004
rect 29260 24948 29316 26462
rect 28924 24946 29316 24948
rect 28924 24894 28926 24946
rect 28978 24894 29316 24946
rect 28924 24892 29316 24894
rect 28924 24882 28980 24892
rect 28140 21970 28196 21980
rect 28252 23100 28420 23156
rect 28476 23212 28644 23268
rect 28700 24724 28756 24734
rect 29260 24724 29316 24892
rect 29372 24948 29428 24958
rect 29428 24892 29540 24948
rect 29372 24882 29428 24892
rect 29372 24724 29428 24734
rect 29260 24722 29428 24724
rect 29260 24670 29374 24722
rect 29426 24670 29428 24722
rect 29260 24668 29428 24670
rect 28028 21858 28084 21868
rect 27692 21810 27972 21812
rect 27692 21758 27694 21810
rect 27746 21758 27972 21810
rect 27692 21756 27972 21758
rect 27692 21746 27748 21756
rect 27692 21028 27748 21038
rect 27692 20802 27748 20972
rect 27692 20750 27694 20802
rect 27746 20750 27748 20802
rect 27692 20738 27748 20750
rect 27916 20802 27972 21756
rect 28140 21698 28196 21710
rect 28140 21646 28142 21698
rect 28194 21646 28196 21698
rect 28140 21588 28196 21646
rect 28028 21364 28084 21374
rect 28028 21270 28084 21308
rect 27916 20750 27918 20802
rect 27970 20750 27972 20802
rect 27916 20738 27972 20750
rect 27580 20524 27748 20580
rect 26908 16548 26964 16558
rect 26908 15876 26964 16492
rect 26908 15874 27076 15876
rect 26908 15822 26910 15874
rect 26962 15822 27076 15874
rect 26908 15820 27076 15822
rect 26908 15810 26964 15820
rect 26908 15316 26964 15326
rect 26628 15314 26964 15316
rect 26628 15262 26910 15314
rect 26962 15262 26964 15314
rect 26628 15260 26964 15262
rect 26572 15222 26628 15260
rect 26908 15250 26964 15260
rect 27020 15316 27076 15820
rect 26404 14924 26740 14980
rect 26348 14914 26404 14924
rect 26012 14532 26068 14542
rect 26572 14532 26628 14542
rect 25732 14530 26628 14532
rect 25732 14478 26014 14530
rect 26066 14478 26574 14530
rect 26626 14478 26628 14530
rect 25732 14476 26628 14478
rect 25676 14466 25732 14476
rect 26012 14466 26068 14476
rect 26572 14466 26628 14476
rect 26684 14418 26740 14924
rect 27020 14756 27076 15260
rect 26684 14366 26686 14418
rect 26738 14366 26740 14418
rect 26684 14354 26740 14366
rect 26796 14700 27076 14756
rect 25676 14308 25732 14318
rect 26124 14308 26180 14318
rect 26348 14308 26404 14318
rect 25676 14306 26124 14308
rect 25676 14254 25678 14306
rect 25730 14254 26124 14306
rect 25676 14252 26124 14254
rect 25676 13972 25732 14252
rect 26124 14214 26180 14252
rect 26236 14306 26404 14308
rect 26236 14254 26350 14306
rect 26402 14254 26404 14306
rect 26236 14252 26404 14254
rect 25676 13906 25732 13916
rect 26012 13860 26068 13870
rect 26012 13766 26068 13804
rect 26236 13412 26292 14252
rect 26348 14242 26404 14252
rect 26348 14084 26404 14094
rect 26348 13858 26404 14028
rect 26348 13806 26350 13858
rect 26402 13806 26404 13858
rect 26348 13794 26404 13806
rect 26460 13860 26516 13870
rect 26460 13766 26516 13804
rect 26236 13346 26292 13356
rect 26684 13746 26740 13758
rect 26684 13694 26686 13746
rect 26738 13694 26740 13746
rect 26684 12964 26740 13694
rect 26684 12898 26740 12908
rect 26348 12404 26404 12414
rect 26348 12310 26404 12348
rect 24332 9996 24836 10052
rect 25116 11788 25620 11844
rect 24332 9604 24388 9996
rect 25116 9940 25172 11788
rect 26796 10164 26852 14700
rect 26908 14420 26964 14430
rect 26908 14326 26964 14364
rect 27132 14418 27188 14430
rect 27132 14366 27134 14418
rect 27186 14366 27188 14418
rect 27132 14196 27188 14366
rect 27132 14130 27188 14140
rect 27244 13860 27300 19292
rect 27356 17108 27412 17118
rect 27580 17108 27636 17118
rect 27412 17106 27636 17108
rect 27412 17054 27582 17106
rect 27634 17054 27636 17106
rect 27412 17052 27636 17054
rect 27356 17014 27412 17052
rect 27580 17042 27636 17052
rect 27580 15876 27636 15886
rect 27580 15426 27636 15820
rect 27580 15374 27582 15426
rect 27634 15374 27636 15426
rect 27580 15362 27636 15374
rect 27356 15316 27412 15326
rect 27356 15222 27412 15260
rect 27468 15204 27524 15214
rect 27356 14420 27412 14430
rect 27356 14326 27412 14364
rect 27468 14196 27524 15148
rect 27692 14644 27748 20524
rect 27804 20578 27860 20590
rect 27804 20526 27806 20578
rect 27858 20526 27860 20578
rect 27804 18564 27860 20526
rect 28028 20132 28084 20142
rect 28028 20038 28084 20076
rect 27804 18498 27860 18508
rect 27916 19794 27972 19806
rect 28140 19796 28196 21532
rect 27916 19742 27918 19794
rect 27970 19742 27972 19794
rect 27916 18340 27972 19742
rect 27804 18284 27972 18340
rect 28028 19740 28196 19796
rect 27804 15428 27860 18284
rect 27916 16994 27972 17006
rect 27916 16942 27918 16994
rect 27970 16942 27972 16994
rect 27916 16772 27972 16942
rect 27916 16706 27972 16716
rect 28028 16100 28084 19740
rect 28140 19236 28196 19246
rect 28140 18338 28196 19180
rect 28140 18286 28142 18338
rect 28194 18286 28196 18338
rect 28140 18274 28196 18286
rect 28028 16034 28084 16044
rect 28140 17108 28196 17118
rect 28140 16210 28196 17052
rect 28140 16158 28142 16210
rect 28194 16158 28196 16210
rect 28140 15876 28196 16158
rect 28140 15810 28196 15820
rect 27804 15372 27972 15428
rect 27804 15204 27860 15242
rect 27804 15138 27860 15148
rect 27916 14644 27972 15372
rect 28252 15316 28308 23100
rect 28364 22930 28420 22942
rect 28364 22878 28366 22930
rect 28418 22878 28420 22930
rect 28364 21924 28420 22878
rect 28476 22372 28532 23212
rect 28700 23156 28756 24668
rect 29372 24658 29428 24668
rect 29484 24164 29540 24892
rect 29372 24108 29540 24164
rect 29372 24052 29428 24108
rect 29372 23958 29428 23996
rect 29708 24052 29764 24062
rect 29708 23938 29764 23996
rect 29708 23886 29710 23938
rect 29762 23886 29764 23938
rect 29708 23874 29764 23886
rect 29484 23828 29540 23838
rect 29820 23828 29876 26852
rect 30156 26850 30212 26862
rect 30156 26798 30158 26850
rect 30210 26798 30212 26850
rect 30156 24836 30212 26798
rect 30156 24770 30212 24780
rect 30268 26852 30436 26908
rect 30156 24610 30212 24622
rect 30156 24558 30158 24610
rect 30210 24558 30212 24610
rect 30156 23828 30212 24558
rect 29820 23772 29988 23828
rect 29484 23378 29540 23772
rect 29484 23326 29486 23378
rect 29538 23326 29540 23378
rect 29484 23314 29540 23326
rect 29596 23492 29652 23502
rect 28588 23154 28756 23156
rect 28588 23102 28702 23154
rect 28754 23102 28756 23154
rect 28588 23100 28756 23102
rect 28588 22484 28644 23100
rect 28700 23090 28756 23100
rect 29036 23156 29092 23166
rect 29036 23062 29092 23100
rect 29372 23156 29428 23166
rect 28700 22932 28756 22942
rect 29260 22932 29316 22942
rect 28700 22930 29316 22932
rect 28700 22878 28702 22930
rect 28754 22878 29262 22930
rect 29314 22878 29316 22930
rect 28700 22876 29316 22878
rect 28700 22866 28756 22876
rect 29260 22866 29316 22876
rect 29372 22484 29428 23100
rect 29596 23154 29652 23436
rect 29596 23102 29598 23154
rect 29650 23102 29652 23154
rect 29484 22932 29540 22942
rect 29484 22594 29540 22876
rect 29484 22542 29486 22594
rect 29538 22542 29540 22594
rect 29484 22530 29540 22542
rect 28588 22428 29316 22484
rect 28476 22316 28644 22372
rect 28588 22258 28644 22316
rect 28588 22206 28590 22258
rect 28642 22206 28644 22258
rect 28364 21698 28420 21868
rect 28364 21646 28366 21698
rect 28418 21646 28420 21698
rect 28364 21634 28420 21646
rect 28476 22148 28532 22158
rect 28364 21028 28420 21038
rect 28364 20914 28420 20972
rect 28364 20862 28366 20914
rect 28418 20862 28420 20914
rect 28364 20850 28420 20862
rect 28476 20692 28532 22092
rect 28588 21812 28644 22206
rect 28588 20916 28644 21756
rect 28812 21588 28868 21598
rect 28812 21494 28868 21532
rect 28588 20850 28644 20860
rect 28812 21028 28868 21038
rect 28364 20636 28532 20692
rect 28364 19794 28420 20636
rect 28364 19742 28366 19794
rect 28418 19742 28420 19794
rect 28364 19730 28420 19742
rect 28476 19906 28532 19918
rect 28476 19854 28478 19906
rect 28530 19854 28532 19906
rect 28476 19796 28532 19854
rect 28476 16212 28532 19740
rect 28588 19348 28644 19358
rect 28588 19254 28644 19292
rect 28700 18338 28756 18350
rect 28700 18286 28702 18338
rect 28754 18286 28756 18338
rect 28588 17780 28644 17790
rect 28588 17686 28644 17724
rect 28700 16884 28756 18286
rect 28812 17108 28868 20972
rect 28812 17042 28868 17052
rect 28700 16818 28756 16828
rect 28924 16772 28980 22428
rect 29148 22258 29204 22270
rect 29148 22206 29150 22258
rect 29202 22206 29204 22258
rect 29148 21924 29204 22206
rect 29148 21858 29204 21868
rect 29260 21700 29316 22428
rect 29372 22418 29428 22428
rect 29372 22146 29428 22158
rect 29372 22094 29374 22146
rect 29426 22094 29428 22146
rect 29372 21924 29428 22094
rect 29596 22148 29652 23102
rect 29820 23156 29876 23166
rect 29820 23062 29876 23100
rect 29708 23044 29764 23054
rect 29708 22820 29764 22988
rect 29932 22932 29988 23772
rect 30156 23762 30212 23772
rect 30044 23714 30100 23726
rect 30044 23662 30046 23714
rect 30098 23662 30100 23714
rect 30044 23380 30100 23662
rect 30044 23314 30100 23324
rect 30156 23156 30212 23166
rect 30156 23062 30212 23100
rect 29932 22876 30212 22932
rect 29708 22764 29988 22820
rect 29932 22482 29988 22764
rect 29932 22430 29934 22482
rect 29986 22430 29988 22482
rect 29932 22418 29988 22430
rect 29596 22082 29652 22092
rect 29372 21858 29428 21868
rect 29932 21924 29988 21934
rect 29260 21644 29876 21700
rect 29372 21476 29428 21486
rect 29260 21474 29428 21476
rect 29260 21422 29374 21474
rect 29426 21422 29428 21474
rect 29260 21420 29428 21422
rect 29260 20804 29316 21420
rect 29372 21410 29428 21420
rect 29148 20748 29260 20804
rect 29036 20132 29092 20142
rect 29036 20038 29092 20076
rect 29148 19796 29204 20748
rect 29260 20710 29316 20748
rect 29596 20692 29652 20702
rect 29372 20636 29596 20692
rect 29260 20244 29316 20254
rect 29372 20244 29428 20636
rect 29596 20598 29652 20636
rect 29820 20690 29876 21644
rect 29932 21026 29988 21868
rect 29932 20974 29934 21026
rect 29986 20974 29988 21026
rect 29932 20962 29988 20974
rect 29820 20638 29822 20690
rect 29874 20638 29876 20690
rect 29820 20626 29876 20638
rect 30044 20692 30100 20702
rect 29260 20242 29428 20244
rect 29260 20190 29262 20242
rect 29314 20190 29428 20242
rect 29260 20188 29428 20190
rect 30044 20242 30100 20636
rect 30044 20190 30046 20242
rect 30098 20190 30100 20242
rect 29260 20178 29316 20188
rect 30044 20178 30100 20190
rect 29484 20020 29540 20030
rect 29708 20020 29764 20030
rect 29484 20018 29764 20020
rect 29484 19966 29486 20018
rect 29538 19966 29710 20018
rect 29762 19966 29764 20018
rect 29484 19964 29764 19966
rect 29372 19908 29428 19918
rect 29372 19814 29428 19852
rect 29260 19796 29316 19806
rect 29148 19740 29260 19796
rect 29260 19730 29316 19740
rect 29484 19796 29540 19964
rect 29708 19954 29764 19964
rect 29484 19730 29540 19740
rect 29148 19348 29204 19358
rect 29148 19234 29204 19292
rect 29148 19182 29150 19234
rect 29202 19182 29204 19234
rect 29148 19170 29204 19182
rect 29260 17108 29316 17118
rect 29260 17014 29316 17052
rect 29148 16884 29204 16894
rect 29148 16790 29204 16828
rect 28980 16716 29092 16772
rect 28924 16706 28980 16716
rect 29036 16436 29092 16716
rect 29036 16380 29316 16436
rect 28476 16146 28532 16156
rect 29148 15988 29204 15998
rect 29148 15894 29204 15932
rect 29260 15986 29316 16380
rect 29596 16156 29988 16212
rect 29484 16100 29540 16110
rect 29596 16100 29652 16156
rect 29484 16098 29652 16100
rect 29484 16046 29486 16098
rect 29538 16046 29652 16098
rect 29484 16044 29652 16046
rect 29932 16098 29988 16156
rect 29932 16046 29934 16098
rect 29986 16046 29988 16098
rect 29484 16034 29540 16044
rect 29932 16034 29988 16046
rect 29708 15988 29764 15998
rect 29260 15934 29262 15986
rect 29314 15934 29316 15986
rect 29260 15922 29316 15934
rect 29596 15986 29764 15988
rect 29596 15934 29710 15986
rect 29762 15934 29764 15986
rect 29596 15932 29764 15934
rect 29596 15652 29652 15932
rect 29708 15922 29764 15932
rect 29932 15876 29988 15886
rect 29932 15874 30100 15876
rect 29932 15822 29934 15874
rect 29986 15822 30100 15874
rect 29932 15820 30100 15822
rect 29932 15810 29988 15820
rect 28924 15596 29652 15652
rect 28924 15538 28980 15596
rect 28924 15486 28926 15538
rect 28978 15486 28980 15538
rect 28924 15474 28980 15486
rect 29708 15540 29764 15550
rect 28700 15426 28756 15438
rect 28700 15374 28702 15426
rect 28754 15374 28756 15426
rect 28140 15260 28308 15316
rect 28588 15314 28644 15326
rect 28588 15262 28590 15314
rect 28642 15262 28644 15314
rect 27916 14588 28084 14644
rect 27692 14578 27748 14588
rect 27692 14420 27748 14430
rect 27916 14420 27972 14430
rect 27692 14418 27972 14420
rect 27692 14366 27694 14418
rect 27746 14366 27918 14418
rect 27970 14366 27972 14418
rect 27692 14364 27972 14366
rect 27692 14354 27748 14364
rect 27916 14354 27972 14364
rect 27132 13804 27300 13860
rect 27356 14140 27524 14196
rect 27580 14306 27636 14318
rect 27580 14254 27582 14306
rect 27634 14254 27636 14306
rect 27020 13748 27076 13758
rect 27020 13654 27076 13692
rect 27132 12404 27188 13804
rect 27244 12964 27300 12974
rect 27244 12870 27300 12908
rect 27132 12178 27188 12348
rect 27132 12126 27134 12178
rect 27186 12126 27188 12178
rect 27132 12114 27188 12126
rect 26124 10108 26852 10164
rect 27244 11732 27300 11742
rect 27244 10610 27300 11676
rect 27244 10558 27246 10610
rect 27298 10558 27300 10610
rect 25116 9874 25172 9884
rect 25340 10052 25396 10062
rect 24332 6130 24388 9548
rect 25340 9042 25396 9996
rect 25340 8990 25342 9042
rect 25394 8990 25396 9042
rect 25340 8978 25396 8990
rect 26124 9938 26180 10108
rect 27244 10052 27300 10558
rect 27244 9986 27300 9996
rect 26124 9886 26126 9938
rect 26178 9886 26180 9938
rect 26012 8932 26068 8942
rect 26012 8838 26068 8876
rect 26124 8372 26180 9886
rect 27356 8428 27412 14140
rect 27580 13860 27636 14254
rect 27804 14196 27860 14206
rect 27692 13860 27748 13870
rect 27580 13858 27748 13860
rect 27580 13806 27694 13858
rect 27746 13806 27748 13858
rect 27580 13804 27748 13806
rect 27692 13794 27748 13804
rect 27468 13412 27524 13422
rect 27468 12962 27524 13356
rect 27468 12910 27470 12962
rect 27522 12910 27524 12962
rect 27468 12898 27524 12910
rect 27804 12962 27860 14140
rect 27804 12910 27806 12962
rect 27858 12910 27860 12962
rect 27804 12898 27860 12910
rect 27468 12738 27524 12750
rect 27468 12686 27470 12738
rect 27522 12686 27524 12738
rect 27468 11620 27524 12686
rect 27468 11564 27972 11620
rect 27916 10722 27972 11564
rect 27916 10670 27918 10722
rect 27970 10670 27972 10722
rect 27916 10658 27972 10670
rect 27916 9940 27972 9950
rect 28028 9940 28084 14588
rect 28140 14308 28196 15260
rect 28140 12852 28196 14252
rect 28252 14420 28308 14430
rect 28588 14420 28644 15262
rect 28700 14756 28756 15374
rect 28700 14690 28756 14700
rect 29372 15314 29428 15326
rect 29372 15262 29374 15314
rect 29426 15262 29428 15314
rect 28252 14418 28644 14420
rect 28252 14366 28254 14418
rect 28306 14366 28644 14418
rect 28252 14364 28644 14366
rect 28252 14084 28308 14364
rect 29260 14308 29316 14318
rect 29260 14214 29316 14252
rect 28252 14018 28308 14028
rect 28140 12786 28196 12796
rect 29372 13748 29428 15262
rect 29708 14756 29764 15484
rect 30044 15428 30100 15820
rect 30156 15652 30212 22876
rect 30268 21028 30324 26852
rect 31388 26516 31444 31892
rect 31500 31556 31556 31566
rect 31500 31108 31556 31500
rect 31836 31218 31892 38668
rect 31948 37828 32004 38782
rect 33068 38834 33124 38846
rect 33068 38782 33070 38834
rect 33122 38782 33124 38834
rect 31948 37762 32004 37772
rect 32396 37940 32452 37950
rect 31948 34580 32004 34590
rect 31948 34130 32004 34524
rect 31948 34078 31950 34130
rect 32002 34078 32004 34130
rect 31948 34020 32004 34078
rect 31948 33954 32004 33964
rect 31836 31166 31838 31218
rect 31890 31166 31892 31218
rect 31836 31154 31892 31166
rect 32060 31890 32116 31902
rect 32060 31838 32062 31890
rect 32114 31838 32116 31890
rect 32060 31108 32116 31838
rect 32284 31108 32340 31118
rect 32060 31052 32284 31108
rect 31500 30994 31556 31052
rect 32284 31014 32340 31052
rect 31500 30942 31502 30994
rect 31554 30942 31556 30994
rect 31500 30930 31556 30942
rect 31948 30100 32004 30110
rect 31948 30006 32004 30044
rect 31836 28644 31892 28654
rect 31500 28418 31556 28430
rect 31500 28366 31502 28418
rect 31554 28366 31556 28418
rect 31500 27972 31556 28366
rect 31500 27906 31556 27916
rect 31388 26450 31444 26460
rect 31500 26962 31556 26974
rect 31500 26910 31502 26962
rect 31554 26910 31556 26962
rect 30940 23380 30996 23390
rect 31500 23380 31556 26910
rect 31724 26180 31780 26190
rect 31612 25620 31668 25630
rect 31612 25506 31668 25564
rect 31612 25454 31614 25506
rect 31666 25454 31668 25506
rect 31612 25442 31668 25454
rect 31724 25282 31780 26124
rect 31724 25230 31726 25282
rect 31778 25230 31780 25282
rect 31724 23492 31780 25230
rect 31724 23426 31780 23436
rect 30940 23378 31556 23380
rect 30940 23326 30942 23378
rect 30994 23326 31556 23378
rect 30940 23324 31556 23326
rect 30940 23314 30996 23324
rect 30380 23268 30436 23278
rect 30380 22372 30436 23212
rect 30380 22306 30436 22316
rect 30492 23154 30548 23166
rect 30492 23102 30494 23154
rect 30546 23102 30548 23154
rect 30492 22708 30548 23102
rect 30716 23154 30772 23166
rect 30716 23102 30718 23154
rect 30770 23102 30772 23154
rect 30716 23044 30772 23102
rect 30716 22978 30772 22988
rect 31388 23044 31444 23054
rect 31836 23044 31892 28588
rect 32172 25620 32228 25630
rect 32172 24612 32228 25564
rect 32396 25508 32452 37884
rect 32508 34356 32564 34366
rect 32508 34262 32564 34300
rect 33068 31780 33124 38782
rect 34972 38724 35028 39454
rect 35084 39060 35140 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35980 41188 36036 41198
rect 35980 41094 36036 41132
rect 36316 41188 36372 41198
rect 35980 40404 36036 40414
rect 35980 40310 36036 40348
rect 35644 40292 35700 40302
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35308 39620 35364 39630
rect 35308 39506 35364 39564
rect 35308 39454 35310 39506
rect 35362 39454 35364 39506
rect 35308 39442 35364 39454
rect 35196 39060 35252 39070
rect 35084 39004 35196 39060
rect 35196 38994 35252 39004
rect 35644 38834 35700 40236
rect 35644 38782 35646 38834
rect 35698 38782 35700 38834
rect 35644 38770 35700 38782
rect 35980 39506 36036 39518
rect 35980 39454 35982 39506
rect 36034 39454 36036 39506
rect 34972 38658 35028 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 33180 34020 33236 34030
rect 33180 31948 33236 33964
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35980 31948 36036 39454
rect 36316 39506 36372 41132
rect 36428 39844 36484 41804
rect 36988 41410 37044 41916
rect 36988 41358 36990 41410
rect 37042 41358 37044 41410
rect 36988 41346 37044 41358
rect 37436 41412 37492 44200
rect 37436 41346 37492 41356
rect 36988 41076 37044 41086
rect 36988 40626 37044 41020
rect 36988 40574 36990 40626
rect 37042 40574 37044 40626
rect 36988 40562 37044 40574
rect 36428 39778 36484 39788
rect 37996 39844 38052 39854
rect 37996 39750 38052 39788
rect 38556 39844 38612 44200
rect 38556 39778 38612 39788
rect 36988 39620 37044 39630
rect 36988 39526 37044 39564
rect 37324 39620 37380 39630
rect 36316 39454 36318 39506
rect 36370 39454 36372 39506
rect 36316 39442 36372 39454
rect 36428 39060 36484 39070
rect 36428 38966 36484 39004
rect 33180 31892 33460 31948
rect 33068 31714 33124 31724
rect 32732 29988 32788 29998
rect 32732 28756 32788 29932
rect 32732 28642 32788 28700
rect 32732 28590 32734 28642
rect 32786 28590 32788 28642
rect 32732 28578 32788 28590
rect 32844 28644 32900 28654
rect 32844 28550 32900 28588
rect 33292 28418 33348 28430
rect 33292 28366 33294 28418
rect 33346 28366 33348 28418
rect 33068 27860 33124 27870
rect 33292 27860 33348 28366
rect 33124 27804 33348 27860
rect 33068 27766 33124 27804
rect 33292 26964 33348 27804
rect 32396 25442 32452 25452
rect 33180 26852 33348 26908
rect 33180 24946 33236 26852
rect 33180 24894 33182 24946
rect 33234 24894 33236 24946
rect 32284 24612 32340 24622
rect 32172 24610 32340 24612
rect 32172 24558 32286 24610
rect 32338 24558 32340 24610
rect 32172 24556 32340 24558
rect 32284 24546 32340 24556
rect 32956 24052 33012 24062
rect 33180 24052 33236 24894
rect 33404 24164 33460 31892
rect 35868 31892 36036 31948
rect 34972 31556 35028 31566
rect 34076 30322 34132 30334
rect 34076 30270 34078 30322
rect 34130 30270 34132 30322
rect 34076 30212 34132 30270
rect 34636 30322 34692 30334
rect 34636 30270 34638 30322
rect 34690 30270 34692 30322
rect 34076 29652 34132 30156
rect 34076 29586 34132 29596
rect 34412 30210 34468 30222
rect 34412 30158 34414 30210
rect 34466 30158 34468 30210
rect 34076 29316 34132 29326
rect 34412 29316 34468 30158
rect 34636 30212 34692 30270
rect 34636 30146 34692 30156
rect 34972 30210 35028 31500
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34972 30158 34974 30210
rect 35026 30158 35028 30210
rect 34972 30146 35028 30158
rect 34076 29314 34468 29316
rect 34076 29262 34078 29314
rect 34130 29262 34468 29314
rect 34076 29260 34468 29262
rect 33740 28756 33796 28766
rect 33628 28700 33740 28756
rect 33628 27186 33684 28700
rect 33740 28662 33796 28700
rect 34076 28644 34132 29260
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34076 28578 34132 28588
rect 33852 28420 33908 28430
rect 33852 27970 33908 28364
rect 33852 27918 33854 27970
rect 33906 27918 33908 27970
rect 33852 27906 33908 27918
rect 34412 27972 34468 27982
rect 33628 27134 33630 27186
rect 33682 27134 33684 27186
rect 33628 27122 33684 27134
rect 34412 27298 34468 27916
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34412 27246 34414 27298
rect 34466 27246 34468 27298
rect 34412 27188 34468 27246
rect 34748 27300 34804 27310
rect 34748 27206 34804 27244
rect 35868 27300 35924 31892
rect 37324 31666 37380 39564
rect 38332 39396 38388 39406
rect 38332 38946 38388 39340
rect 38332 38894 38334 38946
rect 38386 38894 38388 38946
rect 38332 38882 38388 38894
rect 38668 38946 38724 38958
rect 38668 38894 38670 38946
rect 38722 38894 38724 38946
rect 38668 38052 38724 38894
rect 39116 38948 39172 38958
rect 39116 38854 39172 38892
rect 39452 38946 39508 38958
rect 39452 38894 39454 38946
rect 39506 38894 39508 38946
rect 38892 38052 38948 38062
rect 38668 37996 38892 38052
rect 38892 37986 38948 37996
rect 39452 37716 39508 38894
rect 39676 38276 39732 44200
rect 40796 44100 40852 44200
rect 41132 44100 41188 44268
rect 40796 44044 41188 44100
rect 40796 41412 40852 41422
rect 40796 41318 40852 41356
rect 39788 41188 39844 41198
rect 39788 41094 39844 41132
rect 40908 39844 40964 39854
rect 40908 39750 40964 39788
rect 39900 39620 39956 39630
rect 39900 39526 39956 39564
rect 39676 38210 39732 38220
rect 40908 38276 40964 38286
rect 40908 38182 40964 38220
rect 39900 38052 39956 38062
rect 39900 37958 39956 37996
rect 39452 37650 39508 37660
rect 40572 37716 40628 37726
rect 40572 36482 40628 37660
rect 41580 36706 41636 44268
rect 43148 41074 43204 41086
rect 43148 41022 43150 41074
rect 43202 41022 43204 41074
rect 42812 40964 42868 40974
rect 42812 40870 42868 40908
rect 43148 40404 43204 41022
rect 43148 40310 43204 40348
rect 41580 36654 41582 36706
rect 41634 36654 41636 36706
rect 41580 36642 41636 36654
rect 40572 36430 40574 36482
rect 40626 36430 40628 36482
rect 40572 36418 40628 36430
rect 42812 33908 42868 33918
rect 39452 33460 39508 33470
rect 37324 31614 37326 31666
rect 37378 31614 37380 31666
rect 37324 31602 37380 31614
rect 37772 33012 37828 33022
rect 36988 31556 37044 31566
rect 36988 31462 37044 31500
rect 35868 27234 35924 27244
rect 35980 27746 36036 27758
rect 35980 27694 35982 27746
rect 36034 27694 36036 27746
rect 34412 27122 34468 27132
rect 35196 27188 35252 27198
rect 35196 27094 35252 27132
rect 35980 27188 36036 27694
rect 35980 27122 36036 27132
rect 34188 27074 34244 27086
rect 34188 27022 34190 27074
rect 34242 27022 34244 27074
rect 34188 26908 34244 27022
rect 33964 26852 34020 26862
rect 34188 26852 34468 26908
rect 34020 26796 34132 26852
rect 33964 26786 34020 26796
rect 34076 26628 34132 26796
rect 34076 26572 34356 26628
rect 34300 26514 34356 26572
rect 34300 26462 34302 26514
rect 34354 26462 34356 26514
rect 34300 26450 34356 26462
rect 33852 26180 33908 26190
rect 33852 26086 33908 26124
rect 34412 26180 34468 26852
rect 34412 26114 34468 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 33852 25282 33908 25294
rect 33852 25230 33854 25282
rect 33906 25230 33908 25282
rect 33404 24098 33460 24108
rect 33628 24610 33684 24622
rect 33628 24558 33630 24610
rect 33682 24558 33684 24610
rect 33628 24498 33684 24558
rect 33628 24446 33630 24498
rect 33682 24446 33684 24498
rect 32508 24050 33236 24052
rect 32508 23998 32958 24050
rect 33010 23998 33236 24050
rect 32508 23996 33236 23998
rect 32508 23378 32564 23996
rect 32956 23986 33012 23996
rect 33180 23940 33236 23996
rect 33292 23940 33348 23950
rect 33180 23938 33460 23940
rect 33180 23886 33294 23938
rect 33346 23886 33460 23938
rect 33180 23884 33460 23886
rect 33292 23874 33348 23884
rect 32844 23828 32900 23838
rect 32508 23326 32510 23378
rect 32562 23326 32564 23378
rect 32508 23314 32564 23326
rect 32620 23772 32844 23828
rect 31388 23042 31892 23044
rect 31388 22990 31390 23042
rect 31442 22990 31892 23042
rect 31388 22988 31892 22990
rect 30604 22932 30660 22942
rect 30604 22838 30660 22876
rect 31388 22708 31444 22988
rect 30492 22652 31444 22708
rect 30380 22148 30436 22158
rect 30380 22054 30436 22092
rect 30268 20962 30324 20972
rect 30380 20916 30436 20926
rect 30268 20804 30324 20814
rect 30268 20710 30324 20748
rect 30380 20580 30436 20860
rect 30268 20524 30436 20580
rect 30268 20130 30324 20524
rect 30380 20244 30436 20254
rect 30380 20150 30436 20188
rect 30268 20078 30270 20130
rect 30322 20078 30324 20130
rect 30268 20066 30324 20078
rect 30268 17108 30324 17118
rect 30268 16098 30324 17052
rect 30268 16046 30270 16098
rect 30322 16046 30324 16098
rect 30268 16034 30324 16046
rect 30156 15596 30324 15652
rect 30156 15428 30212 15438
rect 30044 15426 30212 15428
rect 30044 15374 30158 15426
rect 30210 15374 30212 15426
rect 30044 15372 30212 15374
rect 30156 15362 30212 15372
rect 30268 15204 30324 15596
rect 29708 14642 29764 14700
rect 29708 14590 29710 14642
rect 29762 14590 29764 14642
rect 29708 14578 29764 14590
rect 30156 15148 30324 15204
rect 30380 15204 30436 15214
rect 29372 12290 29428 13692
rect 29820 14308 29876 14318
rect 29820 13634 29876 14252
rect 29820 13582 29822 13634
rect 29874 13582 29876 13634
rect 29820 13570 29876 13582
rect 30156 13860 30212 15148
rect 29372 12238 29374 12290
rect 29426 12238 29428 12290
rect 28476 11732 28532 11742
rect 29372 11732 29428 12238
rect 28532 11676 28644 11732
rect 28476 11666 28532 11676
rect 27916 9938 28308 9940
rect 27916 9886 27918 9938
rect 27970 9886 28308 9938
rect 27916 9884 28308 9886
rect 27916 9874 27972 9884
rect 28140 9716 28196 9726
rect 28140 8930 28196 9660
rect 28252 9714 28308 9884
rect 28252 9662 28254 9714
rect 28306 9662 28308 9714
rect 28252 9650 28308 9662
rect 28140 8878 28142 8930
rect 28194 8878 28196 8930
rect 28140 8866 28196 8878
rect 28476 9602 28532 9614
rect 28476 9550 28478 9602
rect 28530 9550 28532 9602
rect 27356 8372 27636 8428
rect 26124 8306 26180 8316
rect 24332 6078 24334 6130
rect 24386 6078 24388 6130
rect 24332 6066 24388 6078
rect 24220 5170 24276 5180
rect 23884 4564 23940 4574
rect 23884 4470 23940 4508
rect 22988 4340 23044 4350
rect 22988 4246 23044 4284
rect 26460 4114 26516 4126
rect 26460 4062 26462 4114
rect 26514 4062 26516 4114
rect 21420 3502 21422 3554
rect 21474 3502 21476 3554
rect 21420 3490 21476 3502
rect 24780 3666 24836 3678
rect 24780 3614 24782 3666
rect 24834 3614 24836 3666
rect 20636 3332 21140 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20636 800 20692 3332
rect 22428 3330 22484 3342
rect 22428 3278 22430 3330
rect 22482 3278 22484 3330
rect 22428 800 22484 3278
rect 24220 924 24500 980
rect 24220 800 24276 924
rect 2688 0 2800 800
rect 4480 0 4592 800
rect 6272 0 6384 800
rect 8064 0 8176 800
rect 9856 0 9968 800
rect 11648 0 11760 800
rect 13440 0 13552 800
rect 15232 0 15344 800
rect 17024 0 17136 800
rect 18816 0 18928 800
rect 20608 0 20720 800
rect 22400 0 22512 800
rect 24192 0 24304 800
rect 24444 756 24500 924
rect 24780 756 24836 3614
rect 26460 3388 26516 4062
rect 27580 3668 27636 8372
rect 27132 3666 27636 3668
rect 27132 3614 27582 3666
rect 27634 3614 27636 3666
rect 27132 3612 27636 3614
rect 27132 3554 27188 3612
rect 27580 3602 27636 3612
rect 27804 3668 27860 3678
rect 27132 3502 27134 3554
rect 27186 3502 27188 3554
rect 27132 3490 27188 3502
rect 26012 3332 26516 3388
rect 26012 800 26068 3332
rect 27804 800 27860 3612
rect 28476 3554 28532 9550
rect 28588 9042 28644 11676
rect 29372 11666 29428 11676
rect 30156 10836 30212 13804
rect 30156 10742 30212 10780
rect 29148 10500 29204 10510
rect 29148 9156 29204 10444
rect 29708 9940 29764 9950
rect 29260 9828 29316 9838
rect 29260 9734 29316 9772
rect 29596 9714 29652 9726
rect 29596 9662 29598 9714
rect 29650 9662 29652 9714
rect 29596 9604 29652 9662
rect 29708 9714 29764 9884
rect 29708 9662 29710 9714
rect 29762 9662 29764 9714
rect 29708 9650 29764 9662
rect 29260 9156 29316 9166
rect 29148 9154 29316 9156
rect 29148 9102 29262 9154
rect 29314 9102 29316 9154
rect 29148 9100 29316 9102
rect 29260 9090 29316 9100
rect 28588 8990 28590 9042
rect 28642 8990 28644 9042
rect 28588 8978 28644 8990
rect 29596 9044 29652 9548
rect 29596 8978 29652 8988
rect 29932 9602 29988 9614
rect 29932 9550 29934 9602
rect 29986 9550 29988 9602
rect 28812 4340 28868 4350
rect 28812 4246 28868 4284
rect 29932 4338 29988 9550
rect 30268 9604 30324 9614
rect 30268 9510 30324 9548
rect 29932 4286 29934 4338
rect 29986 4286 29988 4338
rect 29932 4274 29988 4286
rect 30380 4340 30436 15148
rect 30492 15148 30548 22652
rect 30940 22372 30996 22382
rect 30716 20916 30772 20926
rect 30716 20130 30772 20860
rect 30940 20916 30996 22316
rect 31836 21474 31892 21486
rect 31836 21422 31838 21474
rect 31890 21422 31892 21474
rect 30940 20822 30996 20860
rect 31276 21252 31332 21262
rect 31276 20242 31332 21196
rect 31836 21252 31892 21422
rect 31836 21028 31892 21196
rect 32172 21028 32228 21038
rect 31836 21026 32228 21028
rect 31836 20974 31838 21026
rect 31890 20974 32174 21026
rect 32226 20974 32228 21026
rect 31836 20972 32228 20974
rect 31836 20962 31892 20972
rect 32172 20962 32228 20972
rect 31500 20916 31556 20926
rect 31276 20190 31278 20242
rect 31330 20190 31332 20242
rect 31276 20178 31332 20190
rect 31388 20914 31556 20916
rect 31388 20862 31502 20914
rect 31554 20862 31556 20914
rect 31388 20860 31556 20862
rect 30716 20078 30718 20130
rect 30770 20078 30772 20130
rect 30716 20066 30772 20078
rect 30828 18564 30884 18574
rect 30828 18450 30884 18508
rect 30828 18398 30830 18450
rect 30882 18398 30884 18450
rect 30828 18386 30884 18398
rect 30828 17780 30884 17790
rect 30828 17666 30884 17724
rect 30828 17614 30830 17666
rect 30882 17614 30884 17666
rect 30828 17602 30884 17614
rect 31388 17556 31444 20860
rect 31500 20850 31556 20860
rect 31612 20916 31668 20926
rect 31612 20690 31668 20860
rect 31612 20638 31614 20690
rect 31666 20638 31668 20690
rect 31612 20626 31668 20638
rect 32284 20578 32340 20590
rect 32284 20526 32286 20578
rect 32338 20526 32340 20578
rect 32284 20244 32340 20526
rect 32060 20188 32340 20244
rect 32396 20578 32452 20590
rect 32396 20526 32398 20578
rect 32450 20526 32452 20578
rect 32060 20130 32116 20188
rect 32060 20078 32062 20130
rect 32114 20078 32116 20130
rect 32060 20066 32116 20078
rect 31500 20018 31556 20030
rect 31500 19966 31502 20018
rect 31554 19966 31556 20018
rect 31500 19908 31556 19966
rect 31724 20020 31780 20030
rect 31724 19926 31780 19964
rect 31500 19842 31556 19852
rect 31612 19906 31668 19918
rect 31612 19854 31614 19906
rect 31666 19854 31668 19906
rect 31612 18564 31668 19854
rect 31612 18498 31668 18508
rect 32060 19122 32116 19134
rect 32060 19070 32062 19122
rect 32114 19070 32116 19122
rect 31500 18450 31556 18462
rect 31500 18398 31502 18450
rect 31554 18398 31556 18450
rect 31500 18340 31556 18398
rect 32060 18452 32116 19070
rect 32396 19124 32452 20526
rect 32508 20020 32564 20030
rect 32508 19236 32564 19964
rect 32508 19170 32564 19180
rect 32396 19058 32452 19068
rect 32620 18900 32676 23772
rect 32844 23762 32900 23772
rect 33292 23604 33348 23614
rect 33068 23380 33124 23390
rect 33068 23156 33124 23324
rect 33292 23378 33348 23548
rect 33292 23326 33294 23378
rect 33346 23326 33348 23378
rect 33292 23314 33348 23326
rect 33404 23156 33460 23884
rect 33628 23268 33684 24446
rect 33852 24500 33908 25230
rect 34300 24834 34356 24846
rect 34300 24782 34302 24834
rect 34354 24782 34356 24834
rect 33964 24724 34020 24734
rect 34300 24724 34356 24782
rect 33964 24722 34356 24724
rect 33964 24670 33966 24722
rect 34018 24670 34356 24722
rect 33964 24668 34356 24670
rect 33964 24658 34020 24668
rect 34076 24500 34132 24510
rect 33852 24498 34132 24500
rect 33852 24446 34078 24498
rect 34130 24446 34132 24498
rect 33852 24444 34132 24446
rect 33852 23716 33908 23726
rect 33964 23716 34020 24444
rect 34076 24434 34132 24444
rect 34412 24498 34468 24510
rect 34412 24446 34414 24498
rect 34466 24446 34468 24498
rect 33908 23660 34020 23716
rect 34076 23826 34132 23838
rect 34076 23774 34078 23826
rect 34130 23774 34132 23826
rect 33852 23650 33908 23660
rect 34076 23604 34132 23774
rect 34076 23538 34132 23548
rect 33628 23202 33684 23212
rect 33852 23492 33908 23502
rect 33068 23154 33348 23156
rect 33068 23102 33070 23154
rect 33122 23102 33348 23154
rect 33068 23100 33348 23102
rect 33404 23100 33572 23156
rect 33068 23090 33124 23100
rect 32956 20578 33012 20590
rect 32956 20526 32958 20578
rect 33010 20526 33012 20578
rect 32956 20020 33012 20526
rect 33180 20020 33236 20030
rect 32956 20018 33236 20020
rect 32956 19966 33182 20018
rect 33234 19966 33236 20018
rect 32956 19964 33236 19966
rect 32060 18340 32116 18396
rect 31500 18338 32116 18340
rect 31500 18286 32062 18338
rect 32114 18286 32116 18338
rect 31500 18284 32116 18286
rect 31500 17780 31556 18284
rect 31500 17714 31556 17724
rect 31612 17556 31668 17566
rect 31388 17554 31668 17556
rect 31388 17502 31614 17554
rect 31666 17502 31668 17554
rect 31388 17500 31668 17502
rect 31612 17490 31668 17500
rect 32060 16098 32116 18284
rect 32060 16046 32062 16098
rect 32114 16046 32116 16098
rect 32060 16034 32116 16046
rect 32396 18844 32676 18900
rect 32396 15540 32452 18844
rect 33180 18452 33236 19964
rect 33180 18386 33236 18396
rect 33292 19012 33348 23100
rect 33516 23044 33572 23100
rect 33740 23154 33796 23166
rect 33740 23102 33742 23154
rect 33794 23102 33796 23154
rect 33740 23044 33796 23102
rect 33516 22988 33796 23044
rect 33404 22932 33460 22942
rect 33404 22930 33796 22932
rect 33404 22878 33406 22930
rect 33458 22878 33796 22930
rect 33404 22876 33796 22878
rect 33404 22866 33460 22876
rect 33740 22482 33796 22876
rect 33740 22430 33742 22482
rect 33794 22430 33796 22482
rect 33740 22418 33796 22430
rect 33852 22372 33908 23436
rect 34412 23268 34468 24446
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 36204 24050 36260 24062
rect 36204 23998 36206 24050
rect 36258 23998 36260 24050
rect 34860 23716 34916 23726
rect 34524 23268 34580 23278
rect 34412 23266 34580 23268
rect 34412 23214 34526 23266
rect 34578 23214 34580 23266
rect 34412 23212 34580 23214
rect 34524 23202 34580 23212
rect 33852 22278 33908 22316
rect 34076 22596 34132 22606
rect 33628 22258 33684 22270
rect 33628 22206 33630 22258
rect 33682 22206 33684 22258
rect 33628 21924 33684 22206
rect 33628 21858 33684 21868
rect 33852 20802 33908 20814
rect 33852 20750 33854 20802
rect 33906 20750 33908 20802
rect 33852 20244 33908 20750
rect 34076 20804 34132 22540
rect 34748 22484 34804 22494
rect 34188 22482 34804 22484
rect 34188 22430 34750 22482
rect 34802 22430 34804 22482
rect 34188 22428 34804 22430
rect 34188 22370 34244 22428
rect 34748 22418 34804 22428
rect 34188 22318 34190 22370
rect 34242 22318 34244 22370
rect 34188 22306 34244 22318
rect 34636 22260 34692 22270
rect 34860 22260 34916 23660
rect 34972 23044 35028 23054
rect 34972 22370 35028 22988
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34972 22318 34974 22370
rect 35026 22318 35028 22370
rect 34972 22306 35028 22318
rect 35420 22372 35476 22382
rect 35420 22278 35476 22316
rect 36204 22372 36260 23998
rect 36652 23044 36708 23054
rect 36652 22950 36708 22988
rect 36260 22316 36708 22372
rect 36204 22306 36260 22316
rect 34412 22258 34916 22260
rect 34412 22206 34638 22258
rect 34690 22206 34916 22258
rect 34412 22204 34916 22206
rect 34412 21810 34468 22204
rect 34636 22194 34692 22204
rect 34412 21758 34414 21810
rect 34466 21758 34468 21810
rect 34412 21746 34468 21758
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 20916 35140 20926
rect 34412 20914 35140 20916
rect 34412 20862 35086 20914
rect 35138 20862 35140 20914
rect 34412 20860 35140 20862
rect 34188 20804 34244 20814
rect 34412 20804 34468 20860
rect 34076 20802 34468 20804
rect 34076 20750 34190 20802
rect 34242 20750 34468 20802
rect 34076 20748 34468 20750
rect 34188 20738 34244 20748
rect 34524 20692 34580 20702
rect 34524 20690 34916 20692
rect 34524 20638 34526 20690
rect 34578 20638 34916 20690
rect 34524 20636 34916 20638
rect 34524 20626 34580 20636
rect 33852 20178 33908 20188
rect 34188 20578 34244 20590
rect 34188 20526 34190 20578
rect 34242 20526 34244 20578
rect 34188 20132 34244 20526
rect 34188 20066 34244 20076
rect 33964 19908 34020 19918
rect 33964 19906 34804 19908
rect 33964 19854 33966 19906
rect 34018 19854 34804 19906
rect 33964 19852 34804 19854
rect 33964 19842 34020 19852
rect 34748 19458 34804 19852
rect 34748 19406 34750 19458
rect 34802 19406 34804 19458
rect 34748 19394 34804 19406
rect 34860 19460 34916 20636
rect 34972 20020 35028 20860
rect 35084 20850 35140 20860
rect 35644 20916 35700 20926
rect 34972 19954 35028 19964
rect 35084 20356 35140 20366
rect 35084 19460 35140 20300
rect 35420 20132 35476 20142
rect 35476 20076 35588 20132
rect 35420 20066 35476 20076
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34860 19394 34916 19404
rect 34972 19458 35140 19460
rect 34972 19406 35086 19458
rect 35138 19406 35140 19458
rect 34972 19404 35140 19406
rect 34972 19348 35028 19404
rect 35084 19394 35140 19404
rect 35420 19460 35476 19470
rect 35532 19460 35588 20076
rect 35420 19458 35588 19460
rect 35420 19406 35422 19458
rect 35474 19406 35588 19458
rect 35420 19404 35588 19406
rect 35420 19394 35476 19404
rect 33068 18340 33124 18350
rect 33068 16770 33124 18284
rect 33292 17108 33348 18956
rect 33740 19124 33796 19134
rect 34860 19124 34916 19134
rect 33740 17778 33796 19068
rect 34748 19122 34916 19124
rect 34748 19070 34862 19122
rect 34914 19070 34916 19122
rect 34748 19068 34916 19070
rect 34748 19012 34804 19068
rect 34860 19058 34916 19068
rect 34748 18946 34804 18956
rect 34972 18788 35028 19292
rect 34524 18732 35028 18788
rect 35084 19236 35140 19246
rect 34524 18674 34580 18732
rect 34524 18622 34526 18674
rect 34578 18622 34580 18674
rect 34524 18610 34580 18622
rect 33740 17726 33742 17778
rect 33794 17726 33796 17778
rect 33740 17714 33796 17726
rect 34188 18452 34244 18462
rect 34188 17778 34244 18396
rect 34972 18452 35028 18462
rect 34972 18358 35028 18396
rect 34188 17726 34190 17778
rect 34242 17726 34244 17778
rect 34188 17714 34244 17726
rect 33292 17014 33348 17052
rect 33068 16718 33070 16770
rect 33122 16718 33124 16770
rect 33068 16706 33124 16718
rect 33180 16770 33236 16782
rect 33180 16718 33182 16770
rect 33234 16718 33236 16770
rect 33180 16324 33236 16718
rect 32844 16268 33236 16324
rect 32844 16210 32900 16268
rect 32844 16158 32846 16210
rect 32898 16158 32900 16210
rect 32844 16146 32900 16158
rect 35084 16210 35140 19180
rect 35644 19236 35700 20860
rect 36092 19906 36148 19918
rect 36092 19854 36094 19906
rect 36146 19854 36148 19906
rect 35756 19348 35812 19358
rect 35756 19346 36036 19348
rect 35756 19294 35758 19346
rect 35810 19294 36036 19346
rect 35756 19292 36036 19294
rect 35756 19282 35812 19292
rect 35644 19122 35700 19180
rect 35644 19070 35646 19122
rect 35698 19070 35700 19122
rect 35644 19058 35700 19070
rect 35980 18564 36036 19292
rect 36092 19234 36148 19854
rect 36540 19906 36596 19918
rect 36540 19854 36542 19906
rect 36594 19854 36596 19906
rect 36204 19460 36260 19470
rect 36204 19346 36260 19404
rect 36204 19294 36206 19346
rect 36258 19294 36260 19346
rect 36204 19282 36260 19294
rect 36428 19348 36484 19358
rect 36540 19348 36596 19854
rect 36484 19292 36596 19348
rect 36428 19254 36484 19292
rect 36092 19182 36094 19234
rect 36146 19182 36148 19234
rect 36092 19170 36148 19182
rect 36092 18564 36148 18574
rect 35980 18562 36148 18564
rect 35980 18510 36094 18562
rect 36146 18510 36148 18562
rect 35980 18508 36148 18510
rect 36092 18498 36148 18508
rect 35420 18452 35476 18462
rect 35476 18396 35700 18452
rect 35420 18358 35476 18396
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35084 16158 35086 16210
rect 35138 16158 35140 16210
rect 32396 15446 32452 15484
rect 35084 15148 35140 16158
rect 35644 16210 35700 18396
rect 35644 16158 35646 16210
rect 35698 16158 35700 16210
rect 35644 16146 35700 16158
rect 30492 15092 30660 15148
rect 35084 15092 35588 15148
rect 30604 9940 30660 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 33404 13524 33460 13534
rect 32732 13076 32788 13086
rect 30716 9940 30772 9950
rect 30660 9938 30772 9940
rect 30660 9886 30718 9938
rect 30770 9886 30772 9938
rect 30660 9884 30772 9886
rect 30604 9846 30660 9884
rect 30716 9874 30772 9884
rect 31388 9604 31444 9614
rect 31388 8930 31444 9548
rect 31388 8878 31390 8930
rect 31442 8878 31444 8930
rect 31388 8866 31444 8878
rect 30380 4274 30436 4284
rect 29596 4116 29652 4126
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 28476 3502 28478 3554
rect 28530 3502 28532 3554
rect 28476 3490 28532 3502
rect 29596 800 29652 4060
rect 30828 4116 30884 4126
rect 30828 4022 30884 4060
rect 32732 3666 32788 13020
rect 32732 3614 32734 3666
rect 32786 3614 32788 3666
rect 32732 3602 32788 3614
rect 33292 4226 33348 4238
rect 33292 4174 33294 4226
rect 33346 4174 33348 4226
rect 31724 3444 31780 3454
rect 32172 3444 32228 3454
rect 31388 3442 32228 3444
rect 31388 3390 31726 3442
rect 31778 3390 32174 3442
rect 32226 3390 32228 3442
rect 31388 3388 32228 3390
rect 31388 800 31444 3388
rect 31724 3350 31780 3388
rect 32172 3378 32228 3388
rect 33292 2548 33348 4174
rect 33404 3442 33460 13468
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35084 7588 35140 7598
rect 35084 4340 35140 7532
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35084 4274 35140 4284
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34972 3668 35028 3678
rect 33628 3556 33684 3566
rect 33404 3390 33406 3442
rect 33458 3390 33460 3442
rect 33404 3378 33460 3390
rect 33516 3554 33684 3556
rect 33516 3502 33630 3554
rect 33682 3502 33684 3554
rect 33516 3500 33684 3502
rect 33516 2548 33572 3500
rect 33628 3490 33684 3500
rect 33180 2492 33572 2548
rect 33180 800 33236 2492
rect 34972 800 35028 3612
rect 35532 3668 35588 15092
rect 36652 4564 36708 22316
rect 37100 19236 37156 19246
rect 37100 19142 37156 19180
rect 37772 6692 37828 32956
rect 38220 20020 38276 20030
rect 38276 19964 38388 20020
rect 38220 19954 38276 19964
rect 38332 18676 38388 19964
rect 38332 18582 38388 18620
rect 37772 6626 37828 6636
rect 39340 18564 39396 18574
rect 36652 4562 37044 4564
rect 36652 4510 36654 4562
rect 36706 4510 37044 4562
rect 36652 4508 37044 4510
rect 36652 4498 36708 4508
rect 36988 4338 37044 4508
rect 36988 4286 36990 4338
rect 37042 4286 37044 4338
rect 36988 4274 37044 4286
rect 36764 4116 36820 4126
rect 35532 3666 36036 3668
rect 35532 3614 35534 3666
rect 35586 3614 36036 3666
rect 35532 3612 36036 3614
rect 35532 3602 35588 3612
rect 35980 3554 36036 3612
rect 35980 3502 35982 3554
rect 36034 3502 36036 3554
rect 35980 3490 36036 3502
rect 36764 800 36820 4060
rect 37996 4116 38052 4126
rect 37996 4022 38052 4060
rect 36988 3668 37044 3678
rect 36988 3574 37044 3612
rect 38556 3668 38612 3678
rect 38556 800 38612 3612
rect 39340 3668 39396 18508
rect 39452 13972 39508 33404
rect 41132 32900 41188 32910
rect 41132 23380 41188 32844
rect 42812 31666 42868 33852
rect 42812 31614 42814 31666
rect 42866 31614 42868 31666
rect 42812 31602 42868 31614
rect 43148 31666 43204 31678
rect 43148 31614 43150 31666
rect 43202 31614 43204 31666
rect 42588 31554 42644 31566
rect 42588 31502 42590 31554
rect 42642 31502 42644 31554
rect 42588 31444 42644 31502
rect 42588 31378 42644 31388
rect 43148 31444 43204 31614
rect 43148 31378 43204 31388
rect 41132 23314 41188 23324
rect 42812 23380 42868 23390
rect 42812 23286 42868 23324
rect 43148 23154 43204 23166
rect 43148 23102 43150 23154
rect 43202 23102 43204 23154
rect 42588 23044 42644 23054
rect 43148 23044 43204 23102
rect 42588 23042 43204 23044
rect 42588 22990 42590 23042
rect 42642 22990 43204 23042
rect 42588 22988 43204 22990
rect 42588 22978 42644 22988
rect 43148 22484 43204 22988
rect 43148 22418 43204 22428
rect 39452 13906 39508 13916
rect 40348 20580 40404 20590
rect 39340 3666 39844 3668
rect 39340 3614 39342 3666
rect 39394 3614 39844 3666
rect 39340 3612 39844 3614
rect 39340 3602 39396 3612
rect 39788 3554 39844 3612
rect 39788 3502 39790 3554
rect 39842 3502 39844 3554
rect 39788 3490 39844 3502
rect 40348 800 40404 20524
rect 42812 13972 42868 13982
rect 42812 13878 42868 13916
rect 43148 13746 43204 13758
rect 43148 13694 43150 13746
rect 43202 13694 43204 13746
rect 42588 13634 42644 13646
rect 42588 13582 42590 13634
rect 42642 13582 42644 13634
rect 42588 13524 42644 13582
rect 42588 13458 42644 13468
rect 43148 13524 43204 13694
rect 43148 13458 43204 13468
rect 42812 6692 42868 6702
rect 42588 5124 42644 5134
rect 42588 5030 42644 5068
rect 42812 5010 42868 6636
rect 42812 4958 42814 5010
rect 42866 4958 42868 5010
rect 42812 4946 42868 4958
rect 43148 5124 43204 5134
rect 43148 4564 43204 5068
rect 43148 4498 43204 4508
rect 42364 4338 42420 4350
rect 42364 4286 42366 4338
rect 42418 4286 42420 4338
rect 42140 4228 42196 4238
rect 42364 4228 42420 4286
rect 42140 4226 42420 4228
rect 42140 4174 42142 4226
rect 42194 4174 42420 4226
rect 42140 4172 42420 4174
rect 42812 4340 42868 4350
rect 42812 4226 42868 4284
rect 42812 4174 42814 4226
rect 42866 4174 42868 4226
rect 40796 3668 40852 3678
rect 40796 3574 40852 3612
rect 42140 800 42196 4172
rect 42812 4162 42868 4174
rect 24444 700 24836 756
rect 25984 0 26096 800
rect 27776 0 27888 800
rect 29568 0 29680 800
rect 31360 0 31472 800
rect 33152 0 33264 800
rect 34944 0 35056 800
rect 36736 0 36848 800
rect 38528 0 38640 800
rect 40320 0 40432 800
rect 42112 0 42224 800
<< via2 >>
rect 1932 40572 1988 40628
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4732 41244 4788 41300
rect 5404 41916 5460 41972
rect 4284 41020 4340 41076
rect 4396 40908 4452 40964
rect 3836 39676 3892 39732
rect 4172 40684 4228 40740
rect 1932 39564 1988 39620
rect 1932 38834 1988 38836
rect 1932 38782 1934 38834
rect 1934 38782 1986 38834
rect 1986 38782 1988 38834
rect 1932 38780 1988 38782
rect 1372 38668 1428 38724
rect 1260 30044 1316 30100
rect 1932 38162 1988 38164
rect 1932 38110 1934 38162
rect 1934 38110 1986 38162
rect 1986 38110 1988 38162
rect 1932 38108 1988 38110
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 1932 36540 1988 36596
rect 1596 35532 1652 35588
rect 1484 34972 1540 35028
rect 1484 29596 1540 29652
rect 1372 21868 1428 21924
rect 1260 13020 1316 13076
rect 2044 35196 2100 35252
rect 2044 34748 2100 34804
rect 2156 34130 2212 34132
rect 2156 34078 2158 34130
rect 2158 34078 2210 34130
rect 2210 34078 2212 34130
rect 2156 34076 2212 34078
rect 1932 33852 1988 33908
rect 2268 33852 2324 33908
rect 2044 33404 2100 33460
rect 2940 36540 2996 36596
rect 4060 37772 4116 37828
rect 4284 38892 4340 38948
rect 4732 38556 4788 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 5628 41298 5684 41300
rect 5628 41246 5630 41298
rect 5630 41246 5682 41298
rect 5682 41246 5684 41298
rect 5628 41244 5684 41246
rect 7644 40962 7700 40964
rect 7644 40910 7646 40962
rect 7646 40910 7698 40962
rect 7698 40910 7700 40962
rect 7644 40908 7700 40910
rect 7868 40684 7924 40740
rect 8204 40684 8260 40740
rect 4956 40348 5012 40404
rect 5964 40348 6020 40404
rect 5180 38834 5236 38836
rect 5180 38782 5182 38834
rect 5182 38782 5234 38834
rect 5234 38782 5236 38834
rect 5180 38780 5236 38782
rect 5740 38780 5796 38836
rect 4844 38050 4900 38052
rect 4844 37998 4846 38050
rect 4846 37998 4898 38050
rect 4898 37998 4900 38050
rect 4844 37996 4900 37998
rect 5740 38050 5796 38052
rect 5740 37998 5742 38050
rect 5742 37998 5794 38050
rect 5794 37998 5796 38050
rect 5740 37996 5796 37998
rect 4284 37324 4340 37380
rect 4956 37212 5012 37268
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 5068 36876 5124 36932
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4060 34748 4116 34804
rect 2604 34076 2660 34132
rect 2492 33404 2548 33460
rect 1932 32508 1988 32564
rect 1932 31164 1988 31220
rect 1932 30322 1988 30324
rect 1932 30270 1934 30322
rect 1934 30270 1986 30322
rect 1986 30270 1988 30322
rect 1932 30268 1988 30270
rect 1820 29820 1876 29876
rect 2044 29650 2100 29652
rect 2044 29598 2046 29650
rect 2046 29598 2098 29650
rect 2098 29598 2100 29650
rect 2044 29596 2100 29598
rect 3052 32956 3108 33012
rect 3612 32844 3668 32900
rect 4620 33852 4676 33908
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4284 33516 4340 33572
rect 4620 33346 4676 33348
rect 4620 33294 4622 33346
rect 4622 33294 4674 33346
rect 4674 33294 4676 33346
rect 4620 33292 4676 33294
rect 4284 33180 4340 33236
rect 4732 32844 4788 32900
rect 4172 32620 4228 32676
rect 2604 31388 2660 31444
rect 2604 30268 2660 30324
rect 2716 29596 2772 29652
rect 1932 28476 1988 28532
rect 1932 27132 1988 27188
rect 2044 25788 2100 25844
rect 1708 25618 1764 25620
rect 1708 25566 1710 25618
rect 1710 25566 1762 25618
rect 1762 25566 1764 25618
rect 1708 25564 1764 25566
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 1708 23548 1764 23604
rect 1932 23100 1988 23156
rect 1932 21756 1988 21812
rect 1708 20972 1764 21028
rect 1932 20412 1988 20468
rect 1932 19346 1988 19348
rect 1932 19294 1934 19346
rect 1934 19294 1986 19346
rect 1986 19294 1988 19346
rect 1932 19292 1988 19294
rect 1708 18450 1764 18452
rect 1708 18398 1710 18450
rect 1710 18398 1762 18450
rect 1762 18398 1764 18450
rect 1708 18396 1764 18398
rect 2044 18172 2100 18228
rect 2380 18284 2436 18340
rect 1708 17724 1764 17780
rect 1932 17778 1988 17780
rect 1932 17726 1934 17778
rect 1934 17726 1986 17778
rect 1986 17726 1988 17778
rect 1932 17724 1988 17726
rect 2268 17500 2324 17556
rect 2268 16828 2324 16884
rect 2156 16716 2212 16772
rect 1932 16044 1988 16100
rect 1708 15036 1764 15092
rect 1708 13970 1764 13972
rect 1708 13918 1710 13970
rect 1710 13918 1762 13970
rect 1762 13918 1764 13970
rect 1708 13916 1764 13918
rect 2380 16380 2436 16436
rect 1932 15036 1988 15092
rect 3276 29596 3332 29652
rect 3052 27244 3108 27300
rect 2716 21756 2772 21812
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 5068 35922 5124 35924
rect 5068 35870 5070 35922
rect 5070 35870 5122 35922
rect 5122 35870 5124 35922
rect 5068 35868 5124 35870
rect 4956 34860 5012 34916
rect 5852 37436 5908 37492
rect 7196 40402 7252 40404
rect 7196 40350 7198 40402
rect 7198 40350 7250 40402
rect 7250 40350 7252 40402
rect 7196 40348 7252 40350
rect 7196 39730 7252 39732
rect 7196 39678 7198 39730
rect 7198 39678 7250 39730
rect 7250 39678 7252 39730
rect 7196 39676 7252 39678
rect 6412 39340 6468 39396
rect 7644 39394 7700 39396
rect 7644 39342 7646 39394
rect 7646 39342 7698 39394
rect 7698 39342 7700 39394
rect 7644 39340 7700 39342
rect 6412 38780 6468 38836
rect 5852 36594 5908 36596
rect 5852 36542 5854 36594
rect 5854 36542 5906 36594
rect 5906 36542 5908 36594
rect 5852 36540 5908 36542
rect 5964 36482 6020 36484
rect 5964 36430 5966 36482
rect 5966 36430 6018 36482
rect 6018 36430 6020 36482
rect 5964 36428 6020 36430
rect 5964 35420 6020 35476
rect 5516 34914 5572 34916
rect 5516 34862 5518 34914
rect 5518 34862 5570 34914
rect 5570 34862 5572 34914
rect 5516 34860 5572 34862
rect 5292 33516 5348 33572
rect 5068 32956 5124 33012
rect 3724 30156 3780 30212
rect 4172 29650 4228 29652
rect 4172 29598 4174 29650
rect 4174 29598 4226 29650
rect 4226 29598 4228 29650
rect 4172 29596 4228 29598
rect 3836 29426 3892 29428
rect 3836 29374 3838 29426
rect 3838 29374 3890 29426
rect 3890 29374 3892 29426
rect 3836 29372 3892 29374
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4844 29596 4900 29652
rect 4396 29260 4452 29316
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4284 28642 4340 28644
rect 4284 28590 4286 28642
rect 4286 28590 4338 28642
rect 4338 28590 4340 28642
rect 4284 28588 4340 28590
rect 4956 28700 5012 28756
rect 5404 32956 5460 33012
rect 6300 35084 6356 35140
rect 7196 38780 7252 38836
rect 7532 37660 7588 37716
rect 6636 37548 6692 37604
rect 7532 37490 7588 37492
rect 7532 37438 7534 37490
rect 7534 37438 7586 37490
rect 7586 37438 7588 37490
rect 7532 37436 7588 37438
rect 6748 37378 6804 37380
rect 6748 37326 6750 37378
rect 6750 37326 6802 37378
rect 6802 37326 6804 37378
rect 6748 37324 6804 37326
rect 6972 37266 7028 37268
rect 6972 37214 6974 37266
rect 6974 37214 7026 37266
rect 7026 37214 7028 37266
rect 6972 37212 7028 37214
rect 7196 37212 7252 37268
rect 6636 36652 6692 36708
rect 6524 36482 6580 36484
rect 6524 36430 6526 36482
rect 6526 36430 6578 36482
rect 6578 36430 6580 36482
rect 6524 36428 6580 36430
rect 6748 36370 6804 36372
rect 6748 36318 6750 36370
rect 6750 36318 6802 36370
rect 6802 36318 6804 36370
rect 6748 36316 6804 36318
rect 7308 36876 7364 36932
rect 6860 36092 6916 36148
rect 7084 35980 7140 36036
rect 6636 35868 6692 35924
rect 7196 35868 7252 35924
rect 7756 37826 7812 37828
rect 7756 37774 7758 37826
rect 7758 37774 7810 37826
rect 7810 37774 7812 37826
rect 7756 37772 7812 37774
rect 7756 35868 7812 35924
rect 6748 35532 6804 35588
rect 7084 35474 7140 35476
rect 7084 35422 7086 35474
rect 7086 35422 7138 35474
rect 7138 35422 7140 35474
rect 7084 35420 7140 35422
rect 7644 35196 7700 35252
rect 7084 34802 7140 34804
rect 7084 34750 7086 34802
rect 7086 34750 7138 34802
rect 7138 34750 7140 34802
rect 7084 34748 7140 34750
rect 6748 34076 6804 34132
rect 6636 33964 6692 34020
rect 6748 33906 6804 33908
rect 6748 33854 6750 33906
rect 6750 33854 6802 33906
rect 6802 33854 6804 33906
rect 6748 33852 6804 33854
rect 6972 33740 7028 33796
rect 6076 33516 6132 33572
rect 7084 33068 7140 33124
rect 6188 32674 6244 32676
rect 6188 32622 6190 32674
rect 6190 32622 6242 32674
rect 6242 32622 6244 32674
rect 6188 32620 6244 32622
rect 6076 31948 6132 32004
rect 7308 33964 7364 34020
rect 5516 31388 5572 31444
rect 7308 32956 7364 33012
rect 6748 31948 6804 32004
rect 5740 30156 5796 30212
rect 5068 29372 5124 29428
rect 4284 27858 4340 27860
rect 4284 27806 4286 27858
rect 4286 27806 4338 27858
rect 4338 27806 4340 27858
rect 4284 27804 4340 27806
rect 3724 27020 3780 27076
rect 4172 27074 4228 27076
rect 4172 27022 4174 27074
rect 4174 27022 4226 27074
rect 4226 27022 4228 27074
rect 4172 27020 4228 27022
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3836 25228 3892 25284
rect 3836 24050 3892 24052
rect 3836 23998 3838 24050
rect 3838 23998 3890 24050
rect 3890 23998 3892 24050
rect 3836 23996 3892 23998
rect 3612 23042 3668 23044
rect 3612 22990 3614 23042
rect 3614 22990 3666 23042
rect 3666 22990 3668 23042
rect 3612 22988 3668 22990
rect 3500 21644 3556 21700
rect 3164 18338 3220 18340
rect 3164 18286 3166 18338
rect 3166 18286 3218 18338
rect 3218 18286 3220 18338
rect 3164 18284 3220 18286
rect 3276 17778 3332 17780
rect 3276 17726 3278 17778
rect 3278 17726 3330 17778
rect 3330 17726 3332 17778
rect 3276 17724 3332 17726
rect 2940 17052 2996 17108
rect 3948 21308 4004 21364
rect 3836 20914 3892 20916
rect 3836 20862 3838 20914
rect 3838 20862 3890 20914
rect 3890 20862 3892 20914
rect 3836 20860 3892 20862
rect 3836 19852 3892 19908
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4844 25452 4900 25508
rect 4284 25340 4340 25396
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 6748 29708 6804 29764
rect 6076 29260 6132 29316
rect 6636 29148 6692 29204
rect 5852 26460 5908 26516
rect 5852 25618 5908 25620
rect 5852 25566 5854 25618
rect 5854 25566 5906 25618
rect 5906 25566 5908 25618
rect 5852 25564 5908 25566
rect 5740 25394 5796 25396
rect 5740 25342 5742 25394
rect 5742 25342 5794 25394
rect 5794 25342 5796 25394
rect 5740 25340 5796 25342
rect 5068 24444 5124 24500
rect 5740 24556 5796 24612
rect 4284 23772 4340 23828
rect 4172 22988 4228 23044
rect 5628 23826 5684 23828
rect 5628 23774 5630 23826
rect 5630 23774 5682 23826
rect 5682 23774 5684 23826
rect 5628 23772 5684 23774
rect 5740 23660 5796 23716
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4284 20748 4340 20804
rect 5180 21474 5236 21476
rect 5180 21422 5182 21474
rect 5182 21422 5234 21474
rect 5234 21422 5236 21474
rect 5180 21420 5236 21422
rect 5068 20748 5124 20804
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 3500 17836 3556 17892
rect 3836 18284 3892 18340
rect 3276 16940 3332 16996
rect 2604 16156 2660 16212
rect 2604 14924 2660 14980
rect 2268 14700 2324 14756
rect 1820 13692 1876 13748
rect 1596 11564 1652 11620
rect 1708 11676 1764 11732
rect 1708 11004 1764 11060
rect 1708 9714 1764 9716
rect 1708 9662 1710 9714
rect 1710 9662 1762 9714
rect 1762 9662 1764 9714
rect 1708 9660 1764 9662
rect 2156 14252 2212 14308
rect 3052 16098 3108 16100
rect 3052 16046 3054 16098
rect 3054 16046 3106 16098
rect 3106 16046 3108 16098
rect 3052 16044 3108 16046
rect 2940 15986 2996 15988
rect 2940 15934 2942 15986
rect 2942 15934 2994 15986
rect 2994 15934 2996 15986
rect 2940 15932 2996 15934
rect 3276 16098 3332 16100
rect 3276 16046 3278 16098
rect 3278 16046 3330 16098
rect 3330 16046 3332 16098
rect 3276 16044 3332 16046
rect 3388 15820 3444 15876
rect 3052 15090 3108 15092
rect 3052 15038 3054 15090
rect 3054 15038 3106 15090
rect 3106 15038 3108 15090
rect 3052 15036 3108 15038
rect 2492 14140 2548 14196
rect 2716 13970 2772 13972
rect 2716 13918 2718 13970
rect 2718 13918 2770 13970
rect 2770 13918 2772 13970
rect 2716 13916 2772 13918
rect 3164 13804 3220 13860
rect 2268 12178 2324 12180
rect 2268 12126 2270 12178
rect 2270 12126 2322 12178
rect 2322 12126 2324 12178
rect 2268 12124 2324 12126
rect 2268 10610 2324 10612
rect 2268 10558 2270 10610
rect 2270 10558 2322 10610
rect 2322 10558 2324 10610
rect 2268 10556 2324 10558
rect 2268 9938 2324 9940
rect 2268 9886 2270 9938
rect 2270 9886 2322 9938
rect 2322 9886 2324 9938
rect 2268 9884 2324 9886
rect 2044 9324 2100 9380
rect 1708 8316 1764 8372
rect 1708 6972 1764 7028
rect 2604 12796 2660 12852
rect 2492 8316 2548 8372
rect 2492 6972 2548 7028
rect 1708 5628 1764 5684
rect 1708 4844 1764 4900
rect 1708 4284 1764 4340
rect 2156 6076 2212 6132
rect 2492 5628 2548 5684
rect 3500 15260 3556 15316
rect 3836 16882 3892 16884
rect 3836 16830 3838 16882
rect 3838 16830 3890 16882
rect 3890 16830 3892 16882
rect 3836 16828 3892 16830
rect 3948 17836 4004 17892
rect 4732 18396 4788 18452
rect 4508 18284 4564 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 6076 22428 6132 22484
rect 6076 21308 6132 21364
rect 6300 28588 6356 28644
rect 6636 28700 6692 28756
rect 7084 31890 7140 31892
rect 7084 31838 7086 31890
rect 7086 31838 7138 31890
rect 7138 31838 7140 31890
rect 7084 31836 7140 31838
rect 7420 32732 7476 32788
rect 7532 33852 7588 33908
rect 6972 29596 7028 29652
rect 7420 30940 7476 30996
rect 6860 27468 6916 27524
rect 7084 27132 7140 27188
rect 6748 27074 6804 27076
rect 6748 27022 6750 27074
rect 6750 27022 6802 27074
rect 6802 27022 6804 27074
rect 6748 27020 6804 27022
rect 6860 26850 6916 26852
rect 6860 26798 6862 26850
rect 6862 26798 6914 26850
rect 6914 26798 6916 26850
rect 6860 26796 6916 26798
rect 6972 26514 7028 26516
rect 6972 26462 6974 26514
rect 6974 26462 7026 26514
rect 7026 26462 7028 26514
rect 6972 26460 7028 26462
rect 7084 26402 7140 26404
rect 7084 26350 7086 26402
rect 7086 26350 7138 26402
rect 7138 26350 7140 26402
rect 7084 26348 7140 26350
rect 7308 26796 7364 26852
rect 7084 25900 7140 25956
rect 7308 25618 7364 25620
rect 7308 25566 7310 25618
rect 7310 25566 7362 25618
rect 7362 25566 7364 25618
rect 7308 25564 7364 25566
rect 6524 25452 6580 25508
rect 6972 25282 7028 25284
rect 6972 25230 6974 25282
rect 6974 25230 7026 25282
rect 7026 25230 7028 25282
rect 6972 25228 7028 25230
rect 7644 33628 7700 33684
rect 7756 33852 7812 33908
rect 7980 38892 8036 38948
rect 8316 40572 8372 40628
rect 8204 39676 8260 39732
rect 7980 37884 8036 37940
rect 8092 38444 8148 38500
rect 7980 37660 8036 37716
rect 7980 36764 8036 36820
rect 8428 36988 8484 37044
rect 8316 36876 8372 36932
rect 8652 39340 8708 39396
rect 8764 38722 8820 38724
rect 8764 38670 8766 38722
rect 8766 38670 8818 38722
rect 8818 38670 8820 38722
rect 8764 38668 8820 38670
rect 9660 40626 9716 40628
rect 9660 40574 9662 40626
rect 9662 40574 9714 40626
rect 9714 40574 9716 40626
rect 9660 40572 9716 40574
rect 11228 41298 11284 41300
rect 11228 41246 11230 41298
rect 11230 41246 11282 41298
rect 11282 41246 11284 41298
rect 11228 41244 11284 41246
rect 12124 41244 12180 41300
rect 11452 41074 11508 41076
rect 11452 41022 11454 41074
rect 11454 41022 11506 41074
rect 11506 41022 11508 41074
rect 11452 41020 11508 41022
rect 10556 40348 10612 40404
rect 11452 40402 11508 40404
rect 11452 40350 11454 40402
rect 11454 40350 11506 40402
rect 11506 40350 11508 40402
rect 11452 40348 11508 40350
rect 11900 40684 11956 40740
rect 11676 40514 11732 40516
rect 11676 40462 11678 40514
rect 11678 40462 11730 40514
rect 11730 40462 11732 40514
rect 11676 40460 11732 40462
rect 12348 40402 12404 40404
rect 12348 40350 12350 40402
rect 12350 40350 12402 40402
rect 12402 40350 12404 40402
rect 12348 40348 12404 40350
rect 9436 38834 9492 38836
rect 9436 38782 9438 38834
rect 9438 38782 9490 38834
rect 9490 38782 9492 38834
rect 9436 38780 9492 38782
rect 8540 36876 8596 36932
rect 8092 36652 8148 36708
rect 8428 36764 8484 36820
rect 8092 36482 8148 36484
rect 8092 36430 8094 36482
rect 8094 36430 8146 36482
rect 8146 36430 8148 36482
rect 8092 36428 8148 36430
rect 8988 36764 9044 36820
rect 8428 36482 8484 36484
rect 8428 36430 8430 36482
rect 8430 36430 8482 36482
rect 8482 36430 8484 36482
rect 8428 36428 8484 36430
rect 8764 36428 8820 36484
rect 8204 36316 8260 36372
rect 7980 35532 8036 35588
rect 8764 36092 8820 36148
rect 8204 35196 8260 35252
rect 8540 35586 8596 35588
rect 8540 35534 8542 35586
rect 8542 35534 8594 35586
rect 8594 35534 8596 35586
rect 8540 35532 8596 35534
rect 8092 33852 8148 33908
rect 7756 33234 7812 33236
rect 7756 33182 7758 33234
rect 7758 33182 7810 33234
rect 7810 33182 7812 33234
rect 7756 33180 7812 33182
rect 7644 32562 7700 32564
rect 7644 32510 7646 32562
rect 7646 32510 7698 32562
rect 7698 32510 7700 32562
rect 7644 32508 7700 32510
rect 7756 32396 7812 32452
rect 8092 32956 8148 33012
rect 7644 31500 7700 31556
rect 7532 27132 7588 27188
rect 6972 24610 7028 24612
rect 6972 24558 6974 24610
rect 6974 24558 7026 24610
rect 7026 24558 7028 24610
rect 6972 24556 7028 24558
rect 6860 23996 6916 24052
rect 6524 21532 6580 21588
rect 5740 19068 5796 19124
rect 5516 18450 5572 18452
rect 5516 18398 5518 18450
rect 5518 18398 5570 18450
rect 5570 18398 5572 18450
rect 5516 18396 5572 18398
rect 5404 18060 5460 18116
rect 4172 17836 4228 17892
rect 4284 17612 4340 17668
rect 4172 17500 4228 17556
rect 4508 17164 4564 17220
rect 4396 16940 4452 16996
rect 4284 16828 4340 16884
rect 4620 16770 4676 16772
rect 4620 16718 4622 16770
rect 4622 16718 4674 16770
rect 4674 16718 4676 16770
rect 4620 16716 4676 16718
rect 3948 16268 4004 16324
rect 3948 16044 4004 16100
rect 3388 14140 3444 14196
rect 3276 13580 3332 13636
rect 3052 12796 3108 12852
rect 2716 12402 2772 12404
rect 2716 12350 2718 12402
rect 2718 12350 2770 12402
rect 2770 12350 2772 12402
rect 2716 12348 2772 12350
rect 3164 11676 3220 11732
rect 2940 11282 2996 11284
rect 2940 11230 2942 11282
rect 2942 11230 2994 11282
rect 2994 11230 2996 11282
rect 2940 11228 2996 11230
rect 3052 11116 3108 11172
rect 4172 16156 4228 16212
rect 4172 15260 4228 15316
rect 3836 15036 3892 15092
rect 3500 13132 3556 13188
rect 3948 13634 4004 13636
rect 3948 13582 3950 13634
rect 3950 13582 4002 13634
rect 4002 13582 4004 13634
rect 3948 13580 4004 13582
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4844 16268 4900 16324
rect 4508 16210 4564 16212
rect 4508 16158 4510 16210
rect 4510 16158 4562 16210
rect 4562 16158 4564 16210
rect 4508 16156 4564 16158
rect 4732 16098 4788 16100
rect 4732 16046 4734 16098
rect 4734 16046 4786 16098
rect 4786 16046 4788 16098
rect 4732 16044 4788 16046
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4284 14588 4340 14644
rect 4508 14140 4564 14196
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4284 13132 4340 13188
rect 3500 12850 3556 12852
rect 3500 12798 3502 12850
rect 3502 12798 3554 12850
rect 3554 12798 3556 12850
rect 3500 12796 3556 12798
rect 4172 11900 4228 11956
rect 5068 17948 5124 18004
rect 5516 17836 5572 17892
rect 5068 17666 5124 17668
rect 5068 17614 5070 17666
rect 5070 17614 5122 17666
rect 5122 17614 5124 17666
rect 5068 17612 5124 17614
rect 5292 17612 5348 17668
rect 5292 17052 5348 17108
rect 5852 17666 5908 17668
rect 5852 17614 5854 17666
rect 5854 17614 5906 17666
rect 5906 17614 5908 17666
rect 5852 17612 5908 17614
rect 5740 16828 5796 16884
rect 5068 15986 5124 15988
rect 5068 15934 5070 15986
rect 5070 15934 5122 15986
rect 5122 15934 5124 15986
rect 5068 15932 5124 15934
rect 5852 16940 5908 16996
rect 5852 16156 5908 16212
rect 5740 15820 5796 15876
rect 5740 15260 5796 15316
rect 5628 15036 5684 15092
rect 5068 14642 5124 14644
rect 5068 14590 5070 14642
rect 5070 14590 5122 14642
rect 5122 14590 5124 14642
rect 5068 14588 5124 14590
rect 6412 19068 6468 19124
rect 6636 18396 6692 18452
rect 6300 18284 6356 18340
rect 6076 17724 6132 17780
rect 6636 17612 6692 17668
rect 6524 17052 6580 17108
rect 6300 16380 6356 16436
rect 6076 15314 6132 15316
rect 6076 15262 6078 15314
rect 6078 15262 6130 15314
rect 6130 15262 6132 15314
rect 6076 15260 6132 15262
rect 6860 17612 6916 17668
rect 6860 16940 6916 16996
rect 6972 16882 7028 16884
rect 6972 16830 6974 16882
rect 6974 16830 7026 16882
rect 7026 16830 7028 16882
rect 6972 16828 7028 16830
rect 5964 14700 6020 14756
rect 6412 14588 6468 14644
rect 7196 24668 7252 24724
rect 7196 23772 7252 23828
rect 7868 30380 7924 30436
rect 8092 31890 8148 31892
rect 8092 31838 8094 31890
rect 8094 31838 8146 31890
rect 8146 31838 8148 31890
rect 8092 31836 8148 31838
rect 8092 31612 8148 31668
rect 8316 31388 8372 31444
rect 8652 32786 8708 32788
rect 8652 32734 8654 32786
rect 8654 32734 8706 32786
rect 8706 32734 8708 32786
rect 8652 32732 8708 32734
rect 8764 32172 8820 32228
rect 8876 31948 8932 32004
rect 8540 31500 8596 31556
rect 8204 31052 8260 31108
rect 8316 31164 8372 31220
rect 8092 30268 8148 30324
rect 7868 29596 7924 29652
rect 7868 27468 7924 27524
rect 7756 25564 7812 25620
rect 7756 24892 7812 24948
rect 7532 24668 7588 24724
rect 7420 20972 7476 21028
rect 7532 20636 7588 20692
rect 7308 19234 7364 19236
rect 7308 19182 7310 19234
rect 7310 19182 7362 19234
rect 7362 19182 7364 19234
rect 7308 19180 7364 19182
rect 7196 18450 7252 18452
rect 7196 18398 7198 18450
rect 7198 18398 7250 18450
rect 7250 18398 7252 18450
rect 7196 18396 7252 18398
rect 7756 23436 7812 23492
rect 7868 19068 7924 19124
rect 7644 18674 7700 18676
rect 7644 18622 7646 18674
rect 7646 18622 7698 18674
rect 7698 18622 7700 18674
rect 7644 18620 7700 18622
rect 7868 18562 7924 18564
rect 7868 18510 7870 18562
rect 7870 18510 7922 18562
rect 7922 18510 7924 18562
rect 7868 18508 7924 18510
rect 7532 18060 7588 18116
rect 7196 16828 7252 16884
rect 7308 17948 7364 18004
rect 7420 17612 7476 17668
rect 7868 17666 7924 17668
rect 7868 17614 7870 17666
rect 7870 17614 7922 17666
rect 7922 17614 7924 17666
rect 7868 17612 7924 17614
rect 7532 16994 7588 16996
rect 7532 16942 7534 16994
rect 7534 16942 7586 16994
rect 7586 16942 7588 16994
rect 7532 16940 7588 16942
rect 7420 14642 7476 14644
rect 7420 14590 7422 14642
rect 7422 14590 7474 14642
rect 7474 14590 7476 14642
rect 7420 14588 7476 14590
rect 7644 15036 7700 15092
rect 7756 15260 7812 15316
rect 8428 28364 8484 28420
rect 8428 23884 8484 23940
rect 8316 23042 8372 23044
rect 8316 22990 8318 23042
rect 8318 22990 8370 23042
rect 8370 22990 8372 23042
rect 8316 22988 8372 22990
rect 8316 22092 8372 22148
rect 9324 36876 9380 36932
rect 9212 31276 9268 31332
rect 9100 28700 9156 28756
rect 8092 19964 8148 20020
rect 8092 18620 8148 18676
rect 8540 21196 8596 21252
rect 9436 36482 9492 36484
rect 9436 36430 9438 36482
rect 9438 36430 9490 36482
rect 9490 36430 9492 36482
rect 9436 36428 9492 36430
rect 9772 37884 9828 37940
rect 9548 36258 9604 36260
rect 9548 36206 9550 36258
rect 9550 36206 9602 36258
rect 9602 36206 9604 36258
rect 9548 36204 9604 36206
rect 9548 35532 9604 35588
rect 9884 37100 9940 37156
rect 11340 38108 11396 38164
rect 10556 37938 10612 37940
rect 10556 37886 10558 37938
rect 10558 37886 10610 37938
rect 10610 37886 10612 37938
rect 10556 37884 10612 37886
rect 9772 35196 9828 35252
rect 10556 37100 10612 37156
rect 12236 39676 12292 39732
rect 12012 39394 12068 39396
rect 12012 39342 12014 39394
rect 12014 39342 12066 39394
rect 12066 39342 12068 39394
rect 12012 39340 12068 39342
rect 11788 38162 11844 38164
rect 11788 38110 11790 38162
rect 11790 38110 11842 38162
rect 11842 38110 11844 38162
rect 11788 38108 11844 38110
rect 11564 37212 11620 37268
rect 12124 37772 12180 37828
rect 11116 37154 11172 37156
rect 11116 37102 11118 37154
rect 11118 37102 11170 37154
rect 11170 37102 11172 37154
rect 11116 37100 11172 37102
rect 10444 36428 10500 36484
rect 11004 36876 11060 36932
rect 10220 36258 10276 36260
rect 10220 36206 10222 36258
rect 10222 36206 10274 36258
rect 10274 36206 10276 36258
rect 10220 36204 10276 36206
rect 10108 35084 10164 35140
rect 10332 35196 10388 35252
rect 10444 34860 10500 34916
rect 9660 33122 9716 33124
rect 9660 33070 9662 33122
rect 9662 33070 9714 33122
rect 9714 33070 9716 33122
rect 9660 33068 9716 33070
rect 9996 33122 10052 33124
rect 9996 33070 9998 33122
rect 9998 33070 10050 33122
rect 10050 33070 10052 33122
rect 9996 33068 10052 33070
rect 9884 32508 9940 32564
rect 9772 31724 9828 31780
rect 9996 31666 10052 31668
rect 9996 31614 9998 31666
rect 9998 31614 10050 31666
rect 10050 31614 10052 31666
rect 9996 31612 10052 31614
rect 9660 31500 9716 31556
rect 8988 21586 9044 21588
rect 8988 21534 8990 21586
rect 8990 21534 9042 21586
rect 9042 21534 9044 21586
rect 8988 21532 9044 21534
rect 8316 17948 8372 18004
rect 8540 16716 8596 16772
rect 10220 32844 10276 32900
rect 10332 32956 10388 33012
rect 11228 36652 11284 36708
rect 10892 33740 10948 33796
rect 10892 33346 10948 33348
rect 10892 33294 10894 33346
rect 10894 33294 10946 33346
rect 10946 33294 10948 33346
rect 10892 33292 10948 33294
rect 11340 35308 11396 35364
rect 11340 34860 11396 34916
rect 11564 35084 11620 35140
rect 10780 33234 10836 33236
rect 10780 33182 10782 33234
rect 10782 33182 10834 33234
rect 10834 33182 10836 33234
rect 10780 33180 10836 33182
rect 10556 32844 10612 32900
rect 10668 33122 10724 33124
rect 10668 33070 10670 33122
rect 10670 33070 10722 33122
rect 10722 33070 10724 33122
rect 10668 33068 10724 33070
rect 10220 31948 10276 32004
rect 10556 31836 10612 31892
rect 10220 31500 10276 31556
rect 10892 31276 10948 31332
rect 10108 31106 10164 31108
rect 10108 31054 10110 31106
rect 10110 31054 10162 31106
rect 10162 31054 10164 31106
rect 10108 31052 10164 31054
rect 10108 30156 10164 30212
rect 10108 29932 10164 29988
rect 9996 27804 10052 27860
rect 10108 27692 10164 27748
rect 9772 25676 9828 25732
rect 9660 25116 9716 25172
rect 9996 24834 10052 24836
rect 9996 24782 9998 24834
rect 9998 24782 10050 24834
rect 10050 24782 10052 24834
rect 9996 24780 10052 24782
rect 9884 24610 9940 24612
rect 9884 24558 9886 24610
rect 9886 24558 9938 24610
rect 9938 24558 9940 24610
rect 9884 24556 9940 24558
rect 10108 24332 10164 24388
rect 9772 23714 9828 23716
rect 9772 23662 9774 23714
rect 9774 23662 9826 23714
rect 9826 23662 9828 23714
rect 9772 23660 9828 23662
rect 10108 23938 10164 23940
rect 10108 23886 10110 23938
rect 10110 23886 10162 23938
rect 10162 23886 10164 23938
rect 10108 23884 10164 23886
rect 11228 32284 11284 32340
rect 11452 32060 11508 32116
rect 11004 30604 11060 30660
rect 10332 30492 10388 30548
rect 11340 31666 11396 31668
rect 11340 31614 11342 31666
rect 11342 31614 11394 31666
rect 11394 31614 11396 31666
rect 11340 31612 11396 31614
rect 12124 35644 12180 35700
rect 12012 34690 12068 34692
rect 12012 34638 12014 34690
rect 12014 34638 12066 34690
rect 12066 34638 12068 34690
rect 12012 34636 12068 34638
rect 11900 33516 11956 33572
rect 12124 33068 12180 33124
rect 12572 38444 12628 38500
rect 12348 37266 12404 37268
rect 12348 37214 12350 37266
rect 12350 37214 12402 37266
rect 12402 37214 12404 37266
rect 12348 37212 12404 37214
rect 12572 35308 12628 35364
rect 12348 33516 12404 33572
rect 12572 33068 12628 33124
rect 11900 32284 11956 32340
rect 11564 31388 11620 31444
rect 11676 31948 11732 32004
rect 11676 31276 11732 31332
rect 11228 30492 11284 30548
rect 12012 30770 12068 30772
rect 12012 30718 12014 30770
rect 12014 30718 12066 30770
rect 12066 30718 12068 30770
rect 12012 30716 12068 30718
rect 11788 30434 11844 30436
rect 11788 30382 11790 30434
rect 11790 30382 11842 30434
rect 11842 30382 11844 30434
rect 11788 30380 11844 30382
rect 11676 30268 11732 30324
rect 11452 30156 11508 30212
rect 11116 30098 11172 30100
rect 11116 30046 11118 30098
rect 11118 30046 11170 30098
rect 11170 30046 11172 30098
rect 11116 30044 11172 30046
rect 12012 30210 12068 30212
rect 12012 30158 12014 30210
rect 12014 30158 12066 30210
rect 12066 30158 12068 30210
rect 12012 30156 12068 30158
rect 12236 32060 12292 32116
rect 12572 32284 12628 32340
rect 12348 30940 12404 30996
rect 12460 31388 12516 31444
rect 11452 29820 11508 29876
rect 11676 29986 11732 29988
rect 11676 29934 11678 29986
rect 11678 29934 11730 29986
rect 11730 29934 11732 29986
rect 11676 29932 11732 29934
rect 10332 28642 10388 28644
rect 10332 28590 10334 28642
rect 10334 28590 10386 28642
rect 10386 28590 10388 28642
rect 10332 28588 10388 28590
rect 10780 28418 10836 28420
rect 10780 28366 10782 28418
rect 10782 28366 10834 28418
rect 10834 28366 10836 28418
rect 10780 28364 10836 28366
rect 10556 27468 10612 27524
rect 10332 25676 10388 25732
rect 10332 23772 10388 23828
rect 11004 27692 11060 27748
rect 11116 27132 11172 27188
rect 11340 28866 11396 28868
rect 11340 28814 11342 28866
rect 11342 28814 11394 28866
rect 11394 28814 11396 28866
rect 11340 28812 11396 28814
rect 11788 28700 11844 28756
rect 11340 28476 11396 28532
rect 11340 27746 11396 27748
rect 11340 27694 11342 27746
rect 11342 27694 11394 27746
rect 11394 27694 11396 27746
rect 11340 27692 11396 27694
rect 11900 28642 11956 28644
rect 11900 28590 11902 28642
rect 11902 28590 11954 28642
rect 11954 28590 11956 28642
rect 11900 28588 11956 28590
rect 12236 28530 12292 28532
rect 12236 28478 12238 28530
rect 12238 28478 12290 28530
rect 12290 28478 12292 28530
rect 12236 28476 12292 28478
rect 11564 27634 11620 27636
rect 11564 27582 11566 27634
rect 11566 27582 11618 27634
rect 11618 27582 11620 27634
rect 11564 27580 11620 27582
rect 11788 27356 11844 27412
rect 12124 27858 12180 27860
rect 12124 27806 12126 27858
rect 12126 27806 12178 27858
rect 12178 27806 12180 27858
rect 12124 27804 12180 27806
rect 12908 39394 12964 39396
rect 12908 39342 12910 39394
rect 12910 39342 12962 39394
rect 12962 39342 12964 39394
rect 12908 39340 12964 39342
rect 13468 39730 13524 39732
rect 13468 39678 13470 39730
rect 13470 39678 13522 39730
rect 13522 39678 13524 39730
rect 13468 39676 13524 39678
rect 12908 37660 12964 37716
rect 13020 35756 13076 35812
rect 12796 35644 12852 35700
rect 13020 35586 13076 35588
rect 13020 35534 13022 35586
rect 13022 35534 13074 35586
rect 13074 35534 13076 35586
rect 13020 35532 13076 35534
rect 12796 34690 12852 34692
rect 12796 34638 12798 34690
rect 12798 34638 12850 34690
rect 12850 34638 12852 34690
rect 12796 34636 12852 34638
rect 12796 34130 12852 34132
rect 12796 34078 12798 34130
rect 12798 34078 12850 34130
rect 12850 34078 12852 34130
rect 12796 34076 12852 34078
rect 12908 33740 12964 33796
rect 13356 34636 13412 34692
rect 13468 35756 13524 35812
rect 13356 34018 13412 34020
rect 13356 33966 13358 34018
rect 13358 33966 13410 34018
rect 13410 33966 13412 34018
rect 13356 33964 13412 33966
rect 13132 31948 13188 32004
rect 12908 31164 12964 31220
rect 12572 30156 12628 30212
rect 12796 28700 12852 28756
rect 12460 27970 12516 27972
rect 12460 27918 12462 27970
rect 12462 27918 12514 27970
rect 12514 27918 12516 27970
rect 12460 27916 12516 27918
rect 12348 27746 12404 27748
rect 12348 27694 12350 27746
rect 12350 27694 12402 27746
rect 12402 27694 12404 27746
rect 12348 27692 12404 27694
rect 12236 27580 12292 27636
rect 11452 27132 11508 27188
rect 11564 27020 11620 27076
rect 12908 28476 12964 28532
rect 12908 27692 12964 27748
rect 12908 27356 12964 27412
rect 10556 24946 10612 24948
rect 10556 24894 10558 24946
rect 10558 24894 10610 24946
rect 10610 24894 10612 24946
rect 10556 24892 10612 24894
rect 10780 25228 10836 25284
rect 10780 24780 10836 24836
rect 10892 24722 10948 24724
rect 10892 24670 10894 24722
rect 10894 24670 10946 24722
rect 10946 24670 10948 24722
rect 10892 24668 10948 24670
rect 11116 24610 11172 24612
rect 11116 24558 11118 24610
rect 11118 24558 11170 24610
rect 11170 24558 11172 24610
rect 11116 24556 11172 24558
rect 9996 23436 10052 23492
rect 10444 23324 10500 23380
rect 10108 22652 10164 22708
rect 9324 22482 9380 22484
rect 9324 22430 9326 22482
rect 9326 22430 9378 22482
rect 9378 22430 9380 22482
rect 9324 22428 9380 22430
rect 9884 22428 9940 22484
rect 9548 20018 9604 20020
rect 9548 19966 9550 20018
rect 9550 19966 9602 20018
rect 9602 19966 9604 20018
rect 9548 19964 9604 19966
rect 10668 22652 10724 22708
rect 10668 22428 10724 22484
rect 10332 22370 10388 22372
rect 10332 22318 10334 22370
rect 10334 22318 10386 22370
rect 10386 22318 10388 22370
rect 10332 22316 10388 22318
rect 10556 22146 10612 22148
rect 10556 22094 10558 22146
rect 10558 22094 10610 22146
rect 10610 22094 10612 22146
rect 10556 22092 10612 22094
rect 10220 21474 10276 21476
rect 10220 21422 10222 21474
rect 10222 21422 10274 21474
rect 10274 21422 10276 21474
rect 10220 21420 10276 21422
rect 9884 19964 9940 20020
rect 9996 21196 10052 21252
rect 11116 22482 11172 22484
rect 11116 22430 11118 22482
rect 11118 22430 11170 22482
rect 11170 22430 11172 22482
rect 11116 22428 11172 22430
rect 11564 25900 11620 25956
rect 11452 23324 11508 23380
rect 11340 22540 11396 22596
rect 11228 22092 11284 22148
rect 10892 21980 10948 22036
rect 11340 21980 11396 22036
rect 10556 21196 10612 21252
rect 10332 20860 10388 20916
rect 10108 20690 10164 20692
rect 10108 20638 10110 20690
rect 10110 20638 10162 20690
rect 10162 20638 10164 20690
rect 10108 20636 10164 20638
rect 11228 21308 11284 21364
rect 10780 20636 10836 20692
rect 10108 20018 10164 20020
rect 10108 19966 10110 20018
rect 10110 19966 10162 20018
rect 10162 19966 10164 20018
rect 10108 19964 10164 19966
rect 11452 20524 11508 20580
rect 12124 26348 12180 26404
rect 12012 25900 12068 25956
rect 12572 26124 12628 26180
rect 12572 25900 12628 25956
rect 11676 24556 11732 24612
rect 12572 25004 12628 25060
rect 12796 25116 12852 25172
rect 12684 24946 12740 24948
rect 12684 24894 12686 24946
rect 12686 24894 12738 24946
rect 12738 24894 12740 24946
rect 12684 24892 12740 24894
rect 12236 23100 12292 23156
rect 12012 22988 12068 23044
rect 12012 22482 12068 22484
rect 12012 22430 12014 22482
rect 12014 22430 12066 22482
rect 12066 22430 12068 22482
rect 12012 22428 12068 22430
rect 11788 21196 11844 21252
rect 11564 20188 11620 20244
rect 11788 20972 11844 21028
rect 9660 18620 9716 18676
rect 9548 18172 9604 18228
rect 9100 16380 9156 16436
rect 9548 17948 9604 18004
rect 5740 13356 5796 13412
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 5852 13074 5908 13076
rect 5852 13022 5854 13074
rect 5854 13022 5906 13074
rect 5906 13022 5908 13074
rect 5852 13020 5908 13022
rect 5852 12796 5908 12852
rect 5516 11900 5572 11956
rect 5740 12012 5796 12068
rect 4956 11788 5012 11844
rect 4844 11340 4900 11396
rect 6636 13074 6692 13076
rect 6636 13022 6638 13074
rect 6638 13022 6690 13074
rect 6690 13022 6692 13074
rect 6636 13020 6692 13022
rect 6300 12402 6356 12404
rect 6300 12350 6302 12402
rect 6302 12350 6354 12402
rect 6354 12350 6356 12402
rect 6300 12348 6356 12350
rect 6188 12012 6244 12068
rect 5852 11788 5908 11844
rect 6076 11900 6132 11956
rect 5852 11170 5908 11172
rect 5852 11118 5854 11170
rect 5854 11118 5906 11170
rect 5906 11118 5908 11170
rect 5852 11116 5908 11118
rect 4844 10556 4900 10612
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4284 9884 4340 9940
rect 5852 10722 5908 10724
rect 5852 10670 5854 10722
rect 5854 10670 5906 10722
rect 5906 10670 5908 10722
rect 5852 10668 5908 10670
rect 6188 11228 6244 11284
rect 6300 11116 6356 11172
rect 7084 13020 7140 13076
rect 6636 11340 6692 11396
rect 6524 10610 6580 10612
rect 6524 10558 6526 10610
rect 6526 10558 6578 10610
rect 6578 10558 6580 10610
rect 6524 10556 6580 10558
rect 6524 10332 6580 10388
rect 5964 9548 6020 9604
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 6412 9602 6468 9604
rect 6412 9550 6414 9602
rect 6414 9550 6466 9602
rect 6466 9550 6468 9602
rect 6412 9548 6468 9550
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 3276 6076 3332 6132
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 2492 4844 2548 4900
rect 1820 2940 1876 2996
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 6076 4338 6132 4340
rect 6076 4286 6078 4338
rect 6078 4286 6130 4338
rect 6130 4286 6132 4338
rect 6076 4284 6132 4286
rect 7084 12738 7140 12740
rect 7084 12686 7086 12738
rect 7086 12686 7138 12738
rect 7138 12686 7140 12738
rect 7084 12684 7140 12686
rect 7756 12402 7812 12404
rect 7756 12350 7758 12402
rect 7758 12350 7810 12402
rect 7810 12350 7812 12402
rect 7756 12348 7812 12350
rect 6972 12124 7028 12180
rect 7084 11954 7140 11956
rect 7084 11902 7086 11954
rect 7086 11902 7138 11954
rect 7138 11902 7140 11954
rect 7084 11900 7140 11902
rect 7420 11900 7476 11956
rect 7196 11564 7252 11620
rect 6748 10780 6804 10836
rect 6860 11116 6916 11172
rect 7196 10892 7252 10948
rect 8764 14700 8820 14756
rect 8652 14588 8708 14644
rect 9660 17052 9716 17108
rect 9996 18508 10052 18564
rect 10556 18956 10612 19012
rect 10220 18172 10276 18228
rect 9884 16882 9940 16884
rect 9884 16830 9886 16882
rect 9886 16830 9938 16882
rect 9938 16830 9940 16882
rect 9884 16828 9940 16830
rect 9772 15314 9828 15316
rect 9772 15262 9774 15314
rect 9774 15262 9826 15314
rect 9826 15262 9828 15314
rect 9772 15260 9828 15262
rect 10556 16658 10612 16660
rect 10556 16606 10558 16658
rect 10558 16606 10610 16658
rect 10610 16606 10612 16658
rect 10556 16604 10612 16606
rect 11676 19964 11732 20020
rect 11564 19068 11620 19124
rect 11564 18844 11620 18900
rect 11452 18562 11508 18564
rect 11452 18510 11454 18562
rect 11454 18510 11506 18562
rect 11506 18510 11508 18562
rect 11452 18508 11508 18510
rect 10780 16156 10836 16212
rect 10892 16492 10948 16548
rect 11116 16268 11172 16324
rect 11116 15484 11172 15540
rect 11228 16156 11284 16212
rect 12012 20242 12068 20244
rect 12012 20190 12014 20242
rect 12014 20190 12066 20242
rect 12066 20190 12068 20242
rect 12012 20188 12068 20190
rect 12348 19740 12404 19796
rect 12236 19180 12292 19236
rect 12572 24722 12628 24724
rect 12572 24670 12574 24722
rect 12574 24670 12626 24722
rect 12626 24670 12628 24722
rect 12572 24668 12628 24670
rect 13020 26178 13076 26180
rect 13020 26126 13022 26178
rect 13022 26126 13074 26178
rect 13074 26126 13076 26178
rect 13020 26124 13076 26126
rect 12796 21586 12852 21588
rect 12796 21534 12798 21586
rect 12798 21534 12850 21586
rect 12850 21534 12852 21586
rect 12796 21532 12852 21534
rect 12908 21084 12964 21140
rect 12572 20802 12628 20804
rect 12572 20750 12574 20802
rect 12574 20750 12626 20802
rect 12626 20750 12628 20802
rect 12572 20748 12628 20750
rect 12684 19404 12740 19460
rect 12460 18844 12516 18900
rect 13580 35084 13636 35140
rect 13580 32620 13636 32676
rect 13468 28642 13524 28644
rect 13468 28590 13470 28642
rect 13470 28590 13522 28642
rect 13522 28590 13524 28642
rect 13468 28588 13524 28590
rect 13468 27356 13524 27412
rect 13580 27020 13636 27076
rect 14924 39340 14980 39396
rect 14812 38780 14868 38836
rect 14140 38444 14196 38500
rect 14028 38050 14084 38052
rect 14028 37998 14030 38050
rect 14030 37998 14082 38050
rect 14082 37998 14084 38050
rect 14028 37996 14084 37998
rect 15596 39788 15652 39844
rect 15372 39340 15428 39396
rect 15484 38834 15540 38836
rect 15484 38782 15486 38834
rect 15486 38782 15538 38834
rect 15538 38782 15540 38834
rect 15484 38780 15540 38782
rect 13916 37826 13972 37828
rect 13916 37774 13918 37826
rect 13918 37774 13970 37826
rect 13970 37774 13972 37826
rect 13916 37772 13972 37774
rect 14140 37660 14196 37716
rect 13916 36540 13972 36596
rect 13916 36316 13972 36372
rect 14028 32396 14084 32452
rect 13916 31948 13972 32004
rect 14364 37436 14420 37492
rect 15484 38050 15540 38052
rect 15484 37998 15486 38050
rect 15486 37998 15538 38050
rect 15538 37998 15540 38050
rect 15484 37996 15540 37998
rect 15260 37660 15316 37716
rect 15148 37548 15204 37604
rect 16156 39676 16212 39732
rect 16268 39340 16324 39396
rect 16156 38892 16212 38948
rect 14700 36652 14756 36708
rect 15372 36988 15428 37044
rect 14924 36594 14980 36596
rect 14924 36542 14926 36594
rect 14926 36542 14978 36594
rect 14978 36542 14980 36594
rect 14924 36540 14980 36542
rect 14364 35698 14420 35700
rect 14364 35646 14366 35698
rect 14366 35646 14418 35698
rect 14418 35646 14420 35698
rect 14364 35644 14420 35646
rect 15036 34412 15092 34468
rect 14588 33628 14644 33684
rect 14700 33404 14756 33460
rect 14364 32674 14420 32676
rect 14364 32622 14366 32674
rect 14366 32622 14418 32674
rect 14418 32622 14420 32674
rect 14364 32620 14420 32622
rect 14924 32562 14980 32564
rect 14924 32510 14926 32562
rect 14926 32510 14978 32562
rect 14978 32510 14980 32562
rect 14924 32508 14980 32510
rect 15484 36876 15540 36932
rect 15372 36706 15428 36708
rect 15372 36654 15374 36706
rect 15374 36654 15426 36706
rect 15426 36654 15428 36706
rect 15372 36652 15428 36654
rect 15372 36258 15428 36260
rect 15372 36206 15374 36258
rect 15374 36206 15426 36258
rect 15426 36206 15428 36258
rect 15372 36204 15428 36206
rect 15260 35698 15316 35700
rect 15260 35646 15262 35698
rect 15262 35646 15314 35698
rect 15314 35646 15316 35698
rect 15260 35644 15316 35646
rect 15820 38274 15876 38276
rect 15820 38222 15822 38274
rect 15822 38222 15874 38274
rect 15874 38222 15876 38274
rect 15820 38220 15876 38222
rect 16380 39004 16436 39060
rect 16828 39452 16884 39508
rect 16940 39340 16996 39396
rect 16492 38892 16548 38948
rect 16268 38332 16324 38388
rect 16380 38108 16436 38164
rect 16268 37548 16324 37604
rect 15932 37490 15988 37492
rect 15932 37438 15934 37490
rect 15934 37438 15986 37490
rect 15986 37438 15988 37490
rect 15932 37436 15988 37438
rect 15820 36428 15876 36484
rect 16044 36258 16100 36260
rect 16044 36206 16046 36258
rect 16046 36206 16098 36258
rect 16098 36206 16100 36258
rect 16044 36204 16100 36206
rect 15372 34636 15428 34692
rect 15484 34748 15540 34804
rect 15260 34524 15316 34580
rect 15708 34802 15764 34804
rect 15708 34750 15710 34802
rect 15710 34750 15762 34802
rect 15762 34750 15764 34802
rect 15708 34748 15764 34750
rect 16268 34748 16324 34804
rect 15820 34690 15876 34692
rect 15820 34638 15822 34690
rect 15822 34638 15874 34690
rect 15874 34638 15876 34690
rect 15820 34636 15876 34638
rect 15596 33516 15652 33572
rect 15708 34412 15764 34468
rect 15708 33628 15764 33684
rect 14140 31724 14196 31780
rect 14028 31554 14084 31556
rect 14028 31502 14030 31554
rect 14030 31502 14082 31554
rect 14082 31502 14084 31554
rect 14028 31500 14084 31502
rect 13804 31164 13860 31220
rect 14140 30994 14196 30996
rect 14140 30942 14142 30994
rect 14142 30942 14194 30994
rect 14194 30942 14196 30994
rect 14140 30940 14196 30942
rect 13916 29596 13972 29652
rect 13468 24946 13524 24948
rect 13468 24894 13470 24946
rect 13470 24894 13522 24946
rect 13522 24894 13524 24946
rect 13468 24892 13524 24894
rect 13580 26124 13636 26180
rect 13468 24668 13524 24724
rect 13468 24332 13524 24388
rect 13580 23996 13636 24052
rect 13692 25564 13748 25620
rect 13468 20860 13524 20916
rect 13580 21084 13636 21140
rect 13356 20748 13412 20804
rect 13132 20018 13188 20020
rect 13132 19966 13134 20018
rect 13134 19966 13186 20018
rect 13186 19966 13188 20018
rect 13132 19964 13188 19966
rect 13244 19404 13300 19460
rect 13356 20076 13412 20132
rect 13244 18732 13300 18788
rect 11788 17052 11844 17108
rect 11900 16044 11956 16100
rect 11452 15986 11508 15988
rect 11452 15934 11454 15986
rect 11454 15934 11506 15986
rect 11506 15934 11508 15986
rect 11452 15932 11508 15934
rect 11676 15538 11732 15540
rect 11676 15486 11678 15538
rect 11678 15486 11730 15538
rect 11730 15486 11732 15538
rect 11676 15484 11732 15486
rect 9548 13356 9604 13412
rect 8092 11676 8148 11732
rect 7532 11394 7588 11396
rect 7532 11342 7534 11394
rect 7534 11342 7586 11394
rect 7586 11342 7588 11394
rect 7532 11340 7588 11342
rect 7756 10892 7812 10948
rect 6972 10610 7028 10612
rect 6972 10558 6974 10610
rect 6974 10558 7026 10610
rect 7026 10558 7028 10610
rect 6972 10556 7028 10558
rect 6972 9938 7028 9940
rect 6972 9886 6974 9938
rect 6974 9886 7026 9938
rect 7026 9886 7028 9938
rect 6972 9884 7028 9886
rect 7420 9938 7476 9940
rect 7420 9886 7422 9938
rect 7422 9886 7474 9938
rect 7474 9886 7476 9938
rect 7420 9884 7476 9886
rect 8316 12012 8372 12068
rect 9660 12066 9716 12068
rect 9660 12014 9662 12066
rect 9662 12014 9714 12066
rect 9714 12014 9716 12066
rect 9660 12012 9716 12014
rect 8876 11900 8932 11956
rect 8764 11228 8820 11284
rect 8764 10668 8820 10724
rect 8092 9884 8148 9940
rect 9548 9884 9604 9940
rect 7756 9772 7812 9828
rect 10220 15090 10276 15092
rect 10220 15038 10222 15090
rect 10222 15038 10274 15090
rect 10274 15038 10276 15090
rect 10220 15036 10276 15038
rect 11116 15036 11172 15092
rect 9996 14700 10052 14756
rect 10892 14642 10948 14644
rect 10892 14590 10894 14642
rect 10894 14590 10946 14642
rect 10946 14590 10948 14642
rect 10892 14588 10948 14590
rect 9996 14306 10052 14308
rect 9996 14254 9998 14306
rect 9998 14254 10050 14306
rect 10050 14254 10052 14306
rect 9996 14252 10052 14254
rect 9996 13916 10052 13972
rect 10444 13916 10500 13972
rect 10556 12402 10612 12404
rect 10556 12350 10558 12402
rect 10558 12350 10610 12402
rect 10610 12350 10612 12402
rect 10556 12348 10612 12350
rect 10108 11676 10164 11732
rect 10444 11900 10500 11956
rect 10668 11788 10724 11844
rect 11004 14028 11060 14084
rect 10892 13020 10948 13076
rect 10892 11900 10948 11956
rect 9996 10780 10052 10836
rect 9996 9548 10052 9604
rect 10668 11340 10724 11396
rect 10892 11282 10948 11284
rect 10892 11230 10894 11282
rect 10894 11230 10946 11282
rect 10946 11230 10948 11282
rect 10892 11228 10948 11230
rect 11004 11116 11060 11172
rect 11340 15314 11396 15316
rect 11340 15262 11342 15314
rect 11342 15262 11394 15314
rect 11394 15262 11396 15314
rect 11340 15260 11396 15262
rect 11900 15260 11956 15316
rect 11788 15148 11844 15204
rect 11228 13020 11284 13076
rect 11228 12402 11284 12404
rect 11228 12350 11230 12402
rect 11230 12350 11282 12402
rect 11282 12350 11284 12402
rect 11228 12348 11284 12350
rect 11900 14252 11956 14308
rect 11900 14028 11956 14084
rect 11676 12236 11732 12292
rect 12572 16156 12628 16212
rect 12460 15708 12516 15764
rect 12460 14476 12516 14532
rect 13020 16604 13076 16660
rect 12908 16044 12964 16100
rect 13132 15708 13188 15764
rect 12684 15202 12740 15204
rect 12684 15150 12686 15202
rect 12686 15150 12738 15202
rect 12738 15150 12740 15202
rect 12684 15148 12740 15150
rect 12348 14306 12404 14308
rect 12348 14254 12350 14306
rect 12350 14254 12402 14306
rect 12402 14254 12404 14306
rect 12348 14252 12404 14254
rect 13132 12684 13188 12740
rect 12908 11788 12964 11844
rect 9884 8316 9940 8372
rect 10556 8764 10612 8820
rect 9436 8092 9492 8148
rect 7868 7980 7924 8036
rect 7084 6690 7140 6692
rect 7084 6638 7086 6690
rect 7086 6638 7138 6690
rect 7138 6638 7140 6690
rect 7084 6636 7140 6638
rect 9884 8034 9940 8036
rect 9884 7982 9886 8034
rect 9886 7982 9938 8034
rect 9938 7982 9940 8034
rect 9884 7980 9940 7982
rect 9772 7644 9828 7700
rect 9996 7420 10052 7476
rect 8092 6636 8148 6692
rect 8876 6412 8932 6468
rect 10668 8316 10724 8372
rect 10332 7980 10388 8036
rect 10220 7698 10276 7700
rect 10220 7646 10222 7698
rect 10222 7646 10274 7698
rect 10274 7646 10276 7698
rect 10220 7644 10276 7646
rect 10220 6636 10276 6692
rect 11116 8652 11172 8708
rect 11900 11676 11956 11732
rect 12012 11228 12068 11284
rect 12348 11282 12404 11284
rect 12348 11230 12350 11282
rect 12350 11230 12402 11282
rect 12402 11230 12404 11282
rect 12348 11228 12404 11230
rect 11564 11116 11620 11172
rect 10780 8204 10836 8260
rect 10780 7868 10836 7924
rect 11004 8034 11060 8036
rect 11004 7982 11006 8034
rect 11006 7982 11058 8034
rect 11058 7982 11060 8034
rect 11004 7980 11060 7982
rect 10444 7698 10500 7700
rect 10444 7646 10446 7698
rect 10446 7646 10498 7698
rect 10498 7646 10500 7698
rect 10444 7644 10500 7646
rect 11004 7362 11060 7364
rect 11004 7310 11006 7362
rect 11006 7310 11058 7362
rect 11058 7310 11060 7362
rect 11004 7308 11060 7310
rect 11788 9436 11844 9492
rect 11564 8258 11620 8260
rect 11564 8206 11566 8258
rect 11566 8206 11618 8258
rect 11618 8206 11620 8258
rect 11564 8204 11620 8206
rect 13020 9884 13076 9940
rect 12012 8764 12068 8820
rect 11788 7644 11844 7700
rect 13020 8316 13076 8372
rect 12908 8258 12964 8260
rect 12908 8206 12910 8258
rect 12910 8206 12962 8258
rect 12962 8206 12964 8258
rect 12908 8204 12964 8206
rect 12348 8146 12404 8148
rect 12348 8094 12350 8146
rect 12350 8094 12402 8146
rect 12402 8094 12404 8146
rect 12348 8092 12404 8094
rect 12796 8146 12852 8148
rect 12796 8094 12798 8146
rect 12798 8094 12850 8146
rect 12850 8094 12852 8146
rect 12796 8092 12852 8094
rect 12012 7980 12068 8036
rect 11452 7196 11508 7252
rect 11676 7308 11732 7364
rect 11452 6690 11508 6692
rect 11452 6638 11454 6690
rect 11454 6638 11506 6690
rect 11506 6638 11508 6690
rect 11452 6636 11508 6638
rect 10668 6466 10724 6468
rect 10668 6414 10670 6466
rect 10670 6414 10722 6466
rect 10722 6414 10724 6466
rect 10668 6412 10724 6414
rect 11340 6466 11396 6468
rect 11340 6414 11342 6466
rect 11342 6414 11394 6466
rect 11394 6414 11396 6466
rect 11340 6412 11396 6414
rect 10220 5852 10276 5908
rect 10556 5852 10612 5908
rect 10108 4508 10164 4564
rect 10220 5180 10276 5236
rect 10892 5906 10948 5908
rect 10892 5854 10894 5906
rect 10894 5854 10946 5906
rect 10946 5854 10948 5906
rect 10892 5852 10948 5854
rect 12460 7362 12516 7364
rect 12460 7310 12462 7362
rect 12462 7310 12514 7362
rect 12514 7310 12516 7362
rect 12460 7308 12516 7310
rect 11900 6860 11956 6916
rect 13916 24780 13972 24836
rect 13916 24444 13972 24500
rect 14476 31724 14532 31780
rect 14924 31554 14980 31556
rect 14924 31502 14926 31554
rect 14926 31502 14978 31554
rect 14978 31502 14980 31554
rect 14924 31500 14980 31502
rect 14476 31052 14532 31108
rect 15596 32956 15652 33012
rect 15372 31778 15428 31780
rect 15372 31726 15374 31778
rect 15374 31726 15426 31778
rect 15426 31726 15428 31778
rect 15372 31724 15428 31726
rect 15372 30828 15428 30884
rect 14140 26684 14196 26740
rect 14252 21868 14308 21924
rect 14476 27468 14532 27524
rect 15148 29372 15204 29428
rect 16380 34076 16436 34132
rect 15708 31724 15764 31780
rect 15708 31388 15764 31444
rect 16156 31554 16212 31556
rect 16156 31502 16158 31554
rect 16158 31502 16210 31554
rect 16210 31502 16212 31554
rect 16156 31500 16212 31502
rect 16492 33346 16548 33348
rect 16492 33294 16494 33346
rect 16494 33294 16546 33346
rect 16546 33294 16548 33346
rect 16492 33292 16548 33294
rect 16940 37772 16996 37828
rect 16828 36482 16884 36484
rect 16828 36430 16830 36482
rect 16830 36430 16882 36482
rect 16882 36430 16884 36482
rect 16828 36428 16884 36430
rect 16940 36316 16996 36372
rect 16940 34914 16996 34916
rect 16940 34862 16942 34914
rect 16942 34862 16994 34914
rect 16994 34862 16996 34914
rect 16940 34860 16996 34862
rect 16828 33516 16884 33572
rect 16940 33180 16996 33236
rect 17388 39394 17444 39396
rect 17388 39342 17390 39394
rect 17390 39342 17442 39394
rect 17442 39342 17444 39394
rect 17388 39340 17444 39342
rect 17724 39340 17780 39396
rect 17164 38332 17220 38388
rect 17276 38108 17332 38164
rect 17500 38108 17556 38164
rect 17388 37826 17444 37828
rect 17388 37774 17390 37826
rect 17390 37774 17442 37826
rect 17442 37774 17444 37826
rect 17388 37772 17444 37774
rect 18172 39340 18228 39396
rect 17612 37938 17668 37940
rect 17612 37886 17614 37938
rect 17614 37886 17666 37938
rect 17666 37886 17668 37938
rect 17612 37884 17668 37886
rect 18060 37884 18116 37940
rect 18060 37378 18116 37380
rect 18060 37326 18062 37378
rect 18062 37326 18114 37378
rect 18114 37326 18116 37378
rect 18060 37324 18116 37326
rect 17724 37266 17780 37268
rect 17724 37214 17726 37266
rect 17726 37214 17778 37266
rect 17778 37214 17780 37266
rect 17724 37212 17780 37214
rect 17500 36988 17556 37044
rect 17948 36876 18004 36932
rect 18620 38834 18676 38836
rect 18620 38782 18622 38834
rect 18622 38782 18674 38834
rect 18674 38782 18676 38834
rect 18620 38780 18676 38782
rect 18396 37266 18452 37268
rect 18396 37214 18398 37266
rect 18398 37214 18450 37266
rect 18450 37214 18452 37266
rect 18396 37212 18452 37214
rect 17948 36316 18004 36372
rect 17612 34748 17668 34804
rect 17948 34748 18004 34804
rect 17388 33628 17444 33684
rect 17052 32956 17108 33012
rect 17500 33180 17556 33236
rect 16940 32508 16996 32564
rect 16716 32396 16772 32452
rect 16492 31388 16548 31444
rect 16156 30882 16212 30884
rect 16156 30830 16158 30882
rect 16158 30830 16210 30882
rect 16210 30830 16212 30882
rect 16156 30828 16212 30830
rect 16268 30716 16324 30772
rect 15820 30156 15876 30212
rect 15932 30380 15988 30436
rect 15260 28364 15316 28420
rect 15148 27804 15204 27860
rect 15260 27244 15316 27300
rect 14812 27132 14868 27188
rect 14476 26684 14532 26740
rect 15820 28588 15876 28644
rect 15596 28418 15652 28420
rect 15596 28366 15598 28418
rect 15598 28366 15650 28418
rect 15650 28366 15652 28418
rect 15596 28364 15652 28366
rect 15932 28418 15988 28420
rect 15932 28366 15934 28418
rect 15934 28366 15986 28418
rect 15986 28366 15988 28418
rect 15932 28364 15988 28366
rect 16268 29932 16324 29988
rect 16380 28700 16436 28756
rect 16268 28530 16324 28532
rect 16268 28478 16270 28530
rect 16270 28478 16322 28530
rect 16322 28478 16324 28530
rect 16268 28476 16324 28478
rect 16268 28252 16324 28308
rect 16380 28140 16436 28196
rect 15372 26684 15428 26740
rect 15596 27132 15652 27188
rect 15932 27074 15988 27076
rect 15932 27022 15934 27074
rect 15934 27022 15986 27074
rect 15986 27022 15988 27074
rect 15932 27020 15988 27022
rect 18172 36370 18228 36372
rect 18172 36318 18174 36370
rect 18174 36318 18226 36370
rect 18226 36318 18228 36370
rect 18172 36316 18228 36318
rect 18284 36258 18340 36260
rect 18284 36206 18286 36258
rect 18286 36206 18338 36258
rect 18338 36206 18340 36258
rect 18284 36204 18340 36206
rect 18732 34972 18788 35028
rect 18732 34354 18788 34356
rect 18732 34302 18734 34354
rect 18734 34302 18786 34354
rect 18786 34302 18788 34354
rect 18732 34300 18788 34302
rect 19068 38780 19124 38836
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19628 40348 19684 40404
rect 20748 40348 20804 40404
rect 22764 41132 22820 41188
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19516 38722 19572 38724
rect 19516 38670 19518 38722
rect 19518 38670 19570 38722
rect 19570 38670 19572 38722
rect 19516 38668 19572 38670
rect 19068 36316 19124 36372
rect 18844 33292 18900 33348
rect 18956 36258 19012 36260
rect 18956 36206 18958 36258
rect 18958 36206 19010 36258
rect 19010 36206 19012 36258
rect 18956 36204 19012 36206
rect 18060 32562 18116 32564
rect 18060 32510 18062 32562
rect 18062 32510 18114 32562
rect 18114 32510 18116 32562
rect 18060 32508 18116 32510
rect 17052 31500 17108 31556
rect 17276 31052 17332 31108
rect 16940 30210 16996 30212
rect 16940 30158 16942 30210
rect 16942 30158 16994 30210
rect 16994 30158 16996 30210
rect 16940 30156 16996 30158
rect 17052 29932 17108 29988
rect 16604 29426 16660 29428
rect 16604 29374 16606 29426
rect 16606 29374 16658 29426
rect 16658 29374 16660 29426
rect 16604 29372 16660 29374
rect 17052 29484 17108 29540
rect 16940 29426 16996 29428
rect 16940 29374 16942 29426
rect 16942 29374 16994 29426
rect 16994 29374 16996 29426
rect 16940 29372 16996 29374
rect 16604 28418 16660 28420
rect 16604 28366 16606 28418
rect 16606 28366 16658 28418
rect 16658 28366 16660 28418
rect 16604 28364 16660 28366
rect 15708 26908 15764 26964
rect 16156 26908 16212 26964
rect 16716 27186 16772 27188
rect 16716 27134 16718 27186
rect 16718 27134 16770 27186
rect 16770 27134 16772 27186
rect 16716 27132 16772 27134
rect 17724 30268 17780 30324
rect 17388 29708 17444 29764
rect 18060 29932 18116 29988
rect 17612 29820 17668 29876
rect 17500 29596 17556 29652
rect 17836 29538 17892 29540
rect 17836 29486 17838 29538
rect 17838 29486 17890 29538
rect 17890 29486 17892 29538
rect 17836 29484 17892 29486
rect 18060 29538 18116 29540
rect 18060 29486 18062 29538
rect 18062 29486 18114 29538
rect 18114 29486 18116 29538
rect 18060 29484 18116 29486
rect 17612 29260 17668 29316
rect 17948 29148 18004 29204
rect 17388 28642 17444 28644
rect 17388 28590 17390 28642
rect 17390 28590 17442 28642
rect 17442 28590 17444 28642
rect 17388 28588 17444 28590
rect 18620 32562 18676 32564
rect 18620 32510 18622 32562
rect 18622 32510 18674 32562
rect 18674 32510 18676 32562
rect 18620 32508 18676 32510
rect 18396 29986 18452 29988
rect 18396 29934 18398 29986
rect 18398 29934 18450 29986
rect 18450 29934 18452 29986
rect 18396 29932 18452 29934
rect 18508 29314 18564 29316
rect 18508 29262 18510 29314
rect 18510 29262 18562 29314
rect 18562 29262 18564 29314
rect 18508 29260 18564 29262
rect 18508 29036 18564 29092
rect 18284 28642 18340 28644
rect 18284 28590 18286 28642
rect 18286 28590 18338 28642
rect 18338 28590 18340 28642
rect 18284 28588 18340 28590
rect 17276 28140 17332 28196
rect 18060 27916 18116 27972
rect 17612 27692 17668 27748
rect 15932 26572 15988 26628
rect 15820 26402 15876 26404
rect 15820 26350 15822 26402
rect 15822 26350 15874 26402
rect 15874 26350 15876 26402
rect 15820 26348 15876 26350
rect 15596 26236 15652 26292
rect 15820 26124 15876 26180
rect 14924 25004 14980 25060
rect 15484 25004 15540 25060
rect 15260 24946 15316 24948
rect 15260 24894 15262 24946
rect 15262 24894 15314 24946
rect 15314 24894 15316 24946
rect 15260 24892 15316 24894
rect 14812 24722 14868 24724
rect 14812 24670 14814 24722
rect 14814 24670 14866 24722
rect 14866 24670 14868 24722
rect 14812 24668 14868 24670
rect 14476 22764 14532 22820
rect 14700 22540 14756 22596
rect 14476 21644 14532 21700
rect 14588 22204 14644 22260
rect 14588 21868 14644 21924
rect 14364 21420 14420 21476
rect 13804 20188 13860 20244
rect 13916 20130 13972 20132
rect 13916 20078 13918 20130
rect 13918 20078 13970 20130
rect 13970 20078 13972 20130
rect 13916 20076 13972 20078
rect 13692 19404 13748 19460
rect 13804 19740 13860 19796
rect 13580 19234 13636 19236
rect 13580 19182 13582 19234
rect 13582 19182 13634 19234
rect 13634 19182 13636 19234
rect 13580 19180 13636 19182
rect 13692 18844 13748 18900
rect 13468 18396 13524 18452
rect 13916 19292 13972 19348
rect 14476 20578 14532 20580
rect 14476 20526 14478 20578
rect 14478 20526 14530 20578
rect 14530 20526 14532 20578
rect 14476 20524 14532 20526
rect 14364 20076 14420 20132
rect 14028 18620 14084 18676
rect 14252 18450 14308 18452
rect 14252 18398 14254 18450
rect 14254 18398 14306 18450
rect 14306 18398 14308 18450
rect 14252 18396 14308 18398
rect 15148 23436 15204 23492
rect 15148 22764 15204 22820
rect 15036 22428 15092 22484
rect 14924 22258 14980 22260
rect 14924 22206 14926 22258
rect 14926 22206 14978 22258
rect 14978 22206 14980 22258
rect 14924 22204 14980 22206
rect 14812 21644 14868 21700
rect 14924 21420 14980 21476
rect 14812 20748 14868 20804
rect 14924 19964 14980 20020
rect 14700 19740 14756 19796
rect 14700 19404 14756 19460
rect 14364 17948 14420 18004
rect 13356 16770 13412 16772
rect 13356 16718 13358 16770
rect 13358 16718 13410 16770
rect 13410 16718 13412 16770
rect 13356 16716 13412 16718
rect 13580 17442 13636 17444
rect 13580 17390 13582 17442
rect 13582 17390 13634 17442
rect 13634 17390 13636 17442
rect 13580 17388 13636 17390
rect 13356 14476 13412 14532
rect 13692 17106 13748 17108
rect 13692 17054 13694 17106
rect 13694 17054 13746 17106
rect 13746 17054 13748 17106
rect 13692 17052 13748 17054
rect 14140 16098 14196 16100
rect 14140 16046 14142 16098
rect 14142 16046 14194 16098
rect 14194 16046 14196 16098
rect 14140 16044 14196 16046
rect 13580 14364 13636 14420
rect 13692 12684 13748 12740
rect 13916 14530 13972 14532
rect 13916 14478 13918 14530
rect 13918 14478 13970 14530
rect 13970 14478 13972 14530
rect 13916 14476 13972 14478
rect 15260 21196 15316 21252
rect 15260 20018 15316 20020
rect 15260 19966 15262 20018
rect 15262 19966 15314 20018
rect 15314 19966 15316 20018
rect 15260 19964 15316 19966
rect 15036 19346 15092 19348
rect 15036 19294 15038 19346
rect 15038 19294 15090 19346
rect 15090 19294 15092 19346
rect 15036 19292 15092 19294
rect 14700 18508 14756 18564
rect 14812 19180 14868 19236
rect 14700 16828 14756 16884
rect 14700 14754 14756 14756
rect 14700 14702 14702 14754
rect 14702 14702 14754 14754
rect 14754 14702 14756 14754
rect 14700 14700 14756 14702
rect 15596 21474 15652 21476
rect 15596 21422 15598 21474
rect 15598 21422 15650 21474
rect 15650 21422 15652 21474
rect 15596 21420 15652 21422
rect 16268 26514 16324 26516
rect 16268 26462 16270 26514
rect 16270 26462 16322 26514
rect 16322 26462 16324 26514
rect 16268 26460 16324 26462
rect 16604 26460 16660 26516
rect 16380 26402 16436 26404
rect 16380 26350 16382 26402
rect 16382 26350 16434 26402
rect 16434 26350 16436 26402
rect 16380 26348 16436 26350
rect 16268 26236 16324 26292
rect 16828 25676 16884 25732
rect 16940 25788 16996 25844
rect 16492 25282 16548 25284
rect 16492 25230 16494 25282
rect 16494 25230 16546 25282
rect 16546 25230 16548 25282
rect 16492 25228 16548 25230
rect 16604 24946 16660 24948
rect 16604 24894 16606 24946
rect 16606 24894 16658 24946
rect 16658 24894 16660 24946
rect 16604 24892 16660 24894
rect 16380 24722 16436 24724
rect 16380 24670 16382 24722
rect 16382 24670 16434 24722
rect 16434 24670 16436 24722
rect 16380 24668 16436 24670
rect 16492 24610 16548 24612
rect 16492 24558 16494 24610
rect 16494 24558 16546 24610
rect 16546 24558 16548 24610
rect 16492 24556 16548 24558
rect 16492 24050 16548 24052
rect 16492 23998 16494 24050
rect 16494 23998 16546 24050
rect 16546 23998 16548 24050
rect 16492 23996 16548 23998
rect 16044 22092 16100 22148
rect 17052 25282 17108 25284
rect 17052 25230 17054 25282
rect 17054 25230 17106 25282
rect 17106 25230 17108 25282
rect 17052 25228 17108 25230
rect 17164 24892 17220 24948
rect 17164 23938 17220 23940
rect 17164 23886 17166 23938
rect 17166 23886 17218 23938
rect 17218 23886 17220 23938
rect 17164 23884 17220 23886
rect 16828 23826 16884 23828
rect 16828 23774 16830 23826
rect 16830 23774 16882 23826
rect 16882 23774 16884 23826
rect 16828 23772 16884 23774
rect 16716 23436 16772 23492
rect 16604 23212 16660 23268
rect 15932 21756 15988 21812
rect 16492 22092 16548 22148
rect 15372 19068 15428 19124
rect 15596 20860 15652 20916
rect 15708 20802 15764 20804
rect 15708 20750 15710 20802
rect 15710 20750 15762 20802
rect 15762 20750 15764 20802
rect 15708 20748 15764 20750
rect 15708 19852 15764 19908
rect 15708 19010 15764 19012
rect 15708 18958 15710 19010
rect 15710 18958 15762 19010
rect 15762 18958 15764 19010
rect 15708 18956 15764 18958
rect 14924 16882 14980 16884
rect 14924 16830 14926 16882
rect 14926 16830 14978 16882
rect 14978 16830 14980 16882
rect 14924 16828 14980 16830
rect 15148 16716 15204 16772
rect 14924 16492 14980 16548
rect 15932 20972 15988 21028
rect 16268 20972 16324 21028
rect 17388 25900 17444 25956
rect 17500 25676 17556 25732
rect 17724 26460 17780 26516
rect 18060 26402 18116 26404
rect 18060 26350 18062 26402
rect 18062 26350 18114 26402
rect 18114 26350 18116 26402
rect 18060 26348 18116 26350
rect 17724 25564 17780 25620
rect 17612 24946 17668 24948
rect 17612 24894 17614 24946
rect 17614 24894 17666 24946
rect 17666 24894 17668 24946
rect 17612 24892 17668 24894
rect 17724 25228 17780 25284
rect 17500 24668 17556 24724
rect 17500 23996 17556 24052
rect 17500 23436 17556 23492
rect 17612 23212 17668 23268
rect 17388 21868 17444 21924
rect 17612 21868 17668 21924
rect 16828 21474 16884 21476
rect 16828 21422 16830 21474
rect 16830 21422 16882 21474
rect 16882 21422 16884 21474
rect 16828 21420 16884 21422
rect 17500 21420 17556 21476
rect 17612 21362 17668 21364
rect 17612 21310 17614 21362
rect 17614 21310 17666 21362
rect 17666 21310 17668 21362
rect 17612 21308 17668 21310
rect 17388 21084 17444 21140
rect 16044 20018 16100 20020
rect 16044 19966 16046 20018
rect 16046 19966 16098 20018
rect 16098 19966 16100 20018
rect 16044 19964 16100 19966
rect 16044 18732 16100 18788
rect 15820 18620 15876 18676
rect 17164 20636 17220 20692
rect 15484 18508 15540 18564
rect 15708 18060 15764 18116
rect 15372 15708 15428 15764
rect 15596 15426 15652 15428
rect 15596 15374 15598 15426
rect 15598 15374 15650 15426
rect 15650 15374 15652 15426
rect 15596 15372 15652 15374
rect 14476 14252 14532 14308
rect 14588 14588 14644 14644
rect 14812 14530 14868 14532
rect 14812 14478 14814 14530
rect 14814 14478 14866 14530
rect 14866 14478 14868 14530
rect 14812 14476 14868 14478
rect 14700 14418 14756 14420
rect 14700 14366 14702 14418
rect 14702 14366 14754 14418
rect 14754 14366 14756 14418
rect 14700 14364 14756 14366
rect 14700 13244 14756 13300
rect 13916 12178 13972 12180
rect 13916 12126 13918 12178
rect 13918 12126 13970 12178
rect 13970 12126 13972 12178
rect 13916 12124 13972 12126
rect 13692 11340 13748 11396
rect 13692 10668 13748 10724
rect 13580 9938 13636 9940
rect 13580 9886 13582 9938
rect 13582 9886 13634 9938
rect 13634 9886 13636 9938
rect 13580 9884 13636 9886
rect 13356 9436 13412 9492
rect 13356 8316 13412 8372
rect 13468 8258 13524 8260
rect 13468 8206 13470 8258
rect 13470 8206 13522 8258
rect 13522 8206 13524 8258
rect 13468 8204 13524 8206
rect 13580 8034 13636 8036
rect 13580 7982 13582 8034
rect 13582 7982 13634 8034
rect 13634 7982 13636 8034
rect 13580 7980 13636 7982
rect 13356 7084 13412 7140
rect 13244 6860 13300 6916
rect 12684 6690 12740 6692
rect 12684 6638 12686 6690
rect 12686 6638 12738 6690
rect 12738 6638 12740 6690
rect 12684 6636 12740 6638
rect 12796 6578 12852 6580
rect 12796 6526 12798 6578
rect 12798 6526 12850 6578
rect 12850 6526 12852 6578
rect 12796 6524 12852 6526
rect 11900 6412 11956 6468
rect 11004 5234 11060 5236
rect 11004 5182 11006 5234
rect 11006 5182 11058 5234
rect 11058 5182 11060 5234
rect 11004 5180 11060 5182
rect 11788 5180 11844 5236
rect 12684 5234 12740 5236
rect 12684 5182 12686 5234
rect 12686 5182 12738 5234
rect 12738 5182 12740 5234
rect 12684 5180 12740 5182
rect 6300 4060 6356 4116
rect 7420 4114 7476 4116
rect 7420 4062 7422 4114
rect 7422 4062 7474 4114
rect 7474 4062 7476 4114
rect 7420 4060 7476 4062
rect 8764 3554 8820 3556
rect 8764 3502 8766 3554
rect 8766 3502 8818 3554
rect 8818 3502 8820 3554
rect 8764 3500 8820 3502
rect 14028 11228 14084 11284
rect 14252 12796 14308 12852
rect 14140 8316 14196 8372
rect 14476 11340 14532 11396
rect 14364 8092 14420 8148
rect 13916 7084 13972 7140
rect 13692 6524 13748 6580
rect 13804 6466 13860 6468
rect 13804 6414 13806 6466
rect 13806 6414 13858 6466
rect 13858 6414 13860 6466
rect 13804 6412 13860 6414
rect 13468 4060 13524 4116
rect 14140 7420 14196 7476
rect 14700 12124 14756 12180
rect 15260 14364 15316 14420
rect 15260 13468 15316 13524
rect 15596 12908 15652 12964
rect 15036 12850 15092 12852
rect 15036 12798 15038 12850
rect 15038 12798 15090 12850
rect 15090 12798 15092 12850
rect 15036 12796 15092 12798
rect 16828 19906 16884 19908
rect 16828 19854 16830 19906
rect 16830 19854 16882 19906
rect 16882 19854 16884 19906
rect 16828 19852 16884 19854
rect 16268 18396 16324 18452
rect 16492 18732 16548 18788
rect 16156 17500 16212 17556
rect 16268 16716 16324 16772
rect 16268 15708 16324 15764
rect 16940 19010 16996 19012
rect 16940 18958 16942 19010
rect 16942 18958 16994 19010
rect 16994 18958 16996 19010
rect 16940 18956 16996 18958
rect 16716 18172 16772 18228
rect 17612 21084 17668 21140
rect 17500 20748 17556 20804
rect 17500 19740 17556 19796
rect 17612 18956 17668 19012
rect 16940 17836 16996 17892
rect 17948 23884 18004 23940
rect 17836 23714 17892 23716
rect 17836 23662 17838 23714
rect 17838 23662 17890 23714
rect 17890 23662 17892 23714
rect 17836 23660 17892 23662
rect 17836 21644 17892 21700
rect 17836 20802 17892 20804
rect 17836 20750 17838 20802
rect 17838 20750 17890 20802
rect 17890 20750 17892 20802
rect 17836 20748 17892 20750
rect 18284 22988 18340 23044
rect 18396 23324 18452 23380
rect 18172 21868 18228 21924
rect 18172 19068 18228 19124
rect 17164 18396 17220 18452
rect 17388 18450 17444 18452
rect 17388 18398 17390 18450
rect 17390 18398 17442 18450
rect 17442 18398 17444 18450
rect 17388 18396 17444 18398
rect 17948 18844 18004 18900
rect 17500 18060 17556 18116
rect 17948 18284 18004 18340
rect 17388 17666 17444 17668
rect 17388 17614 17390 17666
rect 17390 17614 17442 17666
rect 17442 17614 17444 17666
rect 17388 17612 17444 17614
rect 16716 17500 16772 17556
rect 16604 16492 16660 16548
rect 16604 16156 16660 16212
rect 16828 15148 16884 15204
rect 15820 14530 15876 14532
rect 15820 14478 15822 14530
rect 15822 14478 15874 14530
rect 15874 14478 15876 14530
rect 15820 14476 15876 14478
rect 15820 13468 15876 13524
rect 15708 12460 15764 12516
rect 15932 12236 15988 12292
rect 15260 10722 15316 10724
rect 15260 10670 15262 10722
rect 15262 10670 15314 10722
rect 15314 10670 15316 10722
rect 15260 10668 15316 10670
rect 15372 10834 15428 10836
rect 15372 10782 15374 10834
rect 15374 10782 15426 10834
rect 15426 10782 15428 10834
rect 15372 10780 15428 10782
rect 15484 10444 15540 10500
rect 15148 9772 15204 9828
rect 14700 9324 14756 9380
rect 15372 9266 15428 9268
rect 15372 9214 15374 9266
rect 15374 9214 15426 9266
rect 15426 9214 15428 9266
rect 15372 9212 15428 9214
rect 15036 8876 15092 8932
rect 15036 8092 15092 8148
rect 15484 7980 15540 8036
rect 15372 7698 15428 7700
rect 15372 7646 15374 7698
rect 15374 7646 15426 7698
rect 15426 7646 15428 7698
rect 15372 7644 15428 7646
rect 15708 9548 15764 9604
rect 16604 13468 16660 13524
rect 17836 17890 17892 17892
rect 17836 17838 17838 17890
rect 17838 17838 17890 17890
rect 17890 17838 17892 17890
rect 17836 17836 17892 17838
rect 16940 13356 16996 13412
rect 17052 17052 17108 17108
rect 16716 13020 16772 13076
rect 19068 35644 19124 35700
rect 20188 38220 20244 38276
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19516 37378 19572 37380
rect 19516 37326 19518 37378
rect 19518 37326 19570 37378
rect 19570 37326 19572 37378
rect 19516 37324 19572 37326
rect 20076 37324 20132 37380
rect 19628 36092 19684 36148
rect 19180 33964 19236 34020
rect 19068 33234 19124 33236
rect 19068 33182 19070 33234
rect 19070 33182 19122 33234
rect 19122 33182 19124 33234
rect 19068 33180 19124 33182
rect 19068 29538 19124 29540
rect 19068 29486 19070 29538
rect 19070 29486 19122 29538
rect 19122 29486 19124 29538
rect 19068 29484 19124 29486
rect 18956 29036 19012 29092
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20300 36370 20356 36372
rect 20300 36318 20302 36370
rect 20302 36318 20354 36370
rect 20354 36318 20356 36370
rect 20300 36316 20356 36318
rect 20188 34802 20244 34804
rect 20188 34750 20190 34802
rect 20190 34750 20242 34802
rect 20242 34750 20244 34802
rect 20188 34748 20244 34750
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 21644 39564 21700 39620
rect 20748 38162 20804 38164
rect 20748 38110 20750 38162
rect 20750 38110 20802 38162
rect 20802 38110 20804 38162
rect 20748 38108 20804 38110
rect 20636 36204 20692 36260
rect 22428 39506 22484 39508
rect 22428 39454 22430 39506
rect 22430 39454 22482 39506
rect 22482 39454 22484 39506
rect 22428 39452 22484 39454
rect 23996 41356 24052 41412
rect 24556 41186 24612 41188
rect 24556 41134 24558 41186
rect 24558 41134 24610 41186
rect 24610 41134 24612 41186
rect 24556 41132 24612 41134
rect 25564 41410 25620 41412
rect 25564 41358 25566 41410
rect 25566 41358 25618 41410
rect 25618 41358 25620 41410
rect 25564 41356 25620 41358
rect 26236 41356 26292 41412
rect 25116 40572 25172 40628
rect 26348 40626 26404 40628
rect 26348 40574 26350 40626
rect 26350 40574 26402 40626
rect 26402 40574 26404 40626
rect 26348 40572 26404 40574
rect 27356 40572 27412 40628
rect 27468 41132 27524 41188
rect 24668 40514 24724 40516
rect 24668 40462 24670 40514
rect 24670 40462 24722 40514
rect 24722 40462 24724 40514
rect 24668 40460 24724 40462
rect 25340 40460 25396 40516
rect 22876 39788 22932 39844
rect 24108 39842 24164 39844
rect 24108 39790 24110 39842
rect 24110 39790 24162 39842
rect 24162 39790 24164 39842
rect 24108 39788 24164 39790
rect 23100 39618 23156 39620
rect 23100 39566 23102 39618
rect 23102 39566 23154 39618
rect 23154 39566 23156 39618
rect 23100 39564 23156 39566
rect 23884 39340 23940 39396
rect 24332 39004 24388 39060
rect 21868 38668 21924 38724
rect 21196 36428 21252 36484
rect 20524 35084 20580 35140
rect 20412 34524 20468 34580
rect 19516 33964 19572 34020
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19628 31836 19684 31892
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19292 31052 19348 31108
rect 20076 30434 20132 30436
rect 20076 30382 20078 30434
rect 20078 30382 20130 30434
rect 20130 30382 20132 30434
rect 20076 30380 20132 30382
rect 20300 34300 20356 34356
rect 21532 36092 21588 36148
rect 24108 38722 24164 38724
rect 24108 38670 24110 38722
rect 24110 38670 24162 38722
rect 24162 38670 24164 38722
rect 24108 38668 24164 38670
rect 26236 39730 26292 39732
rect 26236 39678 26238 39730
rect 26238 39678 26290 39730
rect 26290 39678 26292 39730
rect 26236 39676 26292 39678
rect 25788 39452 25844 39508
rect 25228 39340 25284 39396
rect 24668 39116 24724 39172
rect 25116 38668 25172 38724
rect 24668 38108 24724 38164
rect 22428 37100 22484 37156
rect 22092 36428 22148 36484
rect 20860 35756 20916 35812
rect 20860 35420 20916 35476
rect 21980 35810 22036 35812
rect 21980 35758 21982 35810
rect 21982 35758 22034 35810
rect 22034 35758 22036 35810
rect 21980 35756 22036 35758
rect 22204 36316 22260 36372
rect 21868 35084 21924 35140
rect 21980 35196 22036 35252
rect 21756 34524 21812 34580
rect 21532 33180 21588 33236
rect 20300 32172 20356 32228
rect 20300 31724 20356 31780
rect 21308 31836 21364 31892
rect 20972 31612 21028 31668
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20412 29426 20468 29428
rect 20412 29374 20414 29426
rect 20414 29374 20466 29426
rect 20466 29374 20468 29426
rect 20412 29372 20468 29374
rect 19628 29036 19684 29092
rect 18620 23938 18676 23940
rect 18620 23886 18622 23938
rect 18622 23886 18674 23938
rect 18674 23886 18676 23938
rect 18620 23884 18676 23886
rect 18396 18284 18452 18340
rect 18508 18172 18564 18228
rect 17724 17052 17780 17108
rect 17948 16994 18004 16996
rect 17948 16942 17950 16994
rect 17950 16942 18002 16994
rect 18002 16942 18004 16994
rect 17948 16940 18004 16942
rect 17612 16828 17668 16884
rect 17276 16604 17332 16660
rect 17164 15148 17220 15204
rect 17388 16380 17444 16436
rect 17612 16380 17668 16436
rect 17500 15596 17556 15652
rect 17724 15538 17780 15540
rect 17724 15486 17726 15538
rect 17726 15486 17778 15538
rect 17778 15486 17780 15538
rect 17724 15484 17780 15486
rect 18284 15874 18340 15876
rect 18284 15822 18286 15874
rect 18286 15822 18338 15874
rect 18338 15822 18340 15874
rect 18284 15820 18340 15822
rect 18284 15484 18340 15540
rect 18060 15426 18116 15428
rect 18060 15374 18062 15426
rect 18062 15374 18114 15426
rect 18114 15374 18116 15426
rect 18060 15372 18116 15374
rect 17388 15148 17444 15204
rect 18508 16940 18564 16996
rect 18508 15596 18564 15652
rect 16716 12290 16772 12292
rect 16716 12238 16718 12290
rect 16718 12238 16770 12290
rect 16770 12238 16772 12290
rect 16716 12236 16772 12238
rect 17164 13132 17220 13188
rect 16828 12178 16884 12180
rect 16828 12126 16830 12178
rect 16830 12126 16882 12178
rect 16882 12126 16884 12178
rect 16828 12124 16884 12126
rect 17724 13858 17780 13860
rect 17724 13806 17726 13858
rect 17726 13806 17778 13858
rect 17778 13806 17780 13858
rect 17724 13804 17780 13806
rect 18060 13858 18116 13860
rect 18060 13806 18062 13858
rect 18062 13806 18114 13858
rect 18114 13806 18116 13858
rect 18060 13804 18116 13806
rect 17276 12460 17332 12516
rect 17276 11116 17332 11172
rect 16940 10780 16996 10836
rect 17388 10834 17444 10836
rect 17388 10782 17390 10834
rect 17390 10782 17442 10834
rect 17442 10782 17444 10834
rect 17388 10780 17444 10782
rect 15820 9324 15876 9380
rect 17612 13132 17668 13188
rect 17612 12348 17668 12404
rect 17836 12178 17892 12180
rect 17836 12126 17838 12178
rect 17838 12126 17890 12178
rect 17890 12126 17892 12178
rect 17836 12124 17892 12126
rect 17612 10610 17668 10612
rect 17612 10558 17614 10610
rect 17614 10558 17666 10610
rect 17666 10558 17668 10610
rect 17612 10556 17668 10558
rect 18172 10780 18228 10836
rect 18844 24780 18900 24836
rect 18844 24610 18900 24612
rect 18844 24558 18846 24610
rect 18846 24558 18898 24610
rect 18898 24558 18900 24610
rect 18844 24556 18900 24558
rect 18844 20802 18900 20804
rect 18844 20750 18846 20802
rect 18846 20750 18898 20802
rect 18898 20750 18900 20802
rect 18844 20748 18900 20750
rect 18732 19180 18788 19236
rect 18732 18732 18788 18788
rect 20188 28700 20244 28756
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20636 29708 20692 29764
rect 20860 30940 20916 30996
rect 21308 30828 21364 30884
rect 20972 30380 21028 30436
rect 20748 30044 20804 30100
rect 21196 29708 21252 29764
rect 20636 28642 20692 28644
rect 20636 28590 20638 28642
rect 20638 28590 20690 28642
rect 20690 28590 20692 28642
rect 20636 28588 20692 28590
rect 20524 27074 20580 27076
rect 20524 27022 20526 27074
rect 20526 27022 20578 27074
rect 20578 27022 20580 27074
rect 20524 27020 20580 27022
rect 20188 26796 20244 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19628 26178 19684 26180
rect 19628 26126 19630 26178
rect 19630 26126 19682 26178
rect 19682 26126 19684 26178
rect 19628 26124 19684 26126
rect 20860 26236 20916 26292
rect 20636 26124 20692 26180
rect 20524 25506 20580 25508
rect 20524 25454 20526 25506
rect 20526 25454 20578 25506
rect 20578 25454 20580 25506
rect 20524 25452 20580 25454
rect 19628 25340 19684 25396
rect 20412 25340 20468 25396
rect 19068 25228 19124 25284
rect 19852 25282 19908 25284
rect 19852 25230 19854 25282
rect 19854 25230 19906 25282
rect 19906 25230 19908 25282
rect 19852 25228 19908 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20188 25116 20244 25172
rect 19292 23884 19348 23940
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20188 23436 20244 23492
rect 19292 23212 19348 23268
rect 20076 23266 20132 23268
rect 20076 23214 20078 23266
rect 20078 23214 20130 23266
rect 20130 23214 20132 23266
rect 20076 23212 20132 23214
rect 19516 22652 19572 22708
rect 19292 21756 19348 21812
rect 19068 18844 19124 18900
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20188 19852 20244 19908
rect 19628 19628 19684 19684
rect 19516 19122 19572 19124
rect 19516 19070 19518 19122
rect 19518 19070 19570 19122
rect 19570 19070 19572 19122
rect 19516 19068 19572 19070
rect 18844 17612 18900 17668
rect 18732 17106 18788 17108
rect 18732 17054 18734 17106
rect 18734 17054 18786 17106
rect 18786 17054 18788 17106
rect 18732 17052 18788 17054
rect 16156 9266 16212 9268
rect 16156 9214 16158 9266
rect 16158 9214 16210 9266
rect 16210 9214 16212 9266
rect 16156 9212 16212 9214
rect 18396 13356 18452 13412
rect 15820 9154 15876 9156
rect 15820 9102 15822 9154
rect 15822 9102 15874 9154
rect 15874 9102 15876 9154
rect 15820 9100 15876 9102
rect 16716 9154 16772 9156
rect 16716 9102 16718 9154
rect 16718 9102 16770 9154
rect 16770 9102 16772 9154
rect 16716 9100 16772 9102
rect 15820 8652 15876 8708
rect 16268 8370 16324 8372
rect 16268 8318 16270 8370
rect 16270 8318 16322 8370
rect 16322 8318 16324 8370
rect 16268 8316 16324 8318
rect 15932 8092 15988 8148
rect 15820 7698 15876 7700
rect 15820 7646 15822 7698
rect 15822 7646 15874 7698
rect 15874 7646 15876 7698
rect 15820 7644 15876 7646
rect 16604 8316 16660 8372
rect 16716 8652 16772 8708
rect 16604 8146 16660 8148
rect 16604 8094 16606 8146
rect 16606 8094 16658 8146
rect 16658 8094 16660 8146
rect 16604 8092 16660 8094
rect 15148 6690 15204 6692
rect 15148 6638 15150 6690
rect 15150 6638 15202 6690
rect 15202 6638 15204 6690
rect 15148 6636 15204 6638
rect 15596 6412 15652 6468
rect 14700 4114 14756 4116
rect 14700 4062 14702 4114
rect 14702 4062 14754 4114
rect 14754 4062 14756 4114
rect 14700 4060 14756 4062
rect 14028 3500 14084 3556
rect 16828 8092 16884 8148
rect 16940 8034 16996 8036
rect 16940 7982 16942 8034
rect 16942 7982 16994 8034
rect 16994 7982 16996 8034
rect 16940 7980 16996 7982
rect 17164 7532 17220 7588
rect 17388 7868 17444 7924
rect 16828 7474 16884 7476
rect 16828 7422 16830 7474
rect 16830 7422 16882 7474
rect 16882 7422 16884 7474
rect 16828 7420 16884 7422
rect 16604 7308 16660 7364
rect 18508 13074 18564 13076
rect 18508 13022 18510 13074
rect 18510 13022 18562 13074
rect 18562 13022 18564 13074
rect 18508 13020 18564 13022
rect 18732 16828 18788 16884
rect 19292 18226 19348 18228
rect 19292 18174 19294 18226
rect 19294 18174 19346 18226
rect 19346 18174 19348 18226
rect 19292 18172 19348 18174
rect 19068 18060 19124 18116
rect 18844 15708 18900 15764
rect 19068 14028 19124 14084
rect 18732 12684 18788 12740
rect 18620 12402 18676 12404
rect 18620 12350 18622 12402
rect 18622 12350 18674 12402
rect 18674 12350 18676 12402
rect 18620 12348 18676 12350
rect 19180 10108 19236 10164
rect 18508 9884 18564 9940
rect 19404 10610 19460 10612
rect 19404 10558 19406 10610
rect 19406 10558 19458 10610
rect 19458 10558 19460 10610
rect 19404 10556 19460 10558
rect 18508 8540 18564 8596
rect 18732 8316 18788 8372
rect 18508 8258 18564 8260
rect 18508 8206 18510 8258
rect 18510 8206 18562 8258
rect 18562 8206 18564 8258
rect 18508 8204 18564 8206
rect 17836 7756 17892 7812
rect 18620 7980 18676 8036
rect 18172 7644 18228 7700
rect 17724 7586 17780 7588
rect 17724 7534 17726 7586
rect 17726 7534 17778 7586
rect 17778 7534 17780 7586
rect 17724 7532 17780 7534
rect 17948 6802 18004 6804
rect 17948 6750 17950 6802
rect 17950 6750 18002 6802
rect 18002 6750 18004 6802
rect 17948 6748 18004 6750
rect 17836 6636 17892 6692
rect 17052 5628 17108 5684
rect 16380 5122 16436 5124
rect 16380 5070 16382 5122
rect 16382 5070 16434 5122
rect 16434 5070 16436 5122
rect 16380 5068 16436 5070
rect 17500 5068 17556 5124
rect 18396 7644 18452 7700
rect 18284 6748 18340 6804
rect 18396 5682 18452 5684
rect 18396 5630 18398 5682
rect 18398 5630 18450 5682
rect 18450 5630 18452 5682
rect 18396 5628 18452 5630
rect 19180 8540 19236 8596
rect 19068 8428 19124 8484
rect 18956 7644 19012 7700
rect 19292 8316 19348 8372
rect 18956 7308 19012 7364
rect 19292 7756 19348 7812
rect 18844 6636 18900 6692
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16828 19684 16884
rect 20300 19292 20356 19348
rect 20300 18396 20356 18452
rect 20636 25282 20692 25284
rect 20636 25230 20638 25282
rect 20638 25230 20690 25282
rect 20690 25230 20692 25282
rect 20636 25228 20692 25230
rect 20860 25282 20916 25284
rect 20860 25230 20862 25282
rect 20862 25230 20914 25282
rect 20914 25230 20916 25282
rect 20860 25228 20916 25230
rect 20748 22652 20804 22708
rect 20524 19628 20580 19684
rect 20748 19346 20804 19348
rect 20748 19294 20750 19346
rect 20750 19294 20802 19346
rect 20802 19294 20804 19346
rect 20748 19292 20804 19294
rect 20748 19068 20804 19124
rect 21420 27132 21476 27188
rect 21308 27074 21364 27076
rect 21308 27022 21310 27074
rect 21310 27022 21362 27074
rect 21362 27022 21364 27074
rect 21308 27020 21364 27022
rect 21420 25788 21476 25844
rect 21196 25452 21252 25508
rect 21420 25394 21476 25396
rect 21420 25342 21422 25394
rect 21422 25342 21474 25394
rect 21474 25342 21476 25394
rect 21420 25340 21476 25342
rect 21420 22652 21476 22708
rect 20636 18284 20692 18340
rect 20412 17948 20468 18004
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20188 15538 20244 15540
rect 20188 15486 20190 15538
rect 20190 15486 20242 15538
rect 20242 15486 20244 15538
rect 20188 15484 20244 15486
rect 19628 14476 19684 14532
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 20524 14588 20580 14644
rect 20972 16994 21028 16996
rect 20972 16942 20974 16994
rect 20974 16942 21026 16994
rect 21026 16942 21028 16994
rect 20972 16940 21028 16942
rect 20860 15484 20916 15540
rect 21756 29820 21812 29876
rect 21980 34748 22036 34804
rect 22652 36988 22708 37044
rect 22988 36540 23044 36596
rect 23324 36482 23380 36484
rect 23324 36430 23326 36482
rect 23326 36430 23378 36482
rect 23378 36430 23380 36482
rect 23324 36428 23380 36430
rect 23660 36482 23716 36484
rect 23660 36430 23662 36482
rect 23662 36430 23714 36482
rect 23714 36430 23716 36482
rect 23660 36428 23716 36430
rect 22652 36370 22708 36372
rect 22652 36318 22654 36370
rect 22654 36318 22706 36370
rect 22706 36318 22708 36370
rect 22652 36316 22708 36318
rect 22540 36092 22596 36148
rect 22764 35698 22820 35700
rect 22764 35646 22766 35698
rect 22766 35646 22818 35698
rect 22818 35646 22820 35698
rect 22764 35644 22820 35646
rect 22428 35420 22484 35476
rect 22316 35084 22372 35140
rect 23100 35868 23156 35924
rect 22428 34802 22484 34804
rect 22428 34750 22430 34802
rect 22430 34750 22482 34802
rect 22482 34750 22484 34802
rect 22428 34748 22484 34750
rect 22316 34188 22372 34244
rect 22204 32396 22260 32452
rect 22092 31666 22148 31668
rect 22092 31614 22094 31666
rect 22094 31614 22146 31666
rect 22146 31614 22148 31666
rect 22092 31612 22148 31614
rect 22204 30994 22260 30996
rect 22204 30942 22206 30994
rect 22206 30942 22258 30994
rect 22258 30942 22260 30994
rect 22204 30940 22260 30942
rect 21980 30828 22036 30884
rect 22428 30156 22484 30212
rect 22316 30098 22372 30100
rect 22316 30046 22318 30098
rect 22318 30046 22370 30098
rect 22370 30046 22372 30098
rect 22316 30044 22372 30046
rect 22540 30044 22596 30100
rect 21756 27746 21812 27748
rect 21756 27694 21758 27746
rect 21758 27694 21810 27746
rect 21810 27694 21812 27746
rect 21756 27692 21812 27694
rect 21980 27074 22036 27076
rect 21980 27022 21982 27074
rect 21982 27022 22034 27074
rect 22034 27022 22036 27074
rect 21980 27020 22036 27022
rect 22428 29484 22484 29540
rect 22316 27804 22372 27860
rect 22652 27692 22708 27748
rect 24444 36482 24500 36484
rect 24444 36430 24446 36482
rect 24446 36430 24498 36482
rect 24498 36430 24500 36482
rect 24444 36428 24500 36430
rect 24220 36316 24276 36372
rect 23884 36204 23940 36260
rect 24332 35868 24388 35924
rect 24556 35756 24612 35812
rect 23100 34972 23156 35028
rect 23436 35026 23492 35028
rect 23436 34974 23438 35026
rect 23438 34974 23490 35026
rect 23490 34974 23492 35026
rect 23436 34972 23492 34974
rect 24332 35698 24388 35700
rect 24332 35646 24334 35698
rect 24334 35646 24386 35698
rect 24386 35646 24388 35698
rect 24332 35644 24388 35646
rect 24220 35586 24276 35588
rect 24220 35534 24222 35586
rect 24222 35534 24274 35586
rect 24274 35534 24276 35586
rect 24220 35532 24276 35534
rect 24108 35420 24164 35476
rect 24332 35308 24388 35364
rect 23884 34690 23940 34692
rect 23884 34638 23886 34690
rect 23886 34638 23938 34690
rect 23938 34638 23940 34690
rect 23884 34636 23940 34638
rect 24556 34524 24612 34580
rect 23772 34242 23828 34244
rect 23772 34190 23774 34242
rect 23774 34190 23826 34242
rect 23826 34190 23828 34242
rect 23772 34188 23828 34190
rect 23884 33964 23940 34020
rect 24444 34018 24500 34020
rect 24444 33966 24446 34018
rect 24446 33966 24498 34018
rect 24498 33966 24500 34018
rect 24444 33964 24500 33966
rect 25004 36258 25060 36260
rect 25004 36206 25006 36258
rect 25006 36206 25058 36258
rect 25058 36206 25060 36258
rect 25004 36204 25060 36206
rect 24780 34636 24836 34692
rect 24444 33068 24500 33124
rect 23548 31836 23604 31892
rect 23100 31164 23156 31220
rect 22988 30098 23044 30100
rect 22988 30046 22990 30098
rect 22990 30046 23042 30098
rect 23042 30046 23044 30098
rect 22988 30044 23044 30046
rect 23324 27804 23380 27860
rect 21756 26178 21812 26180
rect 21756 26126 21758 26178
rect 21758 26126 21810 26178
rect 21810 26126 21812 26178
rect 21756 26124 21812 26126
rect 22092 23436 22148 23492
rect 21756 23324 21812 23380
rect 22988 27020 23044 27076
rect 22316 26012 22372 26068
rect 22204 22540 22260 22596
rect 22092 20690 22148 20692
rect 22092 20638 22094 20690
rect 22094 20638 22146 20690
rect 22146 20638 22148 20690
rect 22092 20636 22148 20638
rect 21644 20076 21700 20132
rect 21980 19516 22036 19572
rect 21532 19068 21588 19124
rect 21196 18956 21252 19012
rect 21196 18396 21252 18452
rect 21868 18396 21924 18452
rect 22204 19292 22260 19348
rect 22092 19122 22148 19124
rect 22092 19070 22094 19122
rect 22094 19070 22146 19122
rect 22146 19070 22148 19122
rect 22092 19068 22148 19070
rect 21644 17948 21700 18004
rect 22316 19404 22372 19460
rect 22764 26290 22820 26292
rect 22764 26238 22766 26290
rect 22766 26238 22818 26290
rect 22818 26238 22820 26290
rect 22764 26236 22820 26238
rect 22988 26178 23044 26180
rect 22988 26126 22990 26178
rect 22990 26126 23042 26178
rect 23042 26126 23044 26178
rect 22988 26124 23044 26126
rect 22652 25506 22708 25508
rect 22652 25454 22654 25506
rect 22654 25454 22706 25506
rect 22706 25454 22708 25506
rect 22652 25452 22708 25454
rect 24220 31724 24276 31780
rect 24108 31388 24164 31444
rect 23660 31218 23716 31220
rect 23660 31166 23662 31218
rect 23662 31166 23714 31218
rect 23714 31166 23716 31218
rect 23660 31164 23716 31166
rect 23212 25228 23268 25284
rect 23996 28700 24052 28756
rect 23436 25228 23492 25284
rect 23996 25116 24052 25172
rect 22764 22092 22820 22148
rect 22428 19292 22484 19348
rect 22652 20690 22708 20692
rect 22652 20638 22654 20690
rect 22654 20638 22706 20690
rect 22706 20638 22708 20690
rect 22652 20636 22708 20638
rect 22652 19404 22708 19460
rect 22764 19906 22820 19908
rect 22764 19854 22766 19906
rect 22766 19854 22818 19906
rect 22818 19854 22820 19906
rect 22764 19852 22820 19854
rect 22316 18844 22372 18900
rect 22764 18620 22820 18676
rect 23324 24722 23380 24724
rect 23324 24670 23326 24722
rect 23326 24670 23378 24722
rect 23378 24670 23380 24722
rect 23324 24668 23380 24670
rect 22988 23324 23044 23380
rect 23884 25004 23940 25060
rect 23884 24668 23940 24724
rect 23436 23324 23492 23380
rect 23548 24556 23604 24612
rect 23548 23212 23604 23268
rect 23324 20860 23380 20916
rect 23100 20802 23156 20804
rect 23100 20750 23102 20802
rect 23102 20750 23154 20802
rect 23154 20750 23156 20802
rect 23100 20748 23156 20750
rect 24668 32450 24724 32452
rect 24668 32398 24670 32450
rect 24670 32398 24722 32450
rect 24722 32398 24724 32450
rect 24668 32396 24724 32398
rect 26572 39394 26628 39396
rect 26572 39342 26574 39394
rect 26574 39342 26626 39394
rect 26626 39342 26628 39394
rect 26572 39340 26628 39342
rect 28364 41186 28420 41188
rect 28364 41134 28366 41186
rect 28366 41134 28418 41186
rect 28418 41134 28420 41186
rect 28364 41132 28420 41134
rect 27804 39506 27860 39508
rect 27804 39454 27806 39506
rect 27806 39454 27858 39506
rect 27858 39454 27860 39506
rect 27804 39452 27860 39454
rect 26236 38722 26292 38724
rect 26236 38670 26238 38722
rect 26238 38670 26290 38722
rect 26290 38670 26292 38722
rect 26236 38668 26292 38670
rect 25788 36988 25844 37044
rect 25676 36540 25732 36596
rect 25228 35810 25284 35812
rect 25228 35758 25230 35810
rect 25230 35758 25282 35810
rect 25282 35758 25284 35810
rect 25228 35756 25284 35758
rect 25340 35308 25396 35364
rect 25564 35308 25620 35364
rect 25788 35420 25844 35476
rect 26572 36988 26628 37044
rect 26460 36370 26516 36372
rect 26460 36318 26462 36370
rect 26462 36318 26514 36370
rect 26514 36318 26516 36370
rect 26460 36316 26516 36318
rect 25564 34636 25620 34692
rect 25228 33346 25284 33348
rect 25228 33294 25230 33346
rect 25230 33294 25282 33346
rect 25282 33294 25284 33346
rect 25228 33292 25284 33294
rect 24444 31388 24500 31444
rect 24780 31778 24836 31780
rect 24780 31726 24782 31778
rect 24782 31726 24834 31778
rect 24834 31726 24836 31778
rect 24780 31724 24836 31726
rect 25116 31778 25172 31780
rect 25116 31726 25118 31778
rect 25118 31726 25170 31778
rect 25170 31726 25172 31778
rect 25116 31724 25172 31726
rect 25004 31164 25060 31220
rect 24332 30210 24388 30212
rect 24332 30158 24334 30210
rect 24334 30158 24386 30210
rect 24386 30158 24388 30210
rect 24332 30156 24388 30158
rect 24780 27186 24836 27188
rect 24780 27134 24782 27186
rect 24782 27134 24834 27186
rect 24834 27134 24836 27186
rect 24780 27132 24836 27134
rect 25340 29820 25396 29876
rect 25564 28700 25620 28756
rect 25676 27356 25732 27412
rect 25452 27132 25508 27188
rect 25228 27074 25284 27076
rect 25228 27022 25230 27074
rect 25230 27022 25282 27074
rect 25282 27022 25284 27074
rect 25228 27020 25284 27022
rect 24892 24444 24948 24500
rect 24892 21644 24948 21700
rect 24332 21586 24388 21588
rect 24332 21534 24334 21586
rect 24334 21534 24386 21586
rect 24386 21534 24388 21586
rect 24332 21532 24388 21534
rect 24220 21308 24276 21364
rect 23772 20690 23828 20692
rect 23772 20638 23774 20690
rect 23774 20638 23826 20690
rect 23826 20638 23828 20690
rect 23772 20636 23828 20638
rect 22988 20076 23044 20132
rect 23100 20018 23156 20020
rect 23100 19966 23102 20018
rect 23102 19966 23154 20018
rect 23154 19966 23156 20018
rect 23100 19964 23156 19966
rect 23548 20076 23604 20132
rect 23100 19458 23156 19460
rect 23100 19406 23102 19458
rect 23102 19406 23154 19458
rect 23154 19406 23156 19458
rect 23100 19404 23156 19406
rect 22876 19292 22932 19348
rect 23436 19516 23492 19572
rect 21868 17778 21924 17780
rect 21868 17726 21870 17778
rect 21870 17726 21922 17778
rect 21922 17726 21924 17778
rect 21868 17724 21924 17726
rect 22316 17724 22372 17780
rect 22204 17106 22260 17108
rect 22204 17054 22206 17106
rect 22206 17054 22258 17106
rect 22258 17054 22260 17106
rect 22204 17052 22260 17054
rect 21868 16994 21924 16996
rect 21868 16942 21870 16994
rect 21870 16942 21922 16994
rect 21922 16942 21924 16994
rect 21868 16940 21924 16942
rect 22764 16940 22820 16996
rect 22652 16828 22708 16884
rect 23324 18620 23380 18676
rect 21532 15538 21588 15540
rect 21532 15486 21534 15538
rect 21534 15486 21586 15538
rect 21586 15486 21588 15538
rect 21532 15484 21588 15486
rect 20748 13132 20804 13188
rect 20412 12348 20468 12404
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19740 10722 19796 10724
rect 19740 10670 19742 10722
rect 19742 10670 19794 10722
rect 19794 10670 19796 10722
rect 19740 10668 19796 10670
rect 20524 10668 20580 10724
rect 19740 9602 19796 9604
rect 19740 9550 19742 9602
rect 19742 9550 19794 9602
rect 19794 9550 19796 9602
rect 19740 9548 19796 9550
rect 20748 10498 20804 10500
rect 20748 10446 20750 10498
rect 20750 10446 20802 10498
rect 20802 10446 20804 10498
rect 20748 10444 20804 10446
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19516 8428 19572 8484
rect 19516 7980 19572 8036
rect 19852 8316 19908 8372
rect 21196 14530 21252 14532
rect 21196 14478 21198 14530
rect 21198 14478 21250 14530
rect 21250 14478 21252 14530
rect 21196 14476 21252 14478
rect 21644 14476 21700 14532
rect 21308 13132 21364 13188
rect 21868 14140 21924 14196
rect 21756 12236 21812 12292
rect 20972 9660 21028 9716
rect 21196 10892 21252 10948
rect 20636 9602 20692 9604
rect 20636 9550 20638 9602
rect 20638 9550 20690 9602
rect 20690 9550 20692 9602
rect 20636 9548 20692 9550
rect 20748 9436 20804 9492
rect 21868 10610 21924 10612
rect 21868 10558 21870 10610
rect 21870 10558 21922 10610
rect 21922 10558 21924 10610
rect 21868 10556 21924 10558
rect 21644 10444 21700 10500
rect 21196 9436 21252 9492
rect 21420 9714 21476 9716
rect 21420 9662 21422 9714
rect 21422 9662 21474 9714
rect 21474 9662 21476 9714
rect 21420 9660 21476 9662
rect 20860 9324 20916 9380
rect 21308 9324 21364 9380
rect 20748 8652 20804 8708
rect 20524 8316 20580 8372
rect 19964 8204 20020 8260
rect 20188 8258 20244 8260
rect 20188 8206 20190 8258
rect 20190 8206 20242 8258
rect 20242 8206 20244 8258
rect 20188 8204 20244 8206
rect 19964 8034 20020 8036
rect 19964 7982 19966 8034
rect 19966 7982 20018 8034
rect 20018 7982 20020 8034
rect 19964 7980 20020 7982
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20748 8146 20804 8148
rect 20748 8094 20750 8146
rect 20750 8094 20802 8146
rect 20802 8094 20804 8146
rect 20748 8092 20804 8094
rect 20300 7698 20356 7700
rect 20300 7646 20302 7698
rect 20302 7646 20354 7698
rect 20354 7646 20356 7698
rect 20300 7644 20356 7646
rect 19964 7586 20020 7588
rect 19964 7534 19966 7586
rect 19966 7534 20018 7586
rect 20018 7534 20020 7586
rect 19964 7532 20020 7534
rect 20636 7586 20692 7588
rect 20636 7534 20638 7586
rect 20638 7534 20690 7586
rect 20690 7534 20692 7586
rect 20636 7532 20692 7534
rect 19516 7196 19572 7252
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 21196 8988 21252 9044
rect 20972 8652 21028 8708
rect 22092 14140 22148 14196
rect 22092 13746 22148 13748
rect 22092 13694 22094 13746
rect 22094 13694 22146 13746
rect 22146 13694 22148 13746
rect 22092 13692 22148 13694
rect 22652 14812 22708 14868
rect 22540 14530 22596 14532
rect 22540 14478 22542 14530
rect 22542 14478 22594 14530
rect 22594 14478 22596 14530
rect 22540 14476 22596 14478
rect 22540 13858 22596 13860
rect 22540 13806 22542 13858
rect 22542 13806 22594 13858
rect 22594 13806 22596 13858
rect 22540 13804 22596 13806
rect 22652 13692 22708 13748
rect 22876 15538 22932 15540
rect 22876 15486 22878 15538
rect 22878 15486 22930 15538
rect 22930 15486 22932 15538
rect 22876 15484 22932 15486
rect 23884 19852 23940 19908
rect 23772 19404 23828 19460
rect 23884 19234 23940 19236
rect 23884 19182 23886 19234
rect 23886 19182 23938 19234
rect 23938 19182 23940 19234
rect 23884 19180 23940 19182
rect 23772 19122 23828 19124
rect 23772 19070 23774 19122
rect 23774 19070 23826 19122
rect 23826 19070 23828 19122
rect 23772 19068 23828 19070
rect 23548 18508 23604 18564
rect 24556 20802 24612 20804
rect 24556 20750 24558 20802
rect 24558 20750 24610 20802
rect 24610 20750 24612 20802
rect 24556 20748 24612 20750
rect 24556 19628 24612 19684
rect 24108 19516 24164 19572
rect 24332 19346 24388 19348
rect 24332 19294 24334 19346
rect 24334 19294 24386 19346
rect 24386 19294 24388 19346
rect 24332 19292 24388 19294
rect 24780 19234 24836 19236
rect 24780 19182 24782 19234
rect 24782 19182 24834 19234
rect 24834 19182 24836 19234
rect 24780 19180 24836 19182
rect 25564 26796 25620 26852
rect 25228 25228 25284 25284
rect 25788 26514 25844 26516
rect 25788 26462 25790 26514
rect 25790 26462 25842 26514
rect 25842 26462 25844 26514
rect 25788 26460 25844 26462
rect 25564 25340 25620 25396
rect 25452 25004 25508 25060
rect 26348 33964 26404 34020
rect 26124 33122 26180 33124
rect 26124 33070 26126 33122
rect 26126 33070 26178 33122
rect 26178 33070 26180 33122
rect 26124 33068 26180 33070
rect 26236 29426 26292 29428
rect 26236 29374 26238 29426
rect 26238 29374 26290 29426
rect 26290 29374 26292 29426
rect 26236 29372 26292 29374
rect 26908 34860 26964 34916
rect 26908 34354 26964 34356
rect 26908 34302 26910 34354
rect 26910 34302 26962 34354
rect 26962 34302 26964 34354
rect 26908 34300 26964 34302
rect 28364 40348 28420 40404
rect 29372 41410 29428 41412
rect 29372 41358 29374 41410
rect 29374 41358 29426 41410
rect 29426 41358 29428 41410
rect 29372 41356 29428 41358
rect 29596 41356 29652 41412
rect 29708 40796 29764 40852
rect 29260 40626 29316 40628
rect 29260 40574 29262 40626
rect 29262 40574 29314 40626
rect 29314 40574 29316 40626
rect 29260 40572 29316 40574
rect 29484 40012 29540 40068
rect 28476 39788 28532 39844
rect 29372 39842 29428 39844
rect 29372 39790 29374 39842
rect 29374 39790 29426 39842
rect 29426 39790 29428 39842
rect 29372 39788 29428 39790
rect 27916 34300 27972 34356
rect 26572 33346 26628 33348
rect 26572 33294 26574 33346
rect 26574 33294 26626 33346
rect 26626 33294 26628 33346
rect 26572 33292 26628 33294
rect 28700 37938 28756 37940
rect 28700 37886 28702 37938
rect 28702 37886 28754 37938
rect 28754 37886 28756 37938
rect 28700 37884 28756 37886
rect 28700 37436 28756 37492
rect 28588 35868 28644 35924
rect 27692 32844 27748 32900
rect 26684 32396 26740 32452
rect 26460 30156 26516 30212
rect 26572 30044 26628 30100
rect 26796 29820 26852 29876
rect 26572 28812 26628 28868
rect 26012 28642 26068 28644
rect 26012 28590 26014 28642
rect 26014 28590 26066 28642
rect 26066 28590 26068 28642
rect 26012 28588 26068 28590
rect 26348 28588 26404 28644
rect 25900 25004 25956 25060
rect 25900 22204 25956 22260
rect 25452 22092 25508 22148
rect 25340 21644 25396 21700
rect 26012 22146 26068 22148
rect 26012 22094 26014 22146
rect 26014 22094 26066 22146
rect 26066 22094 26068 22146
rect 26012 22092 26068 22094
rect 25676 21532 25732 21588
rect 25676 20524 25732 20580
rect 25564 17778 25620 17780
rect 25564 17726 25566 17778
rect 25566 17726 25618 17778
rect 25618 17726 25620 17778
rect 25564 17724 25620 17726
rect 25116 17500 25172 17556
rect 25564 15260 25620 15316
rect 23324 14812 23380 14868
rect 22092 11116 22148 11172
rect 22876 14252 22932 14308
rect 22092 10892 22148 10948
rect 23212 14140 23268 14196
rect 24220 14588 24276 14644
rect 24220 14028 24276 14084
rect 24108 13244 24164 13300
rect 22204 10834 22260 10836
rect 22204 10782 22206 10834
rect 22206 10782 22258 10834
rect 22258 10782 22260 10834
rect 22204 10780 22260 10782
rect 24108 12348 24164 12404
rect 22316 10668 22372 10724
rect 21980 10220 22036 10276
rect 22652 9996 22708 10052
rect 23100 10610 23156 10612
rect 23100 10558 23102 10610
rect 23102 10558 23154 10610
rect 23154 10558 23156 10610
rect 23100 10556 23156 10558
rect 22988 10498 23044 10500
rect 22988 10446 22990 10498
rect 22990 10446 23042 10498
rect 23042 10446 23044 10498
rect 22988 10444 23044 10446
rect 21868 9714 21924 9716
rect 21868 9662 21870 9714
rect 21870 9662 21922 9714
rect 21922 9662 21924 9714
rect 21868 9660 21924 9662
rect 21420 8876 21476 8932
rect 21980 8652 22036 8708
rect 22316 9436 22372 9492
rect 21644 8316 21700 8372
rect 21420 7698 21476 7700
rect 21420 7646 21422 7698
rect 21422 7646 21474 7698
rect 21474 7646 21476 7698
rect 21420 7644 21476 7646
rect 21756 8258 21812 8260
rect 21756 8206 21758 8258
rect 21758 8206 21810 8258
rect 21810 8206 21812 8258
rect 21756 8204 21812 8206
rect 21868 8092 21924 8148
rect 21756 7698 21812 7700
rect 21756 7646 21758 7698
rect 21758 7646 21810 7698
rect 21810 7646 21812 7698
rect 21756 7644 21812 7646
rect 22428 9100 22484 9156
rect 22764 9714 22820 9716
rect 22764 9662 22766 9714
rect 22766 9662 22818 9714
rect 22818 9662 22820 9714
rect 22764 9660 22820 9662
rect 22652 9212 22708 9268
rect 23996 10834 24052 10836
rect 23996 10782 23998 10834
rect 23998 10782 24050 10834
rect 24050 10782 24052 10834
rect 23996 10780 24052 10782
rect 23212 9772 23268 9828
rect 23324 9996 23380 10052
rect 23100 9436 23156 9492
rect 23996 9714 24052 9716
rect 23996 9662 23998 9714
rect 23998 9662 24050 9714
rect 24050 9662 24052 9714
rect 23996 9660 24052 9662
rect 23996 9266 24052 9268
rect 23996 9214 23998 9266
rect 23998 9214 24050 9266
rect 24050 9214 24052 9266
rect 23996 9212 24052 9214
rect 24220 10780 24276 10836
rect 23436 9100 23492 9156
rect 23100 8930 23156 8932
rect 23100 8878 23102 8930
rect 23102 8878 23154 8930
rect 23154 8878 23156 8930
rect 23100 8876 23156 8878
rect 22988 8764 23044 8820
rect 22316 8316 22372 8372
rect 22540 8316 22596 8372
rect 22204 8092 22260 8148
rect 23548 8370 23604 8372
rect 23548 8318 23550 8370
rect 23550 8318 23602 8370
rect 23602 8318 23604 8370
rect 23548 8316 23604 8318
rect 22876 7980 22932 8036
rect 21308 6636 21364 6692
rect 25340 14924 25396 14980
rect 25452 13244 25508 13300
rect 26012 18450 26068 18452
rect 26012 18398 26014 18450
rect 26014 18398 26066 18450
rect 26066 18398 26068 18450
rect 26012 18396 26068 18398
rect 26348 16044 26404 16100
rect 25900 15820 25956 15876
rect 25788 15148 25844 15204
rect 26908 28754 26964 28756
rect 26908 28702 26910 28754
rect 26910 28702 26962 28754
rect 26962 28702 26964 28754
rect 26908 28700 26964 28702
rect 28476 34636 28532 34692
rect 29260 37884 29316 37940
rect 30716 40460 30772 40516
rect 30044 38834 30100 38836
rect 30044 38782 30046 38834
rect 30046 38782 30098 38834
rect 30098 38782 30100 38834
rect 30044 38780 30100 38782
rect 29148 36988 29204 37044
rect 29148 35868 29204 35924
rect 28700 34524 28756 34580
rect 28812 35308 28868 35364
rect 28588 33404 28644 33460
rect 27804 31948 27860 32004
rect 28252 31948 28308 32004
rect 29596 35586 29652 35588
rect 29596 35534 29598 35586
rect 29598 35534 29650 35586
rect 29650 35534 29652 35586
rect 29596 35532 29652 35534
rect 31164 38834 31220 38836
rect 31164 38782 31166 38834
rect 31166 38782 31218 38834
rect 31218 38782 31220 38834
rect 31164 38780 31220 38782
rect 28924 33740 28980 33796
rect 29372 33740 29428 33796
rect 29260 32844 29316 32900
rect 27244 31836 27300 31892
rect 27692 31500 27748 31556
rect 28140 31500 28196 31556
rect 27916 30210 27972 30212
rect 27916 30158 27918 30210
rect 27918 30158 27970 30210
rect 27970 30158 27972 30210
rect 27916 30156 27972 30158
rect 27356 28700 27412 28756
rect 27244 28642 27300 28644
rect 27244 28590 27246 28642
rect 27246 28590 27298 28642
rect 27298 28590 27300 28642
rect 27244 28588 27300 28590
rect 27692 29820 27748 29876
rect 27692 28812 27748 28868
rect 27580 28588 27636 28644
rect 28700 31836 28756 31892
rect 29260 31836 29316 31892
rect 28700 31612 28756 31668
rect 28140 30044 28196 30100
rect 28252 29820 28308 29876
rect 27804 28530 27860 28532
rect 27804 28478 27806 28530
rect 27806 28478 27858 28530
rect 27858 28478 27860 28530
rect 27804 28476 27860 28478
rect 27356 28140 27412 28196
rect 27132 25730 27188 25732
rect 27132 25678 27134 25730
rect 27134 25678 27186 25730
rect 27186 25678 27188 25730
rect 27132 25676 27188 25678
rect 27020 25394 27076 25396
rect 27020 25342 27022 25394
rect 27022 25342 27074 25394
rect 27074 25342 27076 25394
rect 27020 25340 27076 25342
rect 27020 24556 27076 24612
rect 26684 21586 26740 21588
rect 26684 21534 26686 21586
rect 26686 21534 26738 21586
rect 26738 21534 26740 21586
rect 26684 21532 26740 21534
rect 26684 21308 26740 21364
rect 26908 22370 26964 22372
rect 26908 22318 26910 22370
rect 26910 22318 26962 22370
rect 26962 22318 26964 22370
rect 26908 22316 26964 22318
rect 27132 22204 27188 22260
rect 27132 21980 27188 22036
rect 27020 21868 27076 21924
rect 26796 20748 26852 20804
rect 27916 28252 27972 28308
rect 27916 27244 27972 27300
rect 27692 24610 27748 24612
rect 27692 24558 27694 24610
rect 27694 24558 27746 24610
rect 27746 24558 27748 24610
rect 27692 24556 27748 24558
rect 27356 22428 27412 22484
rect 28028 23042 28084 23044
rect 28028 22990 28030 23042
rect 28030 22990 28082 23042
rect 28082 22990 28084 23042
rect 28028 22988 28084 22990
rect 27804 22428 27860 22484
rect 27692 22316 27748 22372
rect 27356 21698 27412 21700
rect 27356 21646 27358 21698
rect 27358 21646 27410 21698
rect 27410 21646 27412 21698
rect 27356 21644 27412 21646
rect 27244 21420 27300 21476
rect 27132 20802 27188 20804
rect 27132 20750 27134 20802
rect 27134 20750 27186 20802
rect 27186 20750 27188 20802
rect 27132 20748 27188 20750
rect 27020 19180 27076 19236
rect 27468 21308 27524 21364
rect 28812 30156 28868 30212
rect 29260 30156 29316 30212
rect 29036 30044 29092 30100
rect 28588 28252 28644 28308
rect 29260 29596 29316 29652
rect 29036 28588 29092 28644
rect 29148 28364 29204 28420
rect 31164 33906 31220 33908
rect 31164 33854 31166 33906
rect 31166 33854 31218 33906
rect 31218 33854 31220 33906
rect 31164 33852 31220 33854
rect 30380 33740 30436 33796
rect 31500 40236 31556 40292
rect 32956 41916 33012 41972
rect 33180 41410 33236 41412
rect 33180 41358 33182 41410
rect 33182 41358 33234 41410
rect 33234 41358 33236 41410
rect 33180 41356 33236 41358
rect 32172 40348 32228 40404
rect 32396 41132 32452 41188
rect 31836 39788 31892 39844
rect 36988 41916 37044 41972
rect 34076 41020 34132 41076
rect 34076 40626 34132 40628
rect 34076 40574 34078 40626
rect 34078 40574 34130 40626
rect 34130 40574 34132 40626
rect 34076 40572 34132 40574
rect 33068 40012 33124 40068
rect 33404 40348 33460 40404
rect 33068 39842 33124 39844
rect 33068 39790 33070 39842
rect 33070 39790 33122 39842
rect 33122 39790 33124 39842
rect 33068 39788 33124 39790
rect 31836 38668 31892 38724
rect 31500 37826 31556 37828
rect 31500 37774 31502 37826
rect 31502 37774 31554 37826
rect 31554 37774 31556 37826
rect 31500 37772 31556 37774
rect 30156 33458 30212 33460
rect 30156 33406 30158 33458
rect 30158 33406 30210 33458
rect 30210 33406 30212 33458
rect 30156 33404 30212 33406
rect 31724 36204 31780 36260
rect 31724 34300 31780 34356
rect 29932 31666 29988 31668
rect 29932 31614 29934 31666
rect 29934 31614 29986 31666
rect 29986 31614 29988 31666
rect 29932 31612 29988 31614
rect 29932 30098 29988 30100
rect 29932 30046 29934 30098
rect 29934 30046 29986 30098
rect 29986 30046 29988 30098
rect 29932 30044 29988 30046
rect 30268 30210 30324 30212
rect 30268 30158 30270 30210
rect 30270 30158 30322 30210
rect 30322 30158 30324 30210
rect 30268 30156 30324 30158
rect 29708 29036 29764 29092
rect 28588 27074 28644 27076
rect 28588 27022 28590 27074
rect 28590 27022 28642 27074
rect 28642 27022 28644 27074
rect 28588 27020 28644 27022
rect 28812 27244 28868 27300
rect 29372 27298 29428 27300
rect 29372 27246 29374 27298
rect 29374 27246 29426 27298
rect 29426 27246 29428 27298
rect 29372 27244 29428 27246
rect 29148 25676 29204 25732
rect 29260 27020 29316 27076
rect 29820 28700 29876 28756
rect 30268 28700 30324 28756
rect 30044 28364 30100 28420
rect 30268 28418 30324 28420
rect 30268 28366 30270 28418
rect 30270 28366 30322 28418
rect 30322 28366 30324 28418
rect 30268 28364 30324 28366
rect 30716 29036 30772 29092
rect 30716 28530 30772 28532
rect 30716 28478 30718 28530
rect 30718 28478 30770 28530
rect 30770 28478 30772 28530
rect 30716 28476 30772 28478
rect 30716 27916 30772 27972
rect 30828 27804 30884 27860
rect 30828 27074 30884 27076
rect 30828 27022 30830 27074
rect 30830 27022 30882 27074
rect 30882 27022 30884 27074
rect 30828 27020 30884 27022
rect 28476 25004 28532 25060
rect 28924 25004 28980 25060
rect 28140 21980 28196 22036
rect 28700 24668 28756 24724
rect 29372 24892 29428 24948
rect 28028 21868 28084 21924
rect 27692 20972 27748 21028
rect 28140 21532 28196 21588
rect 28028 21362 28084 21364
rect 28028 21310 28030 21362
rect 28030 21310 28082 21362
rect 28082 21310 28084 21362
rect 28028 21308 28084 21310
rect 27244 19292 27300 19348
rect 26908 16492 26964 16548
rect 26572 15260 26628 15316
rect 27020 15260 27076 15316
rect 26348 14924 26404 14980
rect 25676 14476 25732 14532
rect 26124 14306 26180 14308
rect 26124 14254 26126 14306
rect 26126 14254 26178 14306
rect 26178 14254 26180 14306
rect 26124 14252 26180 14254
rect 25676 13916 25732 13972
rect 26012 13858 26068 13860
rect 26012 13806 26014 13858
rect 26014 13806 26066 13858
rect 26066 13806 26068 13858
rect 26012 13804 26068 13806
rect 26348 14028 26404 14084
rect 26460 13858 26516 13860
rect 26460 13806 26462 13858
rect 26462 13806 26514 13858
rect 26514 13806 26516 13858
rect 26460 13804 26516 13806
rect 26236 13356 26292 13412
rect 26684 12908 26740 12964
rect 26348 12402 26404 12404
rect 26348 12350 26350 12402
rect 26350 12350 26402 12402
rect 26402 12350 26404 12402
rect 26348 12348 26404 12350
rect 26908 14418 26964 14420
rect 26908 14366 26910 14418
rect 26910 14366 26962 14418
rect 26962 14366 26964 14418
rect 26908 14364 26964 14366
rect 27132 14140 27188 14196
rect 27356 17106 27412 17108
rect 27356 17054 27358 17106
rect 27358 17054 27410 17106
rect 27410 17054 27412 17106
rect 27356 17052 27412 17054
rect 27580 15820 27636 15876
rect 27356 15314 27412 15316
rect 27356 15262 27358 15314
rect 27358 15262 27410 15314
rect 27410 15262 27412 15314
rect 27356 15260 27412 15262
rect 27468 15148 27524 15204
rect 27356 14418 27412 14420
rect 27356 14366 27358 14418
rect 27358 14366 27410 14418
rect 27410 14366 27412 14418
rect 27356 14364 27412 14366
rect 28028 20130 28084 20132
rect 28028 20078 28030 20130
rect 28030 20078 28082 20130
rect 28082 20078 28084 20130
rect 28028 20076 28084 20078
rect 27804 18508 27860 18564
rect 27916 16716 27972 16772
rect 28140 19180 28196 19236
rect 28028 16044 28084 16100
rect 28140 17052 28196 17108
rect 28140 15820 28196 15876
rect 27804 15202 27860 15204
rect 27804 15150 27806 15202
rect 27806 15150 27858 15202
rect 27858 15150 27860 15202
rect 27804 15148 27860 15150
rect 27692 14588 27748 14644
rect 29372 24050 29428 24052
rect 29372 23998 29374 24050
rect 29374 23998 29426 24050
rect 29426 23998 29428 24050
rect 29372 23996 29428 23998
rect 29708 23996 29764 24052
rect 29484 23772 29540 23828
rect 30156 24780 30212 24836
rect 29596 23436 29652 23492
rect 29036 23154 29092 23156
rect 29036 23102 29038 23154
rect 29038 23102 29090 23154
rect 29090 23102 29092 23154
rect 29036 23100 29092 23102
rect 29372 23100 29428 23156
rect 29484 22876 29540 22932
rect 28364 21868 28420 21924
rect 28476 22092 28532 22148
rect 28364 20972 28420 21028
rect 28588 21756 28644 21812
rect 28812 21586 28868 21588
rect 28812 21534 28814 21586
rect 28814 21534 28866 21586
rect 28866 21534 28868 21586
rect 28812 21532 28868 21534
rect 28588 20860 28644 20916
rect 28812 20972 28868 21028
rect 28476 19740 28532 19796
rect 28588 19346 28644 19348
rect 28588 19294 28590 19346
rect 28590 19294 28642 19346
rect 28642 19294 28644 19346
rect 28588 19292 28644 19294
rect 28588 17778 28644 17780
rect 28588 17726 28590 17778
rect 28590 17726 28642 17778
rect 28642 17726 28644 17778
rect 28588 17724 28644 17726
rect 28812 17052 28868 17108
rect 28700 16828 28756 16884
rect 29148 21868 29204 21924
rect 29372 22428 29428 22484
rect 29820 23154 29876 23156
rect 29820 23102 29822 23154
rect 29822 23102 29874 23154
rect 29874 23102 29876 23154
rect 29820 23100 29876 23102
rect 29708 22988 29764 23044
rect 30156 23772 30212 23828
rect 30044 23324 30100 23380
rect 30156 23154 30212 23156
rect 30156 23102 30158 23154
rect 30158 23102 30210 23154
rect 30210 23102 30212 23154
rect 30156 23100 30212 23102
rect 29596 22092 29652 22148
rect 29372 21868 29428 21924
rect 29932 21868 29988 21924
rect 29260 20802 29316 20804
rect 29260 20750 29262 20802
rect 29262 20750 29314 20802
rect 29314 20750 29316 20802
rect 29260 20748 29316 20750
rect 29036 20130 29092 20132
rect 29036 20078 29038 20130
rect 29038 20078 29090 20130
rect 29090 20078 29092 20130
rect 29036 20076 29092 20078
rect 29596 20690 29652 20692
rect 29596 20638 29598 20690
rect 29598 20638 29650 20690
rect 29650 20638 29652 20690
rect 29596 20636 29652 20638
rect 30044 20636 30100 20692
rect 29372 19906 29428 19908
rect 29372 19854 29374 19906
rect 29374 19854 29426 19906
rect 29426 19854 29428 19906
rect 29372 19852 29428 19854
rect 29260 19740 29316 19796
rect 29484 19740 29540 19796
rect 29148 19292 29204 19348
rect 29260 17106 29316 17108
rect 29260 17054 29262 17106
rect 29262 17054 29314 17106
rect 29314 17054 29316 17106
rect 29260 17052 29316 17054
rect 29148 16882 29204 16884
rect 29148 16830 29150 16882
rect 29150 16830 29202 16882
rect 29202 16830 29204 16882
rect 29148 16828 29204 16830
rect 28924 16716 28980 16772
rect 28476 16156 28532 16212
rect 29148 15986 29204 15988
rect 29148 15934 29150 15986
rect 29150 15934 29202 15986
rect 29202 15934 29204 15986
rect 29148 15932 29204 15934
rect 29708 15484 29764 15540
rect 27020 13746 27076 13748
rect 27020 13694 27022 13746
rect 27022 13694 27074 13746
rect 27074 13694 27076 13746
rect 27020 13692 27076 13694
rect 27244 12962 27300 12964
rect 27244 12910 27246 12962
rect 27246 12910 27298 12962
rect 27298 12910 27300 12962
rect 27244 12908 27300 12910
rect 27132 12348 27188 12404
rect 27244 11676 27300 11732
rect 25116 9884 25172 9940
rect 25340 9996 25396 10052
rect 24332 9548 24388 9604
rect 27244 9996 27300 10052
rect 26012 8930 26068 8932
rect 26012 8878 26014 8930
rect 26014 8878 26066 8930
rect 26066 8878 26068 8930
rect 26012 8876 26068 8878
rect 27804 14140 27860 14196
rect 27468 13356 27524 13412
rect 28140 14306 28196 14308
rect 28140 14254 28142 14306
rect 28142 14254 28194 14306
rect 28194 14254 28196 14306
rect 28140 14252 28196 14254
rect 28700 14700 28756 14756
rect 29260 14306 29316 14308
rect 29260 14254 29262 14306
rect 29262 14254 29314 14306
rect 29314 14254 29316 14306
rect 29260 14252 29316 14254
rect 28252 14028 28308 14084
rect 28140 12796 28196 12852
rect 31500 31500 31556 31556
rect 31948 37772 32004 37828
rect 32396 37884 32452 37940
rect 31948 34524 32004 34580
rect 31948 33964 32004 34020
rect 31500 31052 31556 31108
rect 32284 31106 32340 31108
rect 32284 31054 32286 31106
rect 32286 31054 32338 31106
rect 32338 31054 32340 31106
rect 32284 31052 32340 31054
rect 31948 30098 32004 30100
rect 31948 30046 31950 30098
rect 31950 30046 32002 30098
rect 32002 30046 32004 30098
rect 31948 30044 32004 30046
rect 31836 28588 31892 28644
rect 31500 27916 31556 27972
rect 31388 26460 31444 26516
rect 31724 26124 31780 26180
rect 31612 25564 31668 25620
rect 31724 23436 31780 23492
rect 30380 23212 30436 23268
rect 30380 22316 30436 22372
rect 30716 22988 30772 23044
rect 32172 25618 32228 25620
rect 32172 25566 32174 25618
rect 32174 25566 32226 25618
rect 32226 25566 32228 25618
rect 32172 25564 32228 25566
rect 32508 34354 32564 34356
rect 32508 34302 32510 34354
rect 32510 34302 32562 34354
rect 32562 34302 32564 34354
rect 32508 34300 32564 34302
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35980 41186 36036 41188
rect 35980 41134 35982 41186
rect 35982 41134 36034 41186
rect 36034 41134 36036 41186
rect 35980 41132 36036 41134
rect 36316 41132 36372 41188
rect 35980 40402 36036 40404
rect 35980 40350 35982 40402
rect 35982 40350 36034 40402
rect 36034 40350 36036 40402
rect 35980 40348 36036 40350
rect 35644 40236 35700 40292
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35308 39564 35364 39620
rect 35196 39004 35252 39060
rect 34972 38668 35028 38724
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 33180 34018 33236 34020
rect 33180 33966 33182 34018
rect 33182 33966 33234 34018
rect 33234 33966 33236 34018
rect 33180 33964 33236 33966
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 37436 41356 37492 41412
rect 36988 41020 37044 41076
rect 36428 39788 36484 39844
rect 37996 39842 38052 39844
rect 37996 39790 37998 39842
rect 37998 39790 38050 39842
rect 38050 39790 38052 39842
rect 37996 39788 38052 39790
rect 38556 39788 38612 39844
rect 36988 39618 37044 39620
rect 36988 39566 36990 39618
rect 36990 39566 37042 39618
rect 37042 39566 37044 39618
rect 36988 39564 37044 39566
rect 37324 39564 37380 39620
rect 36428 39058 36484 39060
rect 36428 39006 36430 39058
rect 36430 39006 36482 39058
rect 36482 39006 36484 39058
rect 36428 39004 36484 39006
rect 33068 31724 33124 31780
rect 32732 29932 32788 29988
rect 32732 28700 32788 28756
rect 32844 28642 32900 28644
rect 32844 28590 32846 28642
rect 32846 28590 32898 28642
rect 32898 28590 32900 28642
rect 32844 28588 32900 28590
rect 33068 27858 33124 27860
rect 33068 27806 33070 27858
rect 33070 27806 33122 27858
rect 33122 27806 33124 27858
rect 33068 27804 33124 27806
rect 33292 26908 33348 26964
rect 32396 25452 32452 25508
rect 34972 31500 35028 31556
rect 34076 30156 34132 30212
rect 34076 29596 34132 29652
rect 34636 30156 34692 30212
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 33740 28754 33796 28756
rect 33740 28702 33742 28754
rect 33742 28702 33794 28754
rect 33794 28702 33796 28754
rect 33740 28700 33796 28702
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34076 28588 34132 28644
rect 33852 28364 33908 28420
rect 34412 27916 34468 27972
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34748 27298 34804 27300
rect 34748 27246 34750 27298
rect 34750 27246 34802 27298
rect 34802 27246 34804 27298
rect 34748 27244 34804 27246
rect 38332 39340 38388 39396
rect 39116 38946 39172 38948
rect 39116 38894 39118 38946
rect 39118 38894 39170 38946
rect 39170 38894 39172 38946
rect 39116 38892 39172 38894
rect 38892 37996 38948 38052
rect 40796 41410 40852 41412
rect 40796 41358 40798 41410
rect 40798 41358 40850 41410
rect 40850 41358 40852 41410
rect 40796 41356 40852 41358
rect 39788 41186 39844 41188
rect 39788 41134 39790 41186
rect 39790 41134 39842 41186
rect 39842 41134 39844 41186
rect 39788 41132 39844 41134
rect 40908 39842 40964 39844
rect 40908 39790 40910 39842
rect 40910 39790 40962 39842
rect 40962 39790 40964 39842
rect 40908 39788 40964 39790
rect 39900 39618 39956 39620
rect 39900 39566 39902 39618
rect 39902 39566 39954 39618
rect 39954 39566 39956 39618
rect 39900 39564 39956 39566
rect 39676 38220 39732 38276
rect 40908 38274 40964 38276
rect 40908 38222 40910 38274
rect 40910 38222 40962 38274
rect 40962 38222 40964 38274
rect 40908 38220 40964 38222
rect 39900 38050 39956 38052
rect 39900 37998 39902 38050
rect 39902 37998 39954 38050
rect 39954 37998 39956 38050
rect 39900 37996 39956 37998
rect 39452 37660 39508 37716
rect 40572 37660 40628 37716
rect 42812 40962 42868 40964
rect 42812 40910 42814 40962
rect 42814 40910 42866 40962
rect 42866 40910 42868 40962
rect 42812 40908 42868 40910
rect 43148 40402 43204 40404
rect 43148 40350 43150 40402
rect 43150 40350 43202 40402
rect 43202 40350 43204 40402
rect 43148 40348 43204 40350
rect 42812 33852 42868 33908
rect 39452 33404 39508 33460
rect 37772 32956 37828 33012
rect 36988 31554 37044 31556
rect 36988 31502 36990 31554
rect 36990 31502 37042 31554
rect 37042 31502 37044 31554
rect 36988 31500 37044 31502
rect 35868 27244 35924 27300
rect 34412 27132 34468 27188
rect 35196 27186 35252 27188
rect 35196 27134 35198 27186
rect 35198 27134 35250 27186
rect 35250 27134 35252 27186
rect 35196 27132 35252 27134
rect 35980 27132 36036 27188
rect 33964 26796 34020 26852
rect 33852 26178 33908 26180
rect 33852 26126 33854 26178
rect 33854 26126 33906 26178
rect 33906 26126 33908 26178
rect 33852 26124 33908 26126
rect 34412 26124 34468 26180
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 33404 24108 33460 24164
rect 32844 23772 32900 23828
rect 30604 22930 30660 22932
rect 30604 22878 30606 22930
rect 30606 22878 30658 22930
rect 30658 22878 30660 22930
rect 30604 22876 30660 22878
rect 30380 22146 30436 22148
rect 30380 22094 30382 22146
rect 30382 22094 30434 22146
rect 30434 22094 30436 22146
rect 30380 22092 30436 22094
rect 30268 20972 30324 21028
rect 30380 20860 30436 20916
rect 30268 20802 30324 20804
rect 30268 20750 30270 20802
rect 30270 20750 30322 20802
rect 30322 20750 30324 20802
rect 30268 20748 30324 20750
rect 30380 20242 30436 20244
rect 30380 20190 30382 20242
rect 30382 20190 30434 20242
rect 30434 20190 30436 20242
rect 30380 20188 30436 20190
rect 30268 17052 30324 17108
rect 29708 14700 29764 14756
rect 30380 15148 30436 15204
rect 29372 13692 29428 13748
rect 29820 14252 29876 14308
rect 30156 13804 30212 13860
rect 28476 11676 28532 11732
rect 28140 9714 28196 9716
rect 28140 9662 28142 9714
rect 28142 9662 28194 9714
rect 28194 9662 28196 9714
rect 28140 9660 28196 9662
rect 26124 8316 26180 8372
rect 24220 5180 24276 5236
rect 23884 4562 23940 4564
rect 23884 4510 23886 4562
rect 23886 4510 23938 4562
rect 23938 4510 23940 4562
rect 23884 4508 23940 4510
rect 22988 4338 23044 4340
rect 22988 4286 22990 4338
rect 22990 4286 23042 4338
rect 23042 4286 23044 4338
rect 22988 4284 23044 4286
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 27804 3612 27860 3668
rect 29372 11676 29428 11732
rect 30156 10834 30212 10836
rect 30156 10782 30158 10834
rect 30158 10782 30210 10834
rect 30210 10782 30212 10834
rect 30156 10780 30212 10782
rect 29148 10444 29204 10500
rect 29708 9884 29764 9940
rect 29260 9826 29316 9828
rect 29260 9774 29262 9826
rect 29262 9774 29314 9826
rect 29314 9774 29316 9826
rect 29260 9772 29316 9774
rect 29596 9548 29652 9604
rect 29596 8988 29652 9044
rect 28812 4338 28868 4340
rect 28812 4286 28814 4338
rect 28814 4286 28866 4338
rect 28866 4286 28868 4338
rect 28812 4284 28868 4286
rect 30268 9602 30324 9604
rect 30268 9550 30270 9602
rect 30270 9550 30322 9602
rect 30322 9550 30324 9602
rect 30268 9548 30324 9550
rect 30940 22316 30996 22372
rect 30716 20860 30772 20916
rect 30940 20914 30996 20916
rect 30940 20862 30942 20914
rect 30942 20862 30994 20914
rect 30994 20862 30996 20914
rect 30940 20860 30996 20862
rect 31276 21196 31332 21252
rect 31836 21196 31892 21252
rect 30828 18508 30884 18564
rect 30828 17724 30884 17780
rect 31612 20860 31668 20916
rect 31724 20018 31780 20020
rect 31724 19966 31726 20018
rect 31726 19966 31778 20018
rect 31778 19966 31780 20018
rect 31724 19964 31780 19966
rect 31500 19852 31556 19908
rect 31612 18508 31668 18564
rect 32508 20018 32564 20020
rect 32508 19966 32510 20018
rect 32510 19966 32562 20018
rect 32562 19966 32564 20018
rect 32508 19964 32564 19966
rect 32508 19180 32564 19236
rect 32396 19068 32452 19124
rect 33292 23548 33348 23604
rect 33068 23324 33124 23380
rect 33852 23660 33908 23716
rect 34076 23548 34132 23604
rect 33628 23212 33684 23268
rect 33852 23436 33908 23492
rect 32060 18396 32116 18452
rect 31500 17724 31556 17780
rect 33180 18396 33236 18452
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34860 23660 34916 23716
rect 33852 22370 33908 22372
rect 33852 22318 33854 22370
rect 33854 22318 33906 22370
rect 33906 22318 33908 22370
rect 33852 22316 33908 22318
rect 34076 22540 34132 22596
rect 33628 21868 33684 21924
rect 34972 22988 35028 23044
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35420 22370 35476 22372
rect 35420 22318 35422 22370
rect 35422 22318 35474 22370
rect 35474 22318 35476 22370
rect 35420 22316 35476 22318
rect 36652 23042 36708 23044
rect 36652 22990 36654 23042
rect 36654 22990 36706 23042
rect 36706 22990 36708 23042
rect 36652 22988 36708 22990
rect 36204 22316 36260 22372
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 33852 20188 33908 20244
rect 34188 20076 34244 20132
rect 35644 20860 35700 20916
rect 34972 19964 35028 20020
rect 35084 20300 35140 20356
rect 35420 20076 35476 20132
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34860 19404 34916 19460
rect 34972 19292 35028 19348
rect 33292 18956 33348 19012
rect 33068 18284 33124 18340
rect 33740 19068 33796 19124
rect 34748 18956 34804 19012
rect 35084 19180 35140 19236
rect 34188 18396 34244 18452
rect 34972 18450 35028 18452
rect 34972 18398 34974 18450
rect 34974 18398 35026 18450
rect 35026 18398 35028 18450
rect 34972 18396 35028 18398
rect 33292 17106 33348 17108
rect 33292 17054 33294 17106
rect 33294 17054 33346 17106
rect 33346 17054 33348 17106
rect 33292 17052 33348 17054
rect 35644 19180 35700 19236
rect 36204 19404 36260 19460
rect 36428 19346 36484 19348
rect 36428 19294 36430 19346
rect 36430 19294 36482 19346
rect 36482 19294 36484 19346
rect 36428 19292 36484 19294
rect 35420 18450 35476 18452
rect 35420 18398 35422 18450
rect 35422 18398 35474 18450
rect 35474 18398 35476 18450
rect 35420 18396 35476 18398
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 32396 15538 32452 15540
rect 32396 15486 32398 15538
rect 32398 15486 32450 15538
rect 32450 15486 32452 15538
rect 32396 15484 32452 15486
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 33404 13468 33460 13524
rect 32732 13020 32788 13076
rect 30604 9884 30660 9940
rect 31388 9548 31444 9604
rect 30380 4284 30436 4340
rect 29596 4060 29652 4116
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
rect 30828 4114 30884 4116
rect 30828 4062 30830 4114
rect 30830 4062 30882 4114
rect 30882 4062 30884 4114
rect 30828 4060 30884 4062
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35084 7532 35140 7588
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35084 4284 35140 4340
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34972 3612 35028 3668
rect 37100 19234 37156 19236
rect 37100 19182 37102 19234
rect 37102 19182 37154 19234
rect 37154 19182 37156 19234
rect 37100 19180 37156 19182
rect 38220 19964 38276 20020
rect 38332 18674 38388 18676
rect 38332 18622 38334 18674
rect 38334 18622 38386 18674
rect 38386 18622 38388 18674
rect 38332 18620 38388 18622
rect 37772 6636 37828 6692
rect 39340 18508 39396 18564
rect 36764 4060 36820 4116
rect 37996 4114 38052 4116
rect 37996 4062 37998 4114
rect 37998 4062 38050 4114
rect 38050 4062 38052 4114
rect 37996 4060 38052 4062
rect 36988 3666 37044 3668
rect 36988 3614 36990 3666
rect 36990 3614 37042 3666
rect 37042 3614 37044 3666
rect 36988 3612 37044 3614
rect 38556 3612 38612 3668
rect 41132 32844 41188 32900
rect 42588 31388 42644 31444
rect 43148 31388 43204 31444
rect 41132 23324 41188 23380
rect 42812 23378 42868 23380
rect 42812 23326 42814 23378
rect 42814 23326 42866 23378
rect 42866 23326 42868 23378
rect 42812 23324 42868 23326
rect 43148 22428 43204 22484
rect 39452 13916 39508 13972
rect 40348 20524 40404 20580
rect 42812 13970 42868 13972
rect 42812 13918 42814 13970
rect 42814 13918 42866 13970
rect 42866 13918 42868 13970
rect 42812 13916 42868 13918
rect 42588 13468 42644 13524
rect 43148 13468 43204 13524
rect 42812 6636 42868 6692
rect 42588 5122 42644 5124
rect 42588 5070 42590 5122
rect 42590 5070 42642 5122
rect 42642 5070 42644 5122
rect 42588 5068 42644 5070
rect 43148 5122 43204 5124
rect 43148 5070 43150 5122
rect 43150 5070 43202 5122
rect 43202 5070 43204 5122
rect 43148 5068 43204 5070
rect 43148 4508 43204 4564
rect 42812 4284 42868 4340
rect 40796 3666 40852 3668
rect 40796 3614 40798 3666
rect 40798 3614 40850 3666
rect 40850 3614 40852 3666
rect 40796 3612 40852 3614
<< metal3 >>
rect 0 41972 800 42000
rect 0 41916 5404 41972
rect 5460 41916 5470 41972
rect 32946 41916 32956 41972
rect 33012 41916 36988 41972
rect 37044 41916 37054 41972
rect 0 41888 800 41916
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 23986 41356 23996 41412
rect 24052 41356 25564 41412
rect 25620 41356 25630 41412
rect 26226 41356 26236 41412
rect 26292 41356 29372 41412
rect 29428 41356 29438 41412
rect 29586 41356 29596 41412
rect 29652 41356 33180 41412
rect 33236 41356 33246 41412
rect 37426 41356 37436 41412
rect 37492 41356 40796 41412
rect 40852 41356 40862 41412
rect 4722 41244 4732 41300
rect 4788 41244 5628 41300
rect 5684 41244 5694 41300
rect 11218 41244 11228 41300
rect 11284 41244 12124 41300
rect 12180 41244 12190 41300
rect 22754 41132 22764 41188
rect 22820 41132 24556 41188
rect 24612 41132 24622 41188
rect 27458 41132 27468 41188
rect 27524 41132 28364 41188
rect 28420 41132 28430 41188
rect 32386 41132 32396 41188
rect 32452 41132 35980 41188
rect 36036 41132 36046 41188
rect 36306 41132 36316 41188
rect 36372 41132 39788 41188
rect 39844 41132 39854 41188
rect 4274 41020 4284 41076
rect 4340 41020 11452 41076
rect 11508 41020 11518 41076
rect 34066 41020 34076 41076
rect 34132 41020 36988 41076
rect 37044 41020 37054 41076
rect 4386 40908 4396 40964
rect 4452 40908 7644 40964
rect 7700 40908 7710 40964
rect 31892 40908 42812 40964
rect 42868 40908 42878 40964
rect 31892 40852 31948 40908
rect 29698 40796 29708 40852
rect 29764 40796 31948 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 4162 40684 4172 40740
rect 4228 40684 7868 40740
rect 7924 40684 7934 40740
rect 8194 40684 8204 40740
rect 8260 40684 11900 40740
rect 11956 40684 11966 40740
rect 0 40628 800 40656
rect 0 40572 1932 40628
rect 1988 40572 1998 40628
rect 8306 40572 8316 40628
rect 8372 40572 9660 40628
rect 9716 40572 9726 40628
rect 25106 40572 25116 40628
rect 25172 40572 26348 40628
rect 26404 40572 26414 40628
rect 27346 40572 27356 40628
rect 27412 40572 29260 40628
rect 29316 40572 29326 40628
rect 31892 40572 34076 40628
rect 34132 40572 34142 40628
rect 0 40544 800 40572
rect 31892 40516 31948 40572
rect 8372 40460 11676 40516
rect 11732 40460 11742 40516
rect 24658 40460 24668 40516
rect 24724 40460 25340 40516
rect 25396 40460 25406 40516
rect 30706 40460 30716 40516
rect 30772 40460 31948 40516
rect 8372 40404 8428 40460
rect 44200 40404 45000 40432
rect 4946 40348 4956 40404
rect 5012 40348 5964 40404
rect 6020 40348 6030 40404
rect 7186 40348 7196 40404
rect 7252 40348 8428 40404
rect 10546 40348 10556 40404
rect 10612 40348 11452 40404
rect 11508 40348 12348 40404
rect 12404 40348 12414 40404
rect 19618 40348 19628 40404
rect 19684 40348 20748 40404
rect 20804 40348 20814 40404
rect 28354 40348 28364 40404
rect 28420 40348 32172 40404
rect 32228 40348 32238 40404
rect 33394 40348 33404 40404
rect 33460 40348 35980 40404
rect 36036 40348 36046 40404
rect 43138 40348 43148 40404
rect 43204 40348 45000 40404
rect 44200 40320 45000 40348
rect 31490 40236 31500 40292
rect 31556 40236 35644 40292
rect 35700 40236 35710 40292
rect 29474 40012 29484 40068
rect 29540 40012 33068 40068
rect 33124 40012 33134 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 15586 39788 15596 39844
rect 15652 39788 20188 39844
rect 22866 39788 22876 39844
rect 22932 39788 24108 39844
rect 24164 39788 24174 39844
rect 28466 39788 28476 39844
rect 28532 39788 29372 39844
rect 29428 39788 29438 39844
rect 31826 39788 31836 39844
rect 31892 39788 33068 39844
rect 33124 39788 33134 39844
rect 36418 39788 36428 39844
rect 36484 39788 37996 39844
rect 38052 39788 38062 39844
rect 38546 39788 38556 39844
rect 38612 39788 40908 39844
rect 40964 39788 40974 39844
rect 20132 39732 20188 39788
rect 3826 39676 3836 39732
rect 3892 39676 7196 39732
rect 7252 39676 8204 39732
rect 8260 39676 8270 39732
rect 12226 39676 12236 39732
rect 12292 39676 13468 39732
rect 13524 39676 16156 39732
rect 16212 39676 16222 39732
rect 20132 39676 26236 39732
rect 26292 39676 26302 39732
rect 924 39564 1932 39620
rect 1988 39564 1998 39620
rect 21634 39564 21644 39620
rect 21700 39564 23100 39620
rect 23156 39564 23166 39620
rect 35298 39564 35308 39620
rect 35364 39564 36988 39620
rect 37044 39564 37054 39620
rect 37314 39564 37324 39620
rect 37380 39564 39900 39620
rect 39956 39564 39966 39620
rect 0 39284 800 39312
rect 924 39284 980 39564
rect 16818 39452 16828 39508
rect 16884 39452 22428 39508
rect 22484 39452 22494 39508
rect 25778 39452 25788 39508
rect 25844 39452 27804 39508
rect 27860 39452 27870 39508
rect 6402 39340 6412 39396
rect 6468 39340 7644 39396
rect 7700 39340 8652 39396
rect 8708 39340 12012 39396
rect 12068 39340 12908 39396
rect 12964 39340 14924 39396
rect 14980 39340 15372 39396
rect 15428 39340 16268 39396
rect 16324 39340 16940 39396
rect 16996 39340 17388 39396
rect 17444 39340 17724 39396
rect 17780 39340 17790 39396
rect 18162 39340 18172 39396
rect 18228 39340 23884 39396
rect 23940 39340 25228 39396
rect 25284 39340 25294 39396
rect 26562 39340 26572 39396
rect 26628 39340 38332 39396
rect 38388 39340 38398 39396
rect 0 39228 980 39284
rect 0 39200 800 39228
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 24658 39116 24668 39172
rect 24724 39116 31948 39172
rect 16370 39004 16380 39060
rect 16436 39004 24332 39060
rect 24388 39004 24398 39060
rect 31892 38948 31948 39116
rect 35186 39004 35196 39060
rect 35252 39004 36428 39060
rect 36484 39004 36494 39060
rect 4274 38892 4284 38948
rect 4340 38892 7980 38948
rect 8036 38892 8046 38948
rect 16146 38892 16156 38948
rect 16212 38892 16492 38948
rect 16548 38892 16558 38948
rect 31892 38892 39116 38948
rect 39172 38892 39182 38948
rect 1922 38780 1932 38836
rect 1988 38780 5180 38836
rect 5236 38780 5740 38836
rect 5796 38780 6412 38836
rect 6468 38780 6478 38836
rect 7186 38780 7196 38836
rect 7252 38780 9436 38836
rect 9492 38780 9502 38836
rect 14802 38780 14812 38836
rect 14868 38780 15484 38836
rect 15540 38780 18620 38836
rect 18676 38780 19068 38836
rect 19124 38780 19134 38836
rect 30034 38780 30044 38836
rect 30100 38780 31164 38836
rect 31220 38780 31230 38836
rect 1362 38668 1372 38724
rect 1428 38668 8764 38724
rect 8820 38668 8830 38724
rect 19506 38668 19516 38724
rect 19572 38668 21868 38724
rect 21924 38668 21934 38724
rect 24098 38668 24108 38724
rect 24164 38668 25116 38724
rect 25172 38668 26236 38724
rect 26292 38668 26302 38724
rect 31826 38668 31836 38724
rect 31892 38668 34972 38724
rect 35028 38668 35038 38724
rect 4722 38556 4732 38612
rect 4788 38556 8148 38612
rect 8092 38500 8148 38556
rect 8082 38444 8092 38500
rect 8148 38444 8158 38500
rect 12562 38444 12572 38500
rect 12628 38444 14140 38500
rect 14196 38444 14206 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 16258 38332 16268 38388
rect 16324 38332 17164 38388
rect 17220 38332 17230 38388
rect 15810 38220 15820 38276
rect 15876 38220 20188 38276
rect 20244 38220 20254 38276
rect 39666 38220 39676 38276
rect 39732 38220 40908 38276
rect 40964 38220 40974 38276
rect 1922 38108 1932 38164
rect 1988 38108 1998 38164
rect 11330 38108 11340 38164
rect 11396 38108 11788 38164
rect 11844 38108 11854 38164
rect 15092 38108 16380 38164
rect 16436 38108 17276 38164
rect 17332 38108 17342 38164
rect 17490 38108 17500 38164
rect 17556 38108 20748 38164
rect 20804 38108 24668 38164
rect 24724 38108 24734 38164
rect 0 37940 800 37968
rect 1932 37940 1988 38108
rect 15092 38052 15148 38108
rect 4834 37996 4844 38052
rect 4900 37996 5740 38052
rect 5796 37996 5806 38052
rect 14018 37996 14028 38052
rect 14084 37996 15148 38052
rect 15474 37996 15484 38052
rect 15540 37996 15550 38052
rect 38882 37996 38892 38052
rect 38948 37996 39900 38052
rect 39956 37996 39966 38052
rect 0 37884 1988 37940
rect 7970 37884 7980 37940
rect 8036 37884 8204 37940
rect 8260 37884 8270 37940
rect 9762 37884 9772 37940
rect 9828 37884 10556 37940
rect 10612 37884 10622 37940
rect 0 37856 800 37884
rect 15484 37828 15540 37996
rect 17602 37884 17612 37940
rect 17668 37884 18060 37940
rect 18116 37884 18126 37940
rect 28690 37884 28700 37940
rect 28756 37884 29260 37940
rect 29316 37884 32396 37940
rect 32452 37884 32462 37940
rect 4050 37772 4060 37828
rect 4116 37772 7756 37828
rect 7812 37772 7822 37828
rect 12114 37772 12124 37828
rect 12180 37772 13916 37828
rect 13972 37772 15540 37828
rect 16930 37772 16940 37828
rect 16996 37772 17388 37828
rect 17444 37772 17454 37828
rect 31490 37772 31500 37828
rect 31556 37772 31948 37828
rect 32004 37772 32014 37828
rect 7522 37660 7532 37716
rect 7588 37660 7980 37716
rect 8036 37660 8046 37716
rect 12898 37660 12908 37716
rect 12964 37660 14140 37716
rect 14196 37660 15260 37716
rect 15316 37660 15326 37716
rect 39442 37660 39452 37716
rect 39508 37660 40572 37716
rect 40628 37660 40638 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 6626 37548 6636 37604
rect 6692 37548 15148 37604
rect 15204 37548 16268 37604
rect 16324 37548 16334 37604
rect 5842 37436 5852 37492
rect 5908 37436 7532 37492
rect 7588 37436 7598 37492
rect 14354 37436 14364 37492
rect 14420 37436 15932 37492
rect 15988 37436 28700 37492
rect 28756 37436 28766 37492
rect 4274 37324 4284 37380
rect 4340 37324 6748 37380
rect 6804 37324 6814 37380
rect 18050 37324 18060 37380
rect 18116 37324 19516 37380
rect 19572 37324 20076 37380
rect 20132 37324 20142 37380
rect 4946 37212 4956 37268
rect 5012 37212 6972 37268
rect 7028 37212 7038 37268
rect 7186 37212 7196 37268
rect 7252 37212 11564 37268
rect 11620 37212 12348 37268
rect 12404 37212 12414 37268
rect 17714 37212 17724 37268
rect 17780 37212 18396 37268
rect 18452 37212 18462 37268
rect 9874 37100 9884 37156
rect 9940 37100 10556 37156
rect 10612 37100 10622 37156
rect 11106 37100 11116 37156
rect 11172 37100 22428 37156
rect 22484 37100 22494 37156
rect 8418 36988 8428 37044
rect 8484 36988 11060 37044
rect 15362 36988 15372 37044
rect 15428 36988 17500 37044
rect 17556 36988 17566 37044
rect 22642 36988 22652 37044
rect 22708 36988 25788 37044
rect 25844 36988 25854 37044
rect 26562 36988 26572 37044
rect 26628 36988 29148 37044
rect 29204 36988 29214 37044
rect 11004 36932 11060 36988
rect 5058 36876 5068 36932
rect 5124 36876 7308 36932
rect 7364 36876 7756 36932
rect 7812 36876 8316 36932
rect 8372 36876 8382 36932
rect 8530 36876 8540 36932
rect 8596 36876 9324 36932
rect 9380 36876 9390 36932
rect 10994 36876 11004 36932
rect 11060 36876 11070 36932
rect 15474 36876 15484 36932
rect 15540 36876 17948 36932
rect 18004 36876 18014 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 7970 36764 7980 36820
rect 8036 36764 8092 36820
rect 8148 36764 8158 36820
rect 8418 36764 8428 36820
rect 8484 36764 8988 36820
rect 9044 36764 9054 36820
rect 6626 36652 6636 36708
rect 6692 36652 8092 36708
rect 8148 36652 11228 36708
rect 11284 36652 11294 36708
rect 14690 36652 14700 36708
rect 14756 36652 15372 36708
rect 15428 36652 15438 36708
rect 0 36596 800 36624
rect 0 36540 1932 36596
rect 1988 36540 1998 36596
rect 2930 36540 2940 36596
rect 2996 36540 5852 36596
rect 5908 36540 5918 36596
rect 13906 36540 13916 36596
rect 13972 36540 14924 36596
rect 14980 36540 21924 36596
rect 22978 36540 22988 36596
rect 23044 36540 25676 36596
rect 25732 36540 25742 36596
rect 0 36512 800 36540
rect 5954 36428 5964 36484
rect 6020 36428 6524 36484
rect 6580 36428 6590 36484
rect 8082 36428 8092 36484
rect 8148 36428 8428 36484
rect 8484 36428 8494 36484
rect 8754 36428 8764 36484
rect 8820 36428 9436 36484
rect 9492 36428 10444 36484
rect 10500 36428 10510 36484
rect 15810 36428 15820 36484
rect 15876 36428 16828 36484
rect 16884 36428 21196 36484
rect 21252 36428 21262 36484
rect 6738 36316 6748 36372
rect 6804 36316 6972 36372
rect 7028 36316 7038 36372
rect 8166 36316 8204 36372
rect 8260 36316 8270 36372
rect 13906 36316 13916 36372
rect 13972 36316 16940 36372
rect 16996 36316 17006 36372
rect 17938 36316 17948 36372
rect 18004 36316 18172 36372
rect 18228 36316 18238 36372
rect 19058 36316 19068 36372
rect 19124 36316 20300 36372
rect 20356 36316 20366 36372
rect 9538 36204 9548 36260
rect 9604 36204 10220 36260
rect 10276 36204 10286 36260
rect 15092 36204 15372 36260
rect 15428 36204 16044 36260
rect 16100 36204 16110 36260
rect 6850 36092 6860 36148
rect 6916 36092 8764 36148
rect 8820 36092 8830 36148
rect 6860 35924 6916 36092
rect 15092 36036 15148 36204
rect 16940 36148 16996 36316
rect 21868 36260 21924 36540
rect 22082 36428 22092 36484
rect 22148 36428 23324 36484
rect 23380 36428 23390 36484
rect 23650 36428 23660 36484
rect 23716 36428 24444 36484
rect 24500 36428 24510 36484
rect 22194 36316 22204 36372
rect 22260 36316 22652 36372
rect 22708 36316 22718 36372
rect 24210 36316 24220 36372
rect 24276 36316 26460 36372
rect 26516 36316 26526 36372
rect 18274 36204 18284 36260
rect 18340 36204 18956 36260
rect 19012 36204 19022 36260
rect 19628 36204 20636 36260
rect 20692 36204 20702 36260
rect 21868 36204 23884 36260
rect 23940 36204 25004 36260
rect 25060 36204 31724 36260
rect 31780 36204 31790 36260
rect 19628 36148 19684 36204
rect 16940 36092 19628 36148
rect 19684 36092 19694 36148
rect 21522 36092 21532 36148
rect 21588 36092 22540 36148
rect 22596 36092 22606 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 7074 35980 7084 36036
rect 7140 35980 15148 36036
rect 23100 35980 26908 36036
rect 23100 35924 23156 35980
rect 26852 35924 26908 35980
rect 5058 35868 5068 35924
rect 5124 35868 6636 35924
rect 6692 35868 6702 35924
rect 6860 35868 7196 35924
rect 7252 35868 7262 35924
rect 7718 35868 7756 35924
rect 7812 35868 7822 35924
rect 23090 35868 23100 35924
rect 23156 35868 23166 35924
rect 24322 35868 24332 35924
rect 24388 35868 24398 35924
rect 26852 35868 28588 35924
rect 28644 35868 29148 35924
rect 29204 35868 29214 35924
rect 24332 35812 24388 35868
rect 13010 35756 13020 35812
rect 13076 35756 13468 35812
rect 13524 35756 13534 35812
rect 20850 35756 20860 35812
rect 20916 35756 21980 35812
rect 22036 35756 22046 35812
rect 22428 35756 24388 35812
rect 24546 35756 24556 35812
rect 24612 35756 25228 35812
rect 25284 35756 25294 35812
rect 12114 35644 12124 35700
rect 12180 35644 12796 35700
rect 12852 35644 12862 35700
rect 14354 35644 14364 35700
rect 14420 35644 15260 35700
rect 15316 35644 19068 35700
rect 19124 35644 19134 35700
rect 1586 35532 1596 35588
rect 1652 35532 6748 35588
rect 6804 35532 6814 35588
rect 7970 35532 7980 35588
rect 8036 35532 8540 35588
rect 8596 35532 8606 35588
rect 9538 35532 9548 35588
rect 9604 35532 13020 35588
rect 13076 35532 13086 35588
rect 8540 35476 8596 35532
rect 22428 35476 22484 35756
rect 22754 35644 22764 35700
rect 22820 35644 24332 35700
rect 24388 35644 24398 35700
rect 24210 35532 24220 35588
rect 24276 35532 29596 35588
rect 29652 35532 29662 35588
rect 5954 35420 5964 35476
rect 6020 35420 7084 35476
rect 7140 35420 7150 35476
rect 8540 35420 20860 35476
rect 20916 35420 20926 35476
rect 22418 35420 22428 35476
rect 22484 35420 22494 35476
rect 24098 35420 24108 35476
rect 24164 35420 25788 35476
rect 25844 35420 25854 35476
rect 11330 35308 11340 35364
rect 11396 35308 12572 35364
rect 12628 35308 12638 35364
rect 24322 35308 24332 35364
rect 24388 35308 25340 35364
rect 25396 35308 25406 35364
rect 25554 35308 25564 35364
rect 25620 35308 28812 35364
rect 28868 35308 28878 35364
rect 0 35252 800 35280
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 0 35196 2044 35252
rect 2100 35196 2110 35252
rect 7634 35196 7644 35252
rect 7700 35196 8204 35252
rect 8260 35196 9772 35252
rect 9828 35196 9838 35252
rect 10322 35196 10332 35252
rect 10388 35196 21980 35252
rect 22036 35196 22046 35252
rect 0 35168 800 35196
rect 6290 35084 6300 35140
rect 6356 35084 10108 35140
rect 10164 35084 10174 35140
rect 11554 35084 11564 35140
rect 11620 35084 13580 35140
rect 13636 35084 20356 35140
rect 20514 35084 20524 35140
rect 20580 35084 21868 35140
rect 21924 35084 22316 35140
rect 22372 35084 22382 35140
rect 20300 35028 20356 35084
rect 1474 34972 1484 35028
rect 1540 34972 18732 35028
rect 18788 34972 18798 35028
rect 20300 34972 23100 35028
rect 23156 34972 23436 35028
rect 23492 34972 23502 35028
rect 4946 34860 4956 34916
rect 5012 34860 5516 34916
rect 5572 34860 5582 34916
rect 10434 34860 10444 34916
rect 10500 34860 11340 34916
rect 11396 34860 11406 34916
rect 16930 34860 16940 34916
rect 16996 34860 26908 34916
rect 26964 34860 26974 34916
rect 2034 34748 2044 34804
rect 2100 34748 4060 34804
rect 4116 34748 7084 34804
rect 7140 34748 7150 34804
rect 15474 34748 15484 34804
rect 15540 34748 15708 34804
rect 15764 34748 16268 34804
rect 16324 34748 17612 34804
rect 17668 34748 17678 34804
rect 17938 34748 17948 34804
rect 18004 34748 20188 34804
rect 20244 34748 20254 34804
rect 21970 34748 21980 34804
rect 22036 34748 22428 34804
rect 22484 34748 22494 34804
rect 23884 34748 26908 34804
rect 23884 34692 23940 34748
rect 26852 34692 26908 34748
rect 12002 34636 12012 34692
rect 12068 34636 12796 34692
rect 12852 34636 12862 34692
rect 13346 34636 13356 34692
rect 13412 34636 15372 34692
rect 15428 34636 15820 34692
rect 15876 34636 15886 34692
rect 19628 34636 23884 34692
rect 23940 34636 23950 34692
rect 24770 34636 24780 34692
rect 24836 34636 25564 34692
rect 25620 34636 25630 34692
rect 26852 34636 28476 34692
rect 28532 34636 28542 34692
rect 19628 34580 19684 34636
rect 15250 34524 15260 34580
rect 15316 34524 19684 34580
rect 20402 34524 20412 34580
rect 20468 34524 21756 34580
rect 21812 34524 24556 34580
rect 24612 34524 24622 34580
rect 28690 34524 28700 34580
rect 28756 34524 31948 34580
rect 32004 34524 32014 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 15026 34412 15036 34468
rect 15092 34412 15708 34468
rect 15764 34412 15774 34468
rect 18722 34300 18732 34356
rect 18788 34300 20300 34356
rect 20356 34300 20366 34356
rect 26898 34300 26908 34356
rect 26964 34300 27916 34356
rect 27972 34300 27982 34356
rect 31714 34300 31724 34356
rect 31780 34300 32508 34356
rect 32564 34300 32574 34356
rect 22306 34188 22316 34244
rect 22372 34188 23772 34244
rect 23828 34188 23838 34244
rect 2146 34076 2156 34132
rect 2212 34076 2604 34132
rect 2660 34076 2670 34132
rect 6412 34076 6748 34132
rect 6804 34076 6814 34132
rect 12786 34076 12796 34132
rect 12852 34076 16380 34132
rect 16436 34076 16446 34132
rect 0 33908 800 33936
rect 0 33852 1932 33908
rect 1988 33852 1998 33908
rect 2258 33852 2268 33908
rect 2324 33852 4620 33908
rect 4676 33852 4686 33908
rect 0 33824 800 33852
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 6412 33572 6468 34076
rect 6626 33964 6636 34020
rect 6692 33964 7308 34020
rect 7364 33964 13356 34020
rect 13412 33964 13422 34020
rect 19170 33964 19180 34020
rect 19236 33964 19516 34020
rect 19572 33964 19582 34020
rect 23874 33964 23884 34020
rect 23940 33964 24444 34020
rect 24500 33964 26348 34020
rect 26404 33964 26414 34020
rect 31938 33964 31948 34020
rect 32004 33964 33180 34020
rect 33236 33964 33246 34020
rect 6738 33852 6748 33908
rect 6804 33852 7532 33908
rect 7588 33852 7598 33908
rect 7746 33852 7756 33908
rect 7812 33852 8092 33908
rect 8148 33852 8158 33908
rect 31154 33852 31164 33908
rect 31220 33852 42812 33908
rect 42868 33852 42878 33908
rect 7756 33796 7812 33852
rect 6962 33740 6972 33796
rect 7028 33740 7812 33796
rect 10882 33740 10892 33796
rect 10948 33740 11340 33796
rect 11396 33740 11406 33796
rect 12898 33740 12908 33796
rect 12964 33740 28924 33796
rect 28980 33740 29372 33796
rect 29428 33740 30380 33796
rect 30436 33740 30446 33796
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 7634 33628 7644 33684
rect 7700 33628 14588 33684
rect 14644 33628 14654 33684
rect 15698 33628 15708 33684
rect 15764 33628 17388 33684
rect 17444 33628 17454 33684
rect 4274 33516 4284 33572
rect 4340 33516 5292 33572
rect 5348 33516 5358 33572
rect 6066 33516 6076 33572
rect 6132 33516 6468 33572
rect 11890 33516 11900 33572
rect 11956 33516 12348 33572
rect 12404 33516 15596 33572
rect 15652 33516 15662 33572
rect 16818 33516 16828 33572
rect 16884 33516 16894 33572
rect 16828 33460 16884 33516
rect 2034 33404 2044 33460
rect 2100 33404 2492 33460
rect 2548 33404 3388 33460
rect 14690 33404 14700 33460
rect 14756 33404 16884 33460
rect 28578 33404 28588 33460
rect 28644 33404 30156 33460
rect 30212 33404 39452 33460
rect 39508 33404 39518 33460
rect 3332 33348 3388 33404
rect 3332 33292 4620 33348
rect 4676 33292 4686 33348
rect 9660 33292 10892 33348
rect 10948 33292 10958 33348
rect 16482 33292 16492 33348
rect 16548 33292 18844 33348
rect 18900 33292 18910 33348
rect 25218 33292 25228 33348
rect 25284 33292 26572 33348
rect 26628 33292 26908 33348
rect 4274 33180 4284 33236
rect 4340 33180 7756 33236
rect 7812 33180 7822 33236
rect 9660 33124 9716 33292
rect 10770 33180 10780 33236
rect 10836 33180 16940 33236
rect 16996 33180 17500 33236
rect 17556 33180 17566 33236
rect 19058 33180 19068 33236
rect 19124 33180 21532 33236
rect 21588 33180 21598 33236
rect 7074 33068 7084 33124
rect 7140 33068 9660 33124
rect 9716 33068 9726 33124
rect 9986 33068 9996 33124
rect 10052 33068 10668 33124
rect 10724 33068 12124 33124
rect 12180 33068 12572 33124
rect 12628 33068 12638 33124
rect 24434 33068 24444 33124
rect 24500 33068 26124 33124
rect 26180 33068 26190 33124
rect 26852 33012 26908 33292
rect 3042 32956 3052 33012
rect 3108 32956 5068 33012
rect 5124 32956 5134 33012
rect 5394 32956 5404 33012
rect 5460 32956 7308 33012
rect 7364 32956 7374 33012
rect 8082 32956 8092 33012
rect 8148 32956 10332 33012
rect 10388 32956 10398 33012
rect 15586 32956 15596 33012
rect 15652 32956 17052 33012
rect 17108 32956 17118 33012
rect 26852 32956 37772 33012
rect 37828 32956 37838 33012
rect 8092 32900 8148 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 3602 32844 3612 32900
rect 3668 32844 4732 32900
rect 4788 32844 8148 32900
rect 10210 32844 10220 32900
rect 10276 32844 10556 32900
rect 10612 32844 17444 32900
rect 27682 32844 27692 32900
rect 27748 32844 29260 32900
rect 29316 32844 41132 32900
rect 41188 32844 41198 32900
rect 7410 32732 7420 32788
rect 7476 32732 8652 32788
rect 8708 32732 8718 32788
rect 4162 32620 4172 32676
rect 4228 32620 6188 32676
rect 6244 32620 6254 32676
rect 13570 32620 13580 32676
rect 13636 32620 14364 32676
rect 14420 32620 14430 32676
rect 0 32564 800 32592
rect 17388 32564 17444 32844
rect 0 32508 1932 32564
rect 1988 32508 1998 32564
rect 7634 32508 7644 32564
rect 7700 32508 9884 32564
rect 9940 32508 9950 32564
rect 14914 32508 14924 32564
rect 14980 32508 16940 32564
rect 16996 32508 17006 32564
rect 17378 32508 17388 32564
rect 17444 32508 18060 32564
rect 18116 32508 18620 32564
rect 18676 32508 18686 32564
rect 0 32480 800 32508
rect 7746 32396 7756 32452
rect 7812 32396 14028 32452
rect 14084 32396 14094 32452
rect 16706 32396 16716 32452
rect 16772 32396 22204 32452
rect 22260 32396 22270 32452
rect 24658 32396 24668 32452
rect 24724 32396 26684 32452
rect 26740 32396 26750 32452
rect 11218 32284 11228 32340
rect 11284 32284 11900 32340
rect 11956 32284 12572 32340
rect 12628 32284 12638 32340
rect 8754 32172 8764 32228
rect 8820 32172 20300 32228
rect 20356 32172 20366 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 11442 32060 11452 32116
rect 11508 32060 12236 32116
rect 12292 32060 12302 32116
rect 6066 31948 6076 32004
rect 6132 31948 6748 32004
rect 6804 31948 6814 32004
rect 8866 31948 8876 32004
rect 8932 31948 10220 32004
rect 10276 31948 10286 32004
rect 11666 31948 11676 32004
rect 11732 31948 13132 32004
rect 13188 31948 13916 32004
rect 13972 31948 13982 32004
rect 27794 31948 27804 32004
rect 27860 31948 28252 32004
rect 28308 31948 28318 32004
rect 7074 31836 7084 31892
rect 7140 31836 8092 31892
rect 8148 31836 10556 31892
rect 10612 31836 10622 31892
rect 19618 31836 19628 31892
rect 19684 31836 21308 31892
rect 21364 31836 23548 31892
rect 23604 31836 27244 31892
rect 27300 31836 28700 31892
rect 28756 31836 29260 31892
rect 29316 31836 29326 31892
rect 9762 31724 9772 31780
rect 9828 31724 14140 31780
rect 14196 31724 14206 31780
rect 14466 31724 14476 31780
rect 14532 31724 15372 31780
rect 15428 31724 15708 31780
rect 15764 31724 15774 31780
rect 20290 31724 20300 31780
rect 20356 31724 24220 31780
rect 24276 31724 24780 31780
rect 24836 31724 24846 31780
rect 25106 31724 25116 31780
rect 25172 31724 33068 31780
rect 33124 31724 33134 31780
rect 8054 31612 8092 31668
rect 8148 31612 8158 31668
rect 9986 31612 9996 31668
rect 10052 31612 11340 31668
rect 11396 31612 20804 31668
rect 20962 31612 20972 31668
rect 21028 31612 22092 31668
rect 22148 31612 22158 31668
rect 28690 31612 28700 31668
rect 28756 31612 29932 31668
rect 29988 31612 29998 31668
rect 20748 31556 20804 31612
rect 7634 31500 7644 31556
rect 7700 31500 8540 31556
rect 8596 31500 9660 31556
rect 9716 31500 9726 31556
rect 10210 31500 10220 31556
rect 10276 31500 11452 31556
rect 11508 31500 11518 31556
rect 14018 31500 14028 31556
rect 14084 31500 14924 31556
rect 14980 31500 16156 31556
rect 16212 31500 16222 31556
rect 17042 31500 17052 31556
rect 17108 31500 20692 31556
rect 20748 31500 27692 31556
rect 27748 31500 28140 31556
rect 28196 31500 31500 31556
rect 31556 31500 31566 31556
rect 34962 31500 34972 31556
rect 35028 31500 36988 31556
rect 37044 31500 37054 31556
rect 20636 31444 20692 31500
rect 44200 31444 45000 31472
rect 2594 31388 2604 31444
rect 2660 31388 5516 31444
rect 5572 31388 8316 31444
rect 8372 31388 8382 31444
rect 11554 31388 11564 31444
rect 11620 31388 12460 31444
rect 12516 31388 15708 31444
rect 15764 31388 16492 31444
rect 16548 31388 16558 31444
rect 20636 31388 24108 31444
rect 24164 31388 24444 31444
rect 24500 31388 24510 31444
rect 42578 31388 42588 31444
rect 42644 31388 43148 31444
rect 43204 31388 45000 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 44200 31360 45000 31388
rect 9202 31276 9212 31332
rect 9268 31276 10892 31332
rect 10948 31276 11676 31332
rect 11732 31276 11742 31332
rect 0 31220 800 31248
rect 0 31164 1932 31220
rect 1988 31164 1998 31220
rect 8306 31164 8316 31220
rect 8372 31164 12908 31220
rect 12964 31164 13804 31220
rect 13860 31164 13870 31220
rect 23090 31164 23100 31220
rect 23156 31164 23660 31220
rect 23716 31164 25004 31220
rect 25060 31164 25070 31220
rect 0 31136 800 31164
rect 8194 31052 8204 31108
rect 8260 31052 10108 31108
rect 10164 31052 10174 31108
rect 12124 31052 14476 31108
rect 14532 31052 14542 31108
rect 17266 31052 17276 31108
rect 17332 31052 19292 31108
rect 19348 31052 19358 31108
rect 31490 31052 31500 31108
rect 31556 31052 32284 31108
rect 32340 31052 32350 31108
rect 12124 30996 12180 31052
rect 7410 30940 7420 30996
rect 7476 30940 12180 30996
rect 12338 30940 12348 30996
rect 12404 30940 14140 30996
rect 14196 30940 14206 30996
rect 20850 30940 20860 30996
rect 20916 30940 22204 30996
rect 22260 30940 22270 30996
rect 15362 30828 15372 30884
rect 15428 30828 16156 30884
rect 16212 30828 16222 30884
rect 21298 30828 21308 30884
rect 21364 30828 21980 30884
rect 22036 30828 22046 30884
rect 12002 30716 12012 30772
rect 12068 30716 16268 30772
rect 16324 30716 16334 30772
rect 10966 30604 11004 30660
rect 11060 30604 11070 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 10322 30492 10332 30548
rect 10388 30492 11228 30548
rect 11284 30492 11294 30548
rect 7858 30380 7868 30436
rect 7924 30380 11788 30436
rect 11844 30380 15932 30436
rect 15988 30380 15998 30436
rect 20066 30380 20076 30436
rect 20132 30380 20972 30436
rect 21028 30380 21038 30436
rect 1922 30268 1932 30324
rect 1988 30268 2604 30324
rect 2660 30268 2670 30324
rect 8082 30268 8092 30324
rect 8148 30268 11676 30324
rect 11732 30268 11742 30324
rect 16146 30268 16156 30324
rect 16212 30268 17724 30324
rect 17780 30268 17790 30324
rect 3714 30156 3724 30212
rect 3780 30156 5740 30212
rect 5796 30156 5806 30212
rect 10098 30156 10108 30212
rect 10164 30156 11452 30212
rect 11508 30156 11518 30212
rect 12002 30156 12012 30212
rect 12068 30156 12572 30212
rect 12628 30156 15820 30212
rect 15876 30156 16940 30212
rect 16996 30156 17006 30212
rect 22418 30156 22428 30212
rect 22484 30156 24332 30212
rect 24388 30156 24398 30212
rect 24556 30156 26460 30212
rect 26516 30156 26526 30212
rect 27906 30156 27916 30212
rect 27972 30156 28812 30212
rect 28868 30156 28878 30212
rect 29250 30156 29260 30212
rect 29316 30156 30268 30212
rect 30324 30156 30334 30212
rect 34066 30156 34076 30212
rect 34132 30156 34636 30212
rect 34692 30156 34702 30212
rect 24556 30100 24612 30156
rect 1250 30044 1260 30100
rect 1316 30044 11116 30100
rect 11172 30044 11182 30100
rect 11442 30044 11452 30100
rect 11508 30044 15988 30100
rect 20738 30044 20748 30100
rect 20804 30044 22316 30100
rect 22372 30044 22382 30100
rect 22530 30044 22540 30100
rect 22596 30044 22988 30100
rect 23044 30044 24612 30100
rect 26562 30044 26572 30100
rect 26628 30044 28140 30100
rect 28196 30044 29036 30100
rect 29092 30044 29102 30100
rect 29922 30044 29932 30100
rect 29988 30044 31948 30100
rect 32004 30044 32014 30100
rect 15932 29988 15988 30044
rect 10098 29932 10108 29988
rect 10164 29932 11676 29988
rect 11732 29932 11742 29988
rect 15932 29932 16268 29988
rect 16324 29932 17052 29988
rect 17108 29932 17118 29988
rect 18050 29932 18060 29988
rect 18116 29932 18396 29988
rect 18452 29932 32732 29988
rect 32788 29932 32798 29988
rect 0 29876 800 29904
rect 0 29820 1820 29876
rect 1876 29820 1886 29876
rect 11442 29820 11452 29876
rect 11508 29820 17612 29876
rect 17668 29820 17678 29876
rect 21746 29820 21756 29876
rect 21812 29820 25340 29876
rect 25396 29820 26796 29876
rect 26852 29820 26862 29876
rect 27682 29820 27692 29876
rect 27748 29820 28252 29876
rect 28308 29820 28318 29876
rect 0 29792 800 29820
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 6738 29708 6748 29764
rect 6804 29708 16156 29764
rect 16212 29708 16222 29764
rect 17378 29708 17388 29764
rect 17444 29708 19684 29764
rect 20626 29708 20636 29764
rect 20692 29708 21196 29764
rect 21252 29708 21262 29764
rect 19628 29652 19684 29708
rect 1474 29596 1484 29652
rect 1540 29596 2044 29652
rect 2100 29596 2110 29652
rect 2706 29596 2716 29652
rect 2772 29596 3276 29652
rect 3332 29596 4172 29652
rect 4228 29596 4844 29652
rect 4900 29596 4910 29652
rect 6962 29596 6972 29652
rect 7028 29596 7868 29652
rect 7924 29596 7934 29652
rect 13906 29596 13916 29652
rect 13972 29596 17500 29652
rect 17556 29596 17566 29652
rect 19628 29596 29260 29652
rect 29316 29596 34076 29652
rect 34132 29596 34142 29652
rect 17042 29484 17052 29540
rect 17108 29484 17836 29540
rect 17892 29484 17902 29540
rect 18050 29484 18060 29540
rect 18116 29484 19068 29540
rect 19124 29484 22428 29540
rect 22484 29484 22494 29540
rect 3826 29372 3836 29428
rect 3892 29372 5068 29428
rect 5124 29372 5134 29428
rect 15138 29372 15148 29428
rect 15204 29372 16604 29428
rect 16660 29372 16670 29428
rect 16930 29372 16940 29428
rect 16996 29372 20412 29428
rect 20468 29372 26236 29428
rect 26292 29372 26302 29428
rect 4386 29260 4396 29316
rect 4452 29260 6076 29316
rect 6132 29260 6142 29316
rect 17602 29260 17612 29316
rect 17668 29260 18508 29316
rect 18564 29260 18574 29316
rect 6626 29148 6636 29204
rect 6692 29148 17948 29204
rect 18004 29148 18014 29204
rect 18498 29036 18508 29092
rect 18564 29036 18956 29092
rect 19012 29036 19628 29092
rect 19684 29036 19694 29092
rect 29698 29036 29708 29092
rect 29764 29036 30716 29092
rect 30772 29036 30782 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 11302 28812 11340 28868
rect 11396 28812 11406 28868
rect 26562 28812 26572 28868
rect 26628 28812 27692 28868
rect 27748 28812 27758 28868
rect 4946 28700 4956 28756
rect 5012 28700 6636 28756
rect 6692 28700 9100 28756
rect 9156 28700 11788 28756
rect 11844 28700 12796 28756
rect 12852 28700 12862 28756
rect 16370 28700 16380 28756
rect 16436 28700 20188 28756
rect 20244 28700 20254 28756
rect 23986 28700 23996 28756
rect 24052 28700 25564 28756
rect 25620 28700 26908 28756
rect 26964 28700 26974 28756
rect 27318 28700 27356 28756
rect 27412 28700 29820 28756
rect 29876 28700 30268 28756
rect 30324 28700 30334 28756
rect 32722 28700 32732 28756
rect 32788 28700 33740 28756
rect 33796 28700 33806 28756
rect 4274 28588 4284 28644
rect 4340 28588 6300 28644
rect 6356 28588 10332 28644
rect 10388 28588 10398 28644
rect 11890 28588 11900 28644
rect 11956 28588 13468 28644
rect 13524 28588 13534 28644
rect 15782 28588 15820 28644
rect 15876 28588 15886 28644
rect 16604 28588 17388 28644
rect 17444 28588 17454 28644
rect 18274 28588 18284 28644
rect 18340 28588 20636 28644
rect 20692 28588 26012 28644
rect 26068 28588 26078 28644
rect 26338 28588 26348 28644
rect 26404 28588 27244 28644
rect 27300 28588 27580 28644
rect 27636 28588 27646 28644
rect 29026 28588 29036 28644
rect 29092 28588 29102 28644
rect 31826 28588 31836 28644
rect 31892 28588 32844 28644
rect 32900 28588 34076 28644
rect 34132 28588 34142 28644
rect 0 28532 800 28560
rect 0 28476 1932 28532
rect 1988 28476 1998 28532
rect 11330 28476 11340 28532
rect 11396 28476 12236 28532
rect 12292 28476 12908 28532
rect 12964 28476 12974 28532
rect 16230 28476 16268 28532
rect 16324 28476 16334 28532
rect 0 28448 800 28476
rect 16604 28420 16660 28588
rect 27580 28420 27636 28588
rect 29036 28532 29092 28588
rect 27794 28476 27804 28532
rect 27860 28476 30716 28532
rect 30772 28476 30782 28532
rect 8418 28364 8428 28420
rect 8484 28364 10780 28420
rect 10836 28364 10846 28420
rect 15250 28364 15260 28420
rect 15316 28364 15596 28420
rect 15652 28364 15932 28420
rect 15988 28364 16604 28420
rect 16660 28364 16670 28420
rect 27580 28364 29148 28420
rect 29204 28364 30044 28420
rect 30100 28364 30110 28420
rect 30258 28364 30268 28420
rect 30324 28364 33852 28420
rect 33908 28364 33918 28420
rect 16268 28308 16324 28364
rect 16258 28252 16268 28308
rect 16324 28252 16334 28308
rect 27906 28252 27916 28308
rect 27972 28252 28588 28308
rect 28644 28252 28654 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 16370 28140 16380 28196
rect 16436 28140 17276 28196
rect 17332 28140 17342 28196
rect 27318 28140 27356 28196
rect 27412 28140 27422 28196
rect 9996 27916 12460 27972
rect 12516 27916 12526 27972
rect 18050 27916 18060 27972
rect 18116 27916 30716 27972
rect 30772 27916 31500 27972
rect 31556 27916 34412 27972
rect 34468 27916 34478 27972
rect 9996 27860 10052 27916
rect 4274 27804 4284 27860
rect 4340 27804 9996 27860
rect 10052 27804 10062 27860
rect 12114 27804 12124 27860
rect 12180 27804 15148 27860
rect 15204 27804 15214 27860
rect 22306 27804 22316 27860
rect 22372 27804 23324 27860
rect 23380 27804 23390 27860
rect 30818 27804 30828 27860
rect 30884 27804 33068 27860
rect 33124 27804 33134 27860
rect 10098 27692 10108 27748
rect 10164 27692 11004 27748
rect 11060 27692 11070 27748
rect 11330 27692 11340 27748
rect 11396 27692 12348 27748
rect 12404 27692 12414 27748
rect 12898 27692 12908 27748
rect 12964 27692 17612 27748
rect 17668 27692 17678 27748
rect 21746 27692 21756 27748
rect 21812 27692 22652 27748
rect 22708 27692 22718 27748
rect 11554 27580 11564 27636
rect 11620 27580 12236 27636
rect 12292 27580 12302 27636
rect 6850 27468 6860 27524
rect 6916 27468 7868 27524
rect 7924 27468 10556 27524
rect 10612 27468 14476 27524
rect 14532 27468 14542 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 11778 27356 11788 27412
rect 11844 27356 12908 27412
rect 12964 27356 12974 27412
rect 13458 27356 13468 27412
rect 13524 27356 25676 27412
rect 25732 27356 26908 27412
rect 26852 27300 26908 27356
rect 3042 27244 3052 27300
rect 3108 27244 15260 27300
rect 15316 27244 15326 27300
rect 26852 27244 27916 27300
rect 27972 27244 28812 27300
rect 28868 27244 29372 27300
rect 29428 27244 29438 27300
rect 34738 27244 34748 27300
rect 34804 27244 35868 27300
rect 35924 27244 35934 27300
rect 0 27188 800 27216
rect 0 27132 1932 27188
rect 1988 27132 1998 27188
rect 7074 27132 7084 27188
rect 7140 27132 7532 27188
rect 7588 27132 11116 27188
rect 11172 27132 11182 27188
rect 11414 27132 11452 27188
rect 11508 27132 11518 27188
rect 14802 27132 14812 27188
rect 14868 27132 15596 27188
rect 15652 27132 16716 27188
rect 16772 27132 16782 27188
rect 21410 27132 21420 27188
rect 21476 27132 24780 27188
rect 24836 27132 25452 27188
rect 25508 27132 25518 27188
rect 34402 27132 34412 27188
rect 34468 27132 35196 27188
rect 35252 27132 35980 27188
rect 36036 27132 36046 27188
rect 0 27104 800 27132
rect 3714 27020 3724 27076
rect 3780 27020 4172 27076
rect 4228 27020 6748 27076
rect 6804 27020 6814 27076
rect 10994 27020 11004 27076
rect 11060 27020 11564 27076
rect 11620 27020 11630 27076
rect 13570 27020 13580 27076
rect 13636 27020 15932 27076
rect 15988 27020 15998 27076
rect 20514 27020 20524 27076
rect 20580 27020 21308 27076
rect 21364 27020 21374 27076
rect 21970 27020 21980 27076
rect 22036 27020 22988 27076
rect 23044 27020 25228 27076
rect 25284 27020 28588 27076
rect 28644 27020 29260 27076
rect 29316 27020 30828 27076
rect 30884 27020 30894 27076
rect 15698 26908 15708 26964
rect 15764 26908 16156 26964
rect 16212 26908 16222 26964
rect 33282 26908 33292 26964
rect 33348 26908 33572 26964
rect 33516 26852 33572 26908
rect 6850 26796 6860 26852
rect 6916 26796 7308 26852
rect 7364 26796 7374 26852
rect 20178 26796 20188 26852
rect 20244 26796 25564 26852
rect 25620 26796 25630 26852
rect 33516 26796 33964 26852
rect 34020 26796 34030 26852
rect 14130 26684 14140 26740
rect 14196 26684 14476 26740
rect 14532 26684 14542 26740
rect 15362 26684 15372 26740
rect 15428 26684 15764 26740
rect 15708 26628 15764 26684
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 15708 26572 15932 26628
rect 15988 26572 15998 26628
rect 5842 26460 5852 26516
rect 5908 26460 6972 26516
rect 7028 26460 7038 26516
rect 16230 26460 16268 26516
rect 16324 26460 16334 26516
rect 16594 26460 16604 26516
rect 16660 26460 17724 26516
rect 17780 26460 17790 26516
rect 25778 26460 25788 26516
rect 25844 26460 31388 26516
rect 31444 26460 31454 26516
rect 7074 26348 7084 26404
rect 7140 26348 7150 26404
rect 12114 26348 12124 26404
rect 12180 26348 15820 26404
rect 15876 26348 15886 26404
rect 16370 26348 16380 26404
rect 16436 26348 18060 26404
rect 18116 26348 18126 26404
rect 7084 25956 7140 26348
rect 15586 26236 15596 26292
rect 15652 26236 16268 26292
rect 16324 26236 16334 26292
rect 20850 26236 20860 26292
rect 20916 26236 22764 26292
rect 22820 26236 22830 26292
rect 12562 26124 12572 26180
rect 12628 26124 13020 26180
rect 13076 26124 13580 26180
rect 13636 26124 13646 26180
rect 15810 26124 15820 26180
rect 15876 26124 16604 26180
rect 16660 26124 16670 26180
rect 19618 26124 19628 26180
rect 19684 26124 20636 26180
rect 20692 26124 20702 26180
rect 21746 26124 21756 26180
rect 21812 26124 22988 26180
rect 23044 26124 23054 26180
rect 31714 26124 31724 26180
rect 31780 26124 33852 26180
rect 33908 26124 34412 26180
rect 34468 26124 34478 26180
rect 20636 26068 20692 26124
rect 20636 26012 22316 26068
rect 22372 26012 22382 26068
rect 7074 25900 7084 25956
rect 7140 25900 7150 25956
rect 11442 25900 11452 25956
rect 11508 25900 11564 25956
rect 11620 25900 11630 25956
rect 12002 25900 12012 25956
rect 12068 25900 12572 25956
rect 12628 25900 12638 25956
rect 17350 25900 17388 25956
rect 17444 25900 17454 25956
rect 0 25844 800 25872
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 0 25788 2044 25844
rect 2100 25788 2110 25844
rect 16930 25788 16940 25844
rect 16996 25788 21420 25844
rect 21476 25788 21486 25844
rect 26852 25788 33852 25844
rect 33908 25788 33918 25844
rect 0 25760 800 25788
rect 26852 25732 26908 25788
rect 9762 25676 9772 25732
rect 9828 25676 10332 25732
rect 10388 25676 10398 25732
rect 16818 25676 16828 25732
rect 16884 25676 17500 25732
rect 17556 25676 26908 25732
rect 27122 25676 27132 25732
rect 27188 25676 29148 25732
rect 29204 25676 29214 25732
rect 1698 25564 1708 25620
rect 1764 25564 3388 25620
rect 5842 25564 5852 25620
rect 5908 25564 7308 25620
rect 7364 25564 7374 25620
rect 7746 25564 7756 25620
rect 7812 25564 13692 25620
rect 13748 25564 13758 25620
rect 17714 25564 17724 25620
rect 17780 25564 31612 25620
rect 31668 25564 32172 25620
rect 32228 25564 32238 25620
rect 3332 25396 3388 25564
rect 4834 25452 4844 25508
rect 4900 25452 6524 25508
rect 6580 25452 6590 25508
rect 20514 25452 20524 25508
rect 20580 25452 21196 25508
rect 21252 25452 21262 25508
rect 22642 25452 22652 25508
rect 22708 25452 32396 25508
rect 32452 25452 32462 25508
rect 3332 25340 4284 25396
rect 4340 25340 5740 25396
rect 5796 25340 5806 25396
rect 15484 25340 19628 25396
rect 19684 25340 19694 25396
rect 20402 25340 20412 25396
rect 20468 25340 21420 25396
rect 21476 25340 21486 25396
rect 25554 25340 25564 25396
rect 25620 25340 27020 25396
rect 27076 25340 27086 25396
rect 3826 25228 3836 25284
rect 3892 25228 6972 25284
rect 7028 25228 7038 25284
rect 9660 25228 10780 25284
rect 10836 25228 10846 25284
rect 9660 25172 9716 25228
rect 9650 25116 9660 25172
rect 9716 25116 9726 25172
rect 12786 25116 12796 25172
rect 12852 25116 15316 25172
rect 12562 25004 12572 25060
rect 12628 25004 14924 25060
rect 14980 25004 14990 25060
rect 15260 24948 15316 25116
rect 15484 25060 15540 25340
rect 16482 25228 16492 25284
rect 16548 25228 17052 25284
rect 17108 25228 17118 25284
rect 17686 25228 17724 25284
rect 17780 25228 17790 25284
rect 19058 25228 19068 25284
rect 19124 25228 19852 25284
rect 19908 25228 20636 25284
rect 20692 25228 20702 25284
rect 20850 25228 20860 25284
rect 20916 25228 23212 25284
rect 23268 25228 23278 25284
rect 23426 25228 23436 25284
rect 23492 25228 25228 25284
rect 25284 25228 25294 25284
rect 20178 25116 20188 25172
rect 20244 25116 23996 25172
rect 24052 25116 24062 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 15474 25004 15484 25060
rect 15540 25004 15550 25060
rect 23874 25004 23884 25060
rect 23940 25004 25452 25060
rect 25508 25004 25900 25060
rect 25956 25004 25966 25060
rect 28466 25004 28476 25060
rect 28532 25004 28924 25060
rect 28980 25004 28990 25060
rect 7746 24892 7756 24948
rect 7812 24892 10556 24948
rect 10612 24892 10622 24948
rect 12674 24892 12684 24948
rect 12740 24892 13468 24948
rect 13524 24892 13534 24948
rect 13692 24892 15036 24948
rect 15092 24892 15102 24948
rect 15250 24892 15260 24948
rect 15316 24892 16604 24948
rect 16660 24892 17164 24948
rect 17220 24892 17230 24948
rect 17602 24892 17612 24948
rect 17668 24892 29372 24948
rect 29428 24892 29438 24948
rect 13692 24836 13748 24892
rect 9986 24780 9996 24836
rect 10052 24780 10780 24836
rect 10836 24780 13748 24836
rect 13906 24780 13916 24836
rect 13972 24780 18844 24836
rect 18900 24780 18910 24836
rect 28700 24780 30156 24836
rect 30212 24780 30222 24836
rect 28700 24724 28756 24780
rect 7186 24668 7196 24724
rect 7252 24668 7532 24724
rect 7588 24668 7598 24724
rect 10882 24668 10892 24724
rect 10948 24668 12572 24724
rect 12628 24668 12638 24724
rect 13458 24668 13468 24724
rect 13524 24668 14812 24724
rect 14868 24668 14878 24724
rect 16370 24668 16380 24724
rect 16436 24668 17500 24724
rect 17556 24668 23324 24724
rect 23380 24668 23884 24724
rect 23940 24668 23950 24724
rect 28690 24668 28700 24724
rect 28756 24668 28766 24724
rect 5730 24556 5740 24612
rect 5796 24556 6972 24612
rect 7028 24556 7038 24612
rect 9874 24556 9884 24612
rect 9940 24556 11116 24612
rect 11172 24556 11182 24612
rect 11666 24556 11676 24612
rect 11732 24556 16492 24612
rect 16548 24556 16558 24612
rect 18834 24556 18844 24612
rect 18900 24556 23548 24612
rect 23604 24556 23614 24612
rect 27010 24556 27020 24612
rect 27076 24556 27692 24612
rect 27748 24556 27758 24612
rect 0 24500 800 24528
rect 0 24444 1932 24500
rect 1988 24444 1998 24500
rect 5058 24444 5068 24500
rect 5124 24444 13916 24500
rect 13972 24444 13982 24500
rect 15138 24444 15148 24500
rect 15204 24444 24892 24500
rect 24948 24444 24958 24500
rect 0 24416 800 24444
rect 10070 24332 10108 24388
rect 10164 24332 13468 24388
rect 13524 24332 13534 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 33394 24108 33404 24164
rect 33460 24108 33470 24164
rect 3826 23996 3836 24052
rect 3892 23996 6860 24052
rect 6916 23996 6926 24052
rect 13570 23996 13580 24052
rect 13636 23996 16492 24052
rect 16548 23996 17500 24052
rect 17556 23996 17566 24052
rect 29362 23996 29372 24052
rect 29428 23996 29708 24052
rect 29764 23996 29774 24052
rect 8418 23884 8428 23940
rect 8484 23884 10108 23940
rect 10164 23884 10174 23940
rect 17154 23884 17164 23940
rect 17220 23884 17948 23940
rect 18004 23884 18620 23940
rect 18676 23884 19292 23940
rect 19348 23884 19358 23940
rect 33404 23828 33460 24108
rect 3332 23772 4284 23828
rect 4340 23772 5628 23828
rect 5684 23772 5694 23828
rect 7186 23772 7196 23828
rect 7252 23772 10332 23828
rect 10388 23772 16828 23828
rect 16884 23772 16894 23828
rect 29474 23772 29484 23828
rect 29540 23772 30156 23828
rect 30212 23772 30222 23828
rect 32834 23772 32844 23828
rect 32900 23772 33460 23828
rect 3332 23604 3388 23772
rect 5730 23660 5740 23716
rect 5796 23660 9772 23716
rect 9828 23660 9838 23716
rect 17826 23660 17836 23716
rect 17892 23660 33852 23716
rect 33908 23660 34860 23716
rect 34916 23660 34926 23716
rect 1698 23548 1708 23604
rect 1764 23548 3388 23604
rect 33282 23548 33292 23604
rect 33348 23548 34076 23604
rect 34132 23548 34142 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 7746 23436 7756 23492
rect 7812 23436 9996 23492
rect 10052 23436 10062 23492
rect 15138 23436 15148 23492
rect 15204 23436 16716 23492
rect 16772 23436 17500 23492
rect 17556 23436 17566 23492
rect 20178 23436 20188 23492
rect 20244 23436 22092 23492
rect 22148 23436 22158 23492
rect 29586 23436 29596 23492
rect 29652 23436 31724 23492
rect 31780 23436 31790 23492
rect 33814 23436 33852 23492
rect 33908 23436 33918 23492
rect 20188 23380 20244 23436
rect 10434 23324 10444 23380
rect 10500 23324 11452 23380
rect 11508 23324 11518 23380
rect 18386 23324 18396 23380
rect 18452 23324 20244 23380
rect 21746 23324 21756 23380
rect 21812 23324 22988 23380
rect 23044 23324 23436 23380
rect 23492 23324 23502 23380
rect 30034 23324 30044 23380
rect 30100 23324 33068 23380
rect 33124 23324 33134 23380
rect 41122 23324 41132 23380
rect 41188 23324 42812 23380
rect 42868 23324 42878 23380
rect 16594 23212 16604 23268
rect 16660 23212 17612 23268
rect 17668 23212 19292 23268
rect 19348 23212 20076 23268
rect 20132 23212 20142 23268
rect 23538 23212 23548 23268
rect 23604 23212 30380 23268
rect 30436 23212 33628 23268
rect 33684 23212 33694 23268
rect 0 23156 800 23184
rect 0 23100 1932 23156
rect 1988 23100 1998 23156
rect 12226 23100 12236 23156
rect 12292 23100 13244 23156
rect 13300 23100 13310 23156
rect 29026 23100 29036 23156
rect 29092 23100 29102 23156
rect 29362 23100 29372 23156
rect 29428 23100 29820 23156
rect 29876 23100 30156 23156
rect 30212 23100 30222 23156
rect 0 23072 800 23100
rect 29036 23044 29092 23100
rect 3602 22988 3612 23044
rect 3668 22988 4172 23044
rect 4228 22988 8316 23044
rect 8372 22988 8382 23044
rect 12002 22988 12012 23044
rect 12068 22988 18284 23044
rect 18340 22988 28028 23044
rect 28084 22988 29708 23044
rect 29764 22988 30716 23044
rect 30772 22988 30782 23044
rect 34962 22988 34972 23044
rect 35028 22988 36652 23044
rect 36708 22988 36718 23044
rect 29474 22876 29484 22932
rect 29540 22876 30604 22932
rect 30660 22876 30670 22932
rect 14466 22764 14476 22820
rect 14532 22764 15148 22820
rect 15204 22764 15214 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 10098 22652 10108 22708
rect 10164 22652 10668 22708
rect 10724 22652 19516 22708
rect 19572 22652 20748 22708
rect 20804 22652 21420 22708
rect 21476 22652 21486 22708
rect 5842 22540 5852 22596
rect 5908 22540 11340 22596
rect 11396 22540 11406 22596
rect 14690 22540 14700 22596
rect 14756 22540 22204 22596
rect 22260 22540 22270 22596
rect 26852 22540 34076 22596
rect 34132 22540 34142 22596
rect 26852 22484 26908 22540
rect 44200 22484 45000 22512
rect 6066 22428 6076 22484
rect 6132 22428 9324 22484
rect 9380 22428 9390 22484
rect 9874 22428 9884 22484
rect 9940 22428 10668 22484
rect 10724 22428 10734 22484
rect 11106 22428 11116 22484
rect 11172 22428 12012 22484
rect 12068 22428 12078 22484
rect 15026 22428 15036 22484
rect 15092 22428 26908 22484
rect 27346 22428 27356 22484
rect 27412 22428 27804 22484
rect 27860 22428 29372 22484
rect 29428 22428 29438 22484
rect 43138 22428 43148 22484
rect 43204 22428 45000 22484
rect 44200 22400 45000 22428
rect 10098 22316 10108 22372
rect 10164 22316 10332 22372
rect 10388 22316 10398 22372
rect 26898 22316 26908 22372
rect 26964 22316 27692 22372
rect 27748 22316 27758 22372
rect 30370 22316 30380 22372
rect 30436 22316 30940 22372
rect 30996 22316 31006 22372
rect 33842 22316 33852 22372
rect 33908 22316 35420 22372
rect 35476 22316 36204 22372
rect 36260 22316 36270 22372
rect 14578 22204 14588 22260
rect 14644 22204 14924 22260
rect 14980 22204 14990 22260
rect 25890 22204 25900 22260
rect 25956 22204 27132 22260
rect 27188 22204 27198 22260
rect 8306 22092 8316 22148
rect 8372 22092 10556 22148
rect 10612 22092 10622 22148
rect 11190 22092 11228 22148
rect 11284 22092 11294 22148
rect 16034 22092 16044 22148
rect 16100 22092 16492 22148
rect 16548 22092 16558 22148
rect 22754 22092 22764 22148
rect 22820 22092 25452 22148
rect 25508 22092 26012 22148
rect 26068 22092 26078 22148
rect 28466 22092 28476 22148
rect 28532 22092 29596 22148
rect 29652 22092 30380 22148
rect 30436 22092 30446 22148
rect 10882 21980 10892 22036
rect 10948 21980 11340 22036
rect 11396 21980 11406 22036
rect 27122 21980 27132 22036
rect 27188 21980 28140 22036
rect 28196 21980 28206 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 1362 21868 1372 21924
rect 1428 21868 14252 21924
rect 14308 21868 14588 21924
rect 14644 21868 14654 21924
rect 17350 21868 17388 21924
rect 17444 21868 17454 21924
rect 17602 21868 17612 21924
rect 17668 21868 18172 21924
rect 18228 21868 18238 21924
rect 27010 21868 27020 21924
rect 27076 21868 28028 21924
rect 28084 21868 28364 21924
rect 28420 21868 29148 21924
rect 29204 21868 29214 21924
rect 29362 21868 29372 21924
rect 29428 21868 29438 21924
rect 29922 21868 29932 21924
rect 29988 21868 33628 21924
rect 33684 21868 33694 21924
rect 0 21812 800 21840
rect 29372 21812 29428 21868
rect 0 21756 1932 21812
rect 1988 21756 1998 21812
rect 2706 21756 2716 21812
rect 2772 21756 15708 21812
rect 15764 21756 15774 21812
rect 15922 21756 15932 21812
rect 15988 21756 19292 21812
rect 19348 21756 19358 21812
rect 28578 21756 28588 21812
rect 28644 21756 29428 21812
rect 0 21728 800 21756
rect 3490 21644 3500 21700
rect 3556 21644 14476 21700
rect 14532 21644 14542 21700
rect 14802 21644 14812 21700
rect 14868 21644 17836 21700
rect 17892 21644 17902 21700
rect 6514 21532 6524 21588
rect 6580 21532 8988 21588
rect 9044 21532 12796 21588
rect 12852 21532 12862 21588
rect 19292 21476 19348 21756
rect 24882 21644 24892 21700
rect 24948 21644 25340 21700
rect 25396 21644 25406 21700
rect 26684 21644 27356 21700
rect 27412 21644 27422 21700
rect 26684 21588 26740 21644
rect 24322 21532 24332 21588
rect 24388 21532 25676 21588
rect 25732 21532 25742 21588
rect 26674 21532 26684 21588
rect 26740 21532 26750 21588
rect 28130 21532 28140 21588
rect 28196 21532 28812 21588
rect 28868 21532 28878 21588
rect 5170 21420 5180 21476
rect 5236 21420 10220 21476
rect 10276 21420 10286 21476
rect 14354 21420 14364 21476
rect 14420 21420 14924 21476
rect 14980 21420 15596 21476
rect 15652 21420 15662 21476
rect 16790 21420 16828 21476
rect 16884 21420 17500 21476
rect 17556 21420 17566 21476
rect 19292 21420 27244 21476
rect 27300 21420 27310 21476
rect 3938 21308 3948 21364
rect 4004 21308 6076 21364
rect 6132 21308 11228 21364
rect 11284 21308 11294 21364
rect 17602 21308 17612 21364
rect 17668 21308 22316 21364
rect 22372 21308 24220 21364
rect 24276 21308 26684 21364
rect 26740 21308 26750 21364
rect 27458 21308 27468 21364
rect 27524 21308 28028 21364
rect 28084 21308 28094 21364
rect 8530 21196 8540 21252
rect 8596 21196 9996 21252
rect 10052 21196 10062 21252
rect 10546 21196 10556 21252
rect 10612 21196 11788 21252
rect 11844 21196 11854 21252
rect 15250 21196 15260 21252
rect 15316 21196 31276 21252
rect 31332 21196 31836 21252
rect 31892 21196 31902 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 12898 21084 12908 21140
rect 12964 21084 13580 21140
rect 13636 21084 17388 21140
rect 17444 21084 17454 21140
rect 17602 21084 17612 21140
rect 17668 21084 27524 21140
rect 1698 20972 1708 21028
rect 1764 20972 3388 21028
rect 7410 20972 7420 21028
rect 7476 20972 11788 21028
rect 11844 20972 11854 21028
rect 15922 20972 15932 21028
rect 15988 20972 16268 21028
rect 16324 20972 27412 21028
rect 3332 20804 3388 20972
rect 3826 20860 3836 20916
rect 3892 20860 10332 20916
rect 10388 20860 10398 20916
rect 13458 20860 13468 20916
rect 13524 20860 15596 20916
rect 15652 20860 15662 20916
rect 15810 20860 15820 20916
rect 15876 20860 21868 20916
rect 21924 20860 21934 20916
rect 23314 20860 23324 20916
rect 23380 20860 26852 20916
rect 26796 20804 26852 20860
rect 3332 20748 4284 20804
rect 4340 20748 5068 20804
rect 5124 20748 5134 20804
rect 12562 20748 12572 20804
rect 12628 20748 13356 20804
rect 13412 20748 14812 20804
rect 14868 20748 14878 20804
rect 15698 20748 15708 20804
rect 15764 20748 17500 20804
rect 17556 20748 17566 20804
rect 17826 20748 17836 20804
rect 17892 20748 18844 20804
rect 18900 20748 18910 20804
rect 23090 20748 23100 20804
rect 23156 20748 24556 20804
rect 24612 20748 24622 20804
rect 26786 20748 26796 20804
rect 26852 20748 27132 20804
rect 27188 20748 27198 20804
rect 17836 20692 17892 20748
rect 27356 20692 27412 20972
rect 27468 20916 27524 21084
rect 27682 20972 27692 21028
rect 27748 20972 28364 21028
rect 28420 20972 28812 21028
rect 28868 20972 30268 21028
rect 30324 20972 30334 21028
rect 27468 20860 28588 20916
rect 28644 20860 30380 20916
rect 30436 20860 30716 20916
rect 30772 20860 30782 20916
rect 30930 20860 30940 20916
rect 30996 20860 31612 20916
rect 31668 20860 35644 20916
rect 35700 20860 35710 20916
rect 29250 20748 29260 20804
rect 29316 20748 30268 20804
rect 30324 20748 30334 20804
rect 7522 20636 7532 20692
rect 7588 20636 10108 20692
rect 10164 20636 10780 20692
rect 10836 20636 10846 20692
rect 17154 20636 17164 20692
rect 17220 20636 17892 20692
rect 22082 20636 22092 20692
rect 22148 20636 22652 20692
rect 22708 20636 23772 20692
rect 23828 20636 23838 20692
rect 27356 20636 29596 20692
rect 29652 20636 30044 20692
rect 30100 20636 30110 20692
rect 11442 20524 11452 20580
rect 11508 20524 14476 20580
rect 14532 20524 14542 20580
rect 25666 20524 25676 20580
rect 25732 20524 40348 20580
rect 40404 20524 40414 20580
rect 0 20468 800 20496
rect 0 20412 1932 20468
rect 1988 20412 1998 20468
rect 0 20384 800 20412
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 26852 20300 35084 20356
rect 35140 20300 35150 20356
rect 26852 20244 26908 20300
rect 11554 20188 11564 20244
rect 11620 20188 12012 20244
rect 12068 20188 12078 20244
rect 13794 20188 13804 20244
rect 13860 20188 26908 20244
rect 30370 20188 30380 20244
rect 30436 20188 33852 20244
rect 33908 20188 33918 20244
rect 13346 20076 13356 20132
rect 13412 20076 13916 20132
rect 13972 20076 13982 20132
rect 14354 20076 14364 20132
rect 14420 20076 15148 20132
rect 21634 20076 21644 20132
rect 21700 20076 22988 20132
rect 23044 20076 23054 20132
rect 15092 20020 15148 20076
rect 23492 20020 23548 20132
rect 23604 20076 28028 20132
rect 28084 20076 29036 20132
rect 29092 20076 29102 20132
rect 34178 20076 34188 20132
rect 34244 20076 35420 20132
rect 35476 20076 35486 20132
rect 8082 19964 8092 20020
rect 8148 19964 9548 20020
rect 9604 19964 9614 20020
rect 9874 19964 9884 20020
rect 9940 19964 10108 20020
rect 10164 19964 11676 20020
rect 11732 19964 13132 20020
rect 13188 19964 14924 20020
rect 14980 19964 14990 20020
rect 15092 19964 15260 20020
rect 15316 19964 16044 20020
rect 16100 19964 16110 20020
rect 23090 19964 23100 20020
rect 23156 19964 23548 20020
rect 26852 19964 31724 20020
rect 31780 19964 32508 20020
rect 32564 19964 32574 20020
rect 34962 19964 34972 20020
rect 35028 19964 38220 20020
rect 38276 19964 38286 20020
rect 3826 19852 3836 19908
rect 3892 19852 15148 19908
rect 15698 19852 15708 19908
rect 15764 19852 16828 19908
rect 16884 19852 20188 19908
rect 20244 19852 20254 19908
rect 22754 19852 22764 19908
rect 22820 19852 23884 19908
rect 23940 19852 23950 19908
rect 15092 19796 15148 19852
rect 15708 19796 15764 19852
rect 26852 19796 26908 19964
rect 29362 19852 29372 19908
rect 29428 19852 31500 19908
rect 31556 19852 31566 19908
rect 12338 19740 12348 19796
rect 12404 19740 13804 19796
rect 13860 19740 14700 19796
rect 14756 19740 14766 19796
rect 15092 19740 15764 19796
rect 17490 19740 17500 19796
rect 17556 19740 26908 19796
rect 28466 19740 28476 19796
rect 28532 19740 29260 19796
rect 29316 19740 29484 19796
rect 29540 19740 29550 19796
rect 19618 19628 19628 19684
rect 19684 19628 20524 19684
rect 20580 19628 24556 19684
rect 24612 19628 24622 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 21970 19516 21980 19572
rect 22036 19516 23436 19572
rect 23492 19516 24108 19572
rect 24164 19516 24174 19572
rect 12674 19404 12684 19460
rect 12740 19404 13244 19460
rect 13300 19404 13310 19460
rect 13682 19404 13692 19460
rect 13748 19404 14700 19460
rect 14756 19404 14766 19460
rect 22306 19404 22316 19460
rect 22372 19404 22652 19460
rect 22708 19404 22718 19460
rect 23090 19404 23100 19460
rect 23156 19404 23772 19460
rect 23828 19404 23838 19460
rect 34850 19404 34860 19460
rect 34916 19404 36204 19460
rect 36260 19404 36270 19460
rect 1922 19292 1932 19348
rect 1988 19292 1998 19348
rect 13906 19292 13916 19348
rect 13972 19292 15036 19348
rect 15092 19292 15102 19348
rect 20290 19292 20300 19348
rect 20356 19292 20748 19348
rect 20804 19292 22204 19348
rect 22260 19292 22270 19348
rect 22418 19292 22428 19348
rect 22484 19292 22522 19348
rect 22866 19292 22876 19348
rect 22932 19292 24332 19348
rect 24388 19292 24398 19348
rect 27234 19292 27244 19348
rect 27300 19292 28588 19348
rect 28644 19292 29148 19348
rect 29204 19292 29214 19348
rect 34962 19292 34972 19348
rect 35028 19292 36428 19348
rect 36484 19292 36494 19348
rect 0 19124 800 19152
rect 1932 19124 1988 19292
rect 7298 19180 7308 19236
rect 7364 19180 12236 19236
rect 12292 19180 12302 19236
rect 13570 19180 13580 19236
rect 13636 19180 14812 19236
rect 14868 19180 14878 19236
rect 18722 19180 18732 19236
rect 18788 19180 23884 19236
rect 23940 19180 24780 19236
rect 24836 19180 27020 19236
rect 27076 19180 28140 19236
rect 28196 19180 28206 19236
rect 32498 19180 32508 19236
rect 32564 19180 35084 19236
rect 35140 19180 35150 19236
rect 35634 19180 35644 19236
rect 35700 19180 37100 19236
rect 37156 19180 37166 19236
rect 0 19068 1988 19124
rect 5730 19068 5740 19124
rect 5796 19068 6412 19124
rect 6468 19068 7868 19124
rect 7924 19068 7934 19124
rect 11554 19068 11564 19124
rect 11620 19068 13580 19124
rect 13636 19068 15372 19124
rect 15428 19068 15438 19124
rect 18162 19068 18172 19124
rect 18228 19068 19516 19124
rect 19572 19068 19582 19124
rect 20738 19068 20748 19124
rect 20804 19068 21532 19124
rect 21588 19068 21598 19124
rect 22082 19068 22092 19124
rect 22148 19068 23772 19124
rect 23828 19068 23838 19124
rect 32386 19068 32396 19124
rect 32452 19068 33740 19124
rect 33796 19068 33806 19124
rect 0 19040 800 19068
rect 10546 18956 10556 19012
rect 10612 18956 15708 19012
rect 15764 18956 16940 19012
rect 16996 18956 17612 19012
rect 17668 18956 17678 19012
rect 17948 18956 21196 19012
rect 21252 18956 21262 19012
rect 33282 18956 33292 19012
rect 33348 18956 34748 19012
rect 34804 18956 34814 19012
rect 17948 18900 18004 18956
rect 11554 18844 11564 18900
rect 11620 18844 12460 18900
rect 12516 18844 13692 18900
rect 13748 18844 13758 18900
rect 17938 18844 17948 18900
rect 18004 18844 18014 18900
rect 18508 18844 19068 18900
rect 19124 18844 19134 18900
rect 22278 18844 22316 18900
rect 22372 18844 22382 18900
rect 18508 18788 18564 18844
rect 13206 18732 13244 18788
rect 13300 18732 13310 18788
rect 16034 18732 16044 18788
rect 16100 18732 16492 18788
rect 16548 18732 18564 18788
rect 18694 18732 18732 18788
rect 18788 18732 18798 18788
rect 7634 18620 7644 18676
rect 7700 18620 8092 18676
rect 8148 18620 8158 18676
rect 9650 18620 9660 18676
rect 9716 18620 14028 18676
rect 14084 18620 15820 18676
rect 15876 18620 15886 18676
rect 19068 18564 19124 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 22754 18620 22764 18676
rect 22820 18620 23324 18676
rect 23380 18620 23390 18676
rect 38322 18620 38332 18676
rect 38388 18620 38668 18676
rect 38612 18564 38668 18620
rect 7858 18508 7868 18564
rect 7924 18508 9996 18564
rect 10052 18508 10062 18564
rect 11442 18508 11452 18564
rect 11508 18508 12964 18564
rect 14690 18508 14700 18564
rect 14756 18508 15484 18564
rect 15540 18508 15550 18564
rect 19068 18508 23548 18564
rect 23604 18508 23614 18564
rect 27794 18508 27804 18564
rect 27860 18508 30828 18564
rect 30884 18508 30894 18564
rect 31602 18508 31612 18564
rect 31668 18508 31678 18564
rect 38612 18508 39340 18564
rect 39396 18508 39406 18564
rect 12908 18452 12964 18508
rect 1698 18396 1708 18452
rect 1764 18396 4732 18452
rect 4788 18396 4798 18452
rect 5506 18396 5516 18452
rect 5572 18396 6636 18452
rect 6692 18396 7196 18452
rect 7252 18396 7262 18452
rect 12908 18396 13468 18452
rect 13524 18396 14252 18452
rect 14308 18396 14318 18452
rect 16258 18396 16268 18452
rect 16324 18396 17164 18452
rect 17220 18396 17388 18452
rect 17444 18396 17454 18452
rect 20290 18396 20300 18452
rect 20356 18396 21196 18452
rect 21252 18396 21262 18452
rect 21858 18396 21868 18452
rect 21924 18396 26012 18452
rect 26068 18396 26078 18452
rect 31612 18340 31668 18508
rect 32050 18396 32060 18452
rect 32116 18396 33180 18452
rect 33236 18396 34188 18452
rect 34244 18396 34972 18452
rect 35028 18396 35420 18452
rect 35476 18396 35486 18452
rect 2370 18284 2380 18340
rect 2436 18284 3164 18340
rect 3220 18284 3230 18340
rect 3826 18284 3836 18340
rect 3892 18284 4508 18340
rect 4564 18284 6300 18340
rect 6356 18284 6366 18340
rect 17938 18284 17948 18340
rect 18004 18284 18396 18340
rect 18452 18284 20636 18340
rect 20692 18284 20702 18340
rect 31612 18284 33068 18340
rect 33124 18284 33134 18340
rect 2034 18172 2044 18228
rect 2100 18172 9548 18228
rect 9604 18172 10220 18228
rect 10276 18172 10286 18228
rect 16706 18172 16716 18228
rect 16772 18172 18508 18228
rect 18564 18172 19292 18228
rect 19348 18172 19358 18228
rect 5394 18060 5404 18116
rect 5460 18060 7532 18116
rect 7588 18060 7598 18116
rect 15698 18060 15708 18116
rect 15764 18060 17500 18116
rect 17556 18060 19068 18116
rect 19124 18060 19134 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 5058 17948 5068 18004
rect 5124 17948 7308 18004
rect 7364 17948 8316 18004
rect 8372 17948 8382 18004
rect 9538 17948 9548 18004
rect 9604 17948 14364 18004
rect 14420 17948 14430 18004
rect 20402 17948 20412 18004
rect 20468 17948 21644 18004
rect 21700 17948 21710 18004
rect 3490 17836 3500 17892
rect 3556 17836 3948 17892
rect 4004 17836 4014 17892
rect 4162 17836 4172 17892
rect 4228 17836 5516 17892
rect 5572 17836 5582 17892
rect 16930 17836 16940 17892
rect 16996 17836 17836 17892
rect 17892 17836 17902 17892
rect 0 17780 800 17808
rect 0 17724 1708 17780
rect 1764 17724 1774 17780
rect 1922 17724 1932 17780
rect 1988 17724 3276 17780
rect 3332 17724 6076 17780
rect 6132 17724 6142 17780
rect 21830 17724 21868 17780
rect 21924 17724 21934 17780
rect 22306 17724 22316 17780
rect 22372 17724 25564 17780
rect 25620 17724 28588 17780
rect 28644 17724 30828 17780
rect 30884 17724 31500 17780
rect 31556 17724 31566 17780
rect 0 17696 800 17724
rect 4274 17612 4284 17668
rect 4340 17612 5068 17668
rect 5124 17612 5134 17668
rect 5282 17612 5292 17668
rect 5348 17612 5852 17668
rect 5908 17612 6636 17668
rect 6692 17612 6702 17668
rect 6850 17612 6860 17668
rect 6916 17612 7420 17668
rect 7476 17612 7868 17668
rect 7924 17612 7934 17668
rect 17378 17612 17388 17668
rect 17444 17612 18844 17668
rect 18900 17612 18910 17668
rect 6860 17556 6916 17612
rect 2258 17500 2268 17556
rect 2324 17500 4172 17556
rect 4228 17500 6916 17556
rect 16146 17500 16156 17556
rect 16212 17500 16716 17556
rect 16772 17500 25116 17556
rect 25172 17500 25182 17556
rect 13542 17388 13580 17444
rect 13636 17388 13646 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 4498 17164 4508 17220
rect 4564 17164 6020 17220
rect 5964 17108 6020 17164
rect 2930 17052 2940 17108
rect 2996 17052 5292 17108
rect 5348 17052 5358 17108
rect 5964 17052 6524 17108
rect 6580 17052 9660 17108
rect 9716 17052 9726 17108
rect 11778 17052 11788 17108
rect 11844 17052 13692 17108
rect 13748 17052 13758 17108
rect 17042 17052 17052 17108
rect 17108 17052 17724 17108
rect 17780 17052 18732 17108
rect 18788 17052 18798 17108
rect 22194 17052 22204 17108
rect 22260 17052 27356 17108
rect 27412 17052 27422 17108
rect 28130 17052 28140 17108
rect 28196 17052 28812 17108
rect 28868 17052 29260 17108
rect 29316 17052 29326 17108
rect 30258 17052 30268 17108
rect 30324 17052 33292 17108
rect 33348 17052 33358 17108
rect 3266 16940 3276 16996
rect 3332 16940 4396 16996
rect 4452 16940 4462 16996
rect 5842 16940 5852 16996
rect 5908 16940 6860 16996
rect 6916 16940 7532 16996
rect 7588 16940 7598 16996
rect 17938 16940 17948 16996
rect 18004 16940 18508 16996
rect 18564 16940 18574 16996
rect 20962 16940 20972 16996
rect 21028 16940 21868 16996
rect 21924 16940 22764 16996
rect 22820 16940 22830 16996
rect 2258 16828 2268 16884
rect 2324 16828 3836 16884
rect 3892 16828 3902 16884
rect 4274 16828 4284 16884
rect 4340 16828 4350 16884
rect 5730 16828 5740 16884
rect 5796 16828 6972 16884
rect 7028 16828 7038 16884
rect 7186 16828 7196 16884
rect 7252 16828 9884 16884
rect 9940 16828 9950 16884
rect 14662 16828 14700 16884
rect 14756 16828 14766 16884
rect 14914 16828 14924 16884
rect 14980 16828 17612 16884
rect 17668 16828 17678 16884
rect 18722 16828 18732 16884
rect 18788 16828 19628 16884
rect 19684 16828 19694 16884
rect 22418 16828 22428 16884
rect 22484 16828 22652 16884
rect 22708 16828 22718 16884
rect 23548 16828 28700 16884
rect 28756 16828 29148 16884
rect 29204 16828 29214 16884
rect 4284 16772 4340 16828
rect 23548 16772 23604 16828
rect 2146 16716 2156 16772
rect 2212 16716 4340 16772
rect 4610 16716 4620 16772
rect 4676 16716 8540 16772
rect 8596 16716 8606 16772
rect 13346 16716 13356 16772
rect 13412 16716 15148 16772
rect 15204 16716 15214 16772
rect 16258 16716 16268 16772
rect 16324 16716 23604 16772
rect 27906 16716 27916 16772
rect 27972 16716 28924 16772
rect 28980 16716 28990 16772
rect 10546 16604 10556 16660
rect 10612 16604 13020 16660
rect 13076 16604 17276 16660
rect 17332 16604 17342 16660
rect 10892 16548 10948 16604
rect 10882 16492 10892 16548
rect 10948 16492 10958 16548
rect 14914 16492 14924 16548
rect 14980 16492 16604 16548
rect 16660 16492 26908 16548
rect 26964 16492 26974 16548
rect 0 16436 800 16464
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16380 2380 16436
rect 2436 16380 2446 16436
rect 6290 16380 6300 16436
rect 6356 16380 9100 16436
rect 9156 16380 17388 16436
rect 17444 16380 17454 16436
rect 17602 16380 17612 16436
rect 17668 16380 17706 16436
rect 0 16352 800 16380
rect 3938 16268 3948 16324
rect 4004 16268 4844 16324
rect 4900 16268 4910 16324
rect 10098 16268 10108 16324
rect 10164 16268 11116 16324
rect 11172 16268 11182 16324
rect 2594 16156 2604 16212
rect 2660 16156 4172 16212
rect 4228 16156 4238 16212
rect 4498 16156 4508 16212
rect 4564 16156 5852 16212
rect 5908 16156 5918 16212
rect 10770 16156 10780 16212
rect 10836 16156 11228 16212
rect 11284 16156 11294 16212
rect 12562 16156 12572 16212
rect 12628 16156 16604 16212
rect 16660 16156 28476 16212
rect 28532 16156 28542 16212
rect 1922 16044 1932 16100
rect 1988 16044 3052 16100
rect 3108 16044 3118 16100
rect 3266 16044 3276 16100
rect 3332 16044 3948 16100
rect 4004 16044 4014 16100
rect 4722 16044 4732 16100
rect 4788 16044 4798 16100
rect 11890 16044 11900 16100
rect 11956 16044 12908 16100
rect 12964 16044 14140 16100
rect 14196 16044 14206 16100
rect 26338 16044 26348 16100
rect 26404 16044 28028 16100
rect 28084 16044 28094 16100
rect 4732 15988 4788 16044
rect 2930 15932 2940 15988
rect 2996 15932 4788 15988
rect 5058 15932 5068 15988
rect 5124 15932 11452 15988
rect 11508 15932 11518 15988
rect 26852 15932 29148 15988
rect 29204 15932 29214 15988
rect 26852 15876 26908 15932
rect 3378 15820 3388 15876
rect 3444 15820 5740 15876
rect 5796 15820 5806 15876
rect 18274 15820 18284 15876
rect 18340 15820 25900 15876
rect 25956 15820 26908 15876
rect 27570 15820 27580 15876
rect 27636 15820 28140 15876
rect 28196 15820 28206 15876
rect 3500 15316 3556 15820
rect 12450 15708 12460 15764
rect 12516 15708 13132 15764
rect 13188 15708 15372 15764
rect 15428 15708 16268 15764
rect 16324 15708 16334 15764
rect 18722 15708 18732 15764
rect 18788 15708 18844 15764
rect 18900 15708 18910 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 17490 15596 17500 15652
rect 17556 15596 18508 15652
rect 18564 15596 18574 15652
rect 11106 15484 11116 15540
rect 11172 15484 11676 15540
rect 11732 15484 11742 15540
rect 17714 15484 17724 15540
rect 17780 15484 18284 15540
rect 18340 15484 20188 15540
rect 20244 15484 20254 15540
rect 20850 15484 20860 15540
rect 20916 15484 21532 15540
rect 21588 15484 22876 15540
rect 22932 15484 22942 15540
rect 29698 15484 29708 15540
rect 29764 15484 32396 15540
rect 32452 15484 32462 15540
rect 15586 15372 15596 15428
rect 15652 15372 16828 15428
rect 16884 15372 18060 15428
rect 18116 15372 18126 15428
rect 3490 15260 3500 15316
rect 3556 15260 3566 15316
rect 4162 15260 4172 15316
rect 4228 15260 5740 15316
rect 5796 15260 6076 15316
rect 6132 15260 6142 15316
rect 7746 15260 7756 15316
rect 7812 15260 9772 15316
rect 9828 15260 9838 15316
rect 11330 15260 11340 15316
rect 11396 15260 11900 15316
rect 11956 15260 11966 15316
rect 25554 15260 25564 15316
rect 25620 15260 26572 15316
rect 26628 15260 26638 15316
rect 27010 15260 27020 15316
rect 27076 15260 27356 15316
rect 27412 15260 27422 15316
rect 11778 15148 11788 15204
rect 11844 15148 12684 15204
rect 12740 15148 12750 15204
rect 16818 15148 16828 15204
rect 16884 15148 17164 15204
rect 17220 15148 17388 15204
rect 17444 15148 17454 15204
rect 25778 15148 25788 15204
rect 25844 15148 27468 15204
rect 27524 15148 27534 15204
rect 27794 15148 27804 15204
rect 27860 15148 30380 15204
rect 30436 15148 30446 15204
rect 0 15092 800 15120
rect 0 15036 1708 15092
rect 1764 15036 1774 15092
rect 1922 15036 1932 15092
rect 1988 15036 3052 15092
rect 3108 15036 3118 15092
rect 3276 15036 3836 15092
rect 3892 15036 5628 15092
rect 5684 15036 7644 15092
rect 7700 15036 7710 15092
rect 10210 15036 10220 15092
rect 10276 15036 11116 15092
rect 11172 15036 11182 15092
rect 0 15008 800 15036
rect 3276 14980 3332 15036
rect 2594 14924 2604 14980
rect 2660 14924 3332 14980
rect 15092 14924 25340 14980
rect 25396 14924 26348 14980
rect 26404 14924 26414 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 15092 14868 15148 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 8372 14812 15148 14868
rect 22642 14812 22652 14868
rect 22708 14812 23324 14868
rect 23380 14812 23390 14868
rect 8372 14756 8428 14812
rect 2258 14700 2268 14756
rect 2324 14700 5964 14756
rect 6020 14700 8428 14756
rect 8754 14700 8764 14756
rect 8820 14700 9996 14756
rect 10052 14700 14700 14756
rect 14756 14700 14766 14756
rect 15092 14700 28700 14756
rect 28756 14700 29708 14756
rect 29764 14700 29774 14756
rect 15092 14644 15148 14700
rect 4274 14588 4284 14644
rect 4340 14588 5068 14644
rect 5124 14588 6412 14644
rect 6468 14588 7420 14644
rect 7476 14588 8652 14644
rect 8708 14588 8718 14644
rect 10882 14588 10892 14644
rect 10948 14588 11228 14644
rect 11284 14588 11294 14644
rect 13916 14588 14588 14644
rect 14644 14588 15148 14644
rect 20514 14588 20524 14644
rect 20580 14588 24220 14644
rect 24276 14588 24286 14644
rect 27682 14588 27692 14644
rect 27748 14588 27758 14644
rect 13916 14532 13972 14588
rect 12450 14476 12460 14532
rect 12516 14476 13356 14532
rect 13412 14476 13422 14532
rect 13906 14476 13916 14532
rect 13972 14476 13982 14532
rect 14802 14476 14812 14532
rect 14868 14476 15820 14532
rect 15876 14476 15886 14532
rect 19618 14476 19628 14532
rect 19684 14476 21196 14532
rect 21252 14476 21262 14532
rect 21634 14476 21644 14532
rect 21700 14476 22540 14532
rect 22596 14476 25676 14532
rect 25732 14476 25742 14532
rect 13570 14364 13580 14420
rect 13636 14364 14700 14420
rect 14756 14364 15260 14420
rect 15316 14364 15326 14420
rect 26898 14364 26908 14420
rect 26964 14364 27356 14420
rect 27412 14364 27422 14420
rect 27692 14308 27748 14588
rect 2146 14252 2156 14308
rect 2212 14252 9996 14308
rect 10052 14252 10062 14308
rect 11890 14252 11900 14308
rect 11956 14252 12348 14308
rect 12404 14252 12414 14308
rect 14466 14252 14476 14308
rect 14532 14252 22876 14308
rect 22932 14252 22942 14308
rect 26114 14252 26124 14308
rect 26180 14252 27748 14308
rect 28130 14252 28140 14308
rect 28196 14252 29260 14308
rect 29316 14252 29820 14308
rect 29876 14252 29886 14308
rect 2482 14140 2492 14196
rect 2548 14140 3388 14196
rect 3444 14140 4508 14196
rect 4564 14140 4574 14196
rect 21858 14140 21868 14196
rect 21924 14140 22092 14196
rect 22148 14140 23212 14196
rect 23268 14140 27132 14196
rect 27188 14140 27804 14196
rect 27860 14140 27870 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 10994 14028 11004 14084
rect 11060 14028 11900 14084
rect 11956 14028 19068 14084
rect 19124 14028 19134 14084
rect 24210 14028 24220 14084
rect 24276 14028 26348 14084
rect 26404 14028 28252 14084
rect 28308 14028 28318 14084
rect 1698 13916 1708 13972
rect 1764 13916 2716 13972
rect 2772 13916 2782 13972
rect 9986 13916 9996 13972
rect 10052 13916 10444 13972
rect 10500 13916 25676 13972
rect 25732 13916 25742 13972
rect 39442 13916 39452 13972
rect 39508 13916 42812 13972
rect 42868 13916 42878 13972
rect 3154 13804 3164 13860
rect 3220 13804 17724 13860
rect 17780 13804 18060 13860
rect 18116 13804 22540 13860
rect 22596 13804 22606 13860
rect 26002 13804 26012 13860
rect 26068 13804 26460 13860
rect 26516 13804 30156 13860
rect 30212 13804 30222 13860
rect 0 13748 800 13776
rect 0 13692 1820 13748
rect 1876 13692 1886 13748
rect 22082 13692 22092 13748
rect 22148 13692 22652 13748
rect 22708 13692 27020 13748
rect 27076 13692 29372 13748
rect 29428 13692 29438 13748
rect 0 13664 800 13692
rect 3266 13580 3276 13636
rect 3332 13580 3948 13636
rect 4004 13580 4014 13636
rect 44200 13524 45000 13552
rect 15250 13468 15260 13524
rect 15316 13468 15820 13524
rect 15876 13468 16604 13524
rect 16660 13468 33404 13524
rect 33460 13468 33470 13524
rect 42578 13468 42588 13524
rect 42644 13468 43148 13524
rect 43204 13468 45000 13524
rect 44200 13440 45000 13468
rect 5730 13356 5740 13412
rect 5796 13356 9548 13412
rect 9604 13356 9614 13412
rect 16930 13356 16940 13412
rect 16996 13356 18396 13412
rect 18452 13356 18462 13412
rect 26226 13356 26236 13412
rect 26292 13356 27468 13412
rect 27524 13356 27534 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 14690 13244 14700 13300
rect 14756 13244 24108 13300
rect 24164 13244 25452 13300
rect 25508 13244 25518 13300
rect 3490 13132 3500 13188
rect 3556 13132 4284 13188
rect 4340 13132 17164 13188
rect 17220 13132 17612 13188
rect 17668 13132 20748 13188
rect 20804 13132 21308 13188
rect 21364 13132 21374 13188
rect 1250 13020 1260 13076
rect 1316 13020 5852 13076
rect 5908 13020 5918 13076
rect 6626 13020 6636 13076
rect 6692 13020 6972 13076
rect 7028 13020 7084 13076
rect 7140 13020 7150 13076
rect 10882 13020 10892 13076
rect 10948 13020 11228 13076
rect 11284 13020 11294 13076
rect 16706 13020 16716 13076
rect 16772 13020 18508 13076
rect 18564 13020 18574 13076
rect 23492 13020 32732 13076
rect 32788 13020 32798 13076
rect 23492 12964 23548 13020
rect 15586 12908 15596 12964
rect 15652 12908 23548 12964
rect 26674 12908 26684 12964
rect 26740 12908 27244 12964
rect 27300 12908 27310 12964
rect 2594 12796 2604 12852
rect 2660 12796 3052 12852
rect 3108 12796 3500 12852
rect 3556 12796 3566 12852
rect 5814 12796 5852 12852
rect 5908 12796 5918 12852
rect 7084 12796 14084 12852
rect 14242 12796 14252 12852
rect 14308 12796 15036 12852
rect 15092 12796 28140 12852
rect 28196 12796 28206 12852
rect 7084 12740 7140 12796
rect 14028 12740 14084 12796
rect 7074 12684 7084 12740
rect 7140 12684 7150 12740
rect 13122 12684 13132 12740
rect 13188 12684 13692 12740
rect 13748 12684 13758 12740
rect 14028 12684 18732 12740
rect 18788 12684 18798 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 8372 12460 15708 12516
rect 15764 12460 15774 12516
rect 17266 12460 17276 12516
rect 17332 12460 17612 12516
rect 17668 12460 17678 12516
rect 0 12404 800 12432
rect 8372 12404 8428 12460
rect 0 12348 2716 12404
rect 2772 12348 2782 12404
rect 6290 12348 6300 12404
rect 6356 12348 7756 12404
rect 7812 12348 8428 12404
rect 10546 12348 10556 12404
rect 10612 12348 11228 12404
rect 11284 12348 17444 12404
rect 17602 12348 17612 12404
rect 17668 12348 18620 12404
rect 18676 12348 20412 12404
rect 20468 12348 20478 12404
rect 24098 12348 24108 12404
rect 24164 12348 26348 12404
rect 26404 12348 27132 12404
rect 27188 12348 27198 12404
rect 0 12320 800 12348
rect 17388 12292 17444 12348
rect 11666 12236 11676 12292
rect 11732 12236 15932 12292
rect 15988 12236 16716 12292
rect 16772 12236 16782 12292
rect 17388 12236 21756 12292
rect 21812 12236 21822 12292
rect 2258 12124 2268 12180
rect 2324 12124 6972 12180
rect 7028 12124 7038 12180
rect 13906 12124 13916 12180
rect 13972 12124 14700 12180
rect 14756 12124 14766 12180
rect 16818 12124 16828 12180
rect 16884 12124 17836 12180
rect 17892 12124 17902 12180
rect 5730 12012 5740 12068
rect 5796 12012 6188 12068
rect 6244 12012 6254 12068
rect 8306 12012 8316 12068
rect 8372 12012 9660 12068
rect 9716 12012 9726 12068
rect 4162 11900 4172 11956
rect 4228 11900 5516 11956
rect 5572 11900 5582 11956
rect 6066 11900 6076 11956
rect 6132 11900 7084 11956
rect 7140 11900 7150 11956
rect 7410 11900 7420 11956
rect 7476 11900 8428 11956
rect 8866 11900 8876 11956
rect 8932 11900 10444 11956
rect 10500 11900 10892 11956
rect 10948 11900 10958 11956
rect 8372 11844 8428 11900
rect 4946 11788 4956 11844
rect 5012 11788 5852 11844
rect 5908 11788 5918 11844
rect 8372 11788 10668 11844
rect 10724 11788 12908 11844
rect 12964 11788 12974 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 11900 11732 11956 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 1698 11676 1708 11732
rect 1764 11676 3164 11732
rect 3220 11676 3230 11732
rect 8082 11676 8092 11732
rect 8148 11676 10108 11732
rect 10164 11676 10174 11732
rect 11890 11676 11900 11732
rect 11956 11676 11966 11732
rect 27234 11676 27244 11732
rect 27300 11676 28476 11732
rect 28532 11676 29372 11732
rect 29428 11676 29438 11732
rect 1586 11564 1596 11620
rect 1652 11564 7196 11620
rect 7252 11564 7262 11620
rect 4834 11340 4844 11396
rect 4900 11340 6636 11396
rect 6692 11340 7532 11396
rect 7588 11340 10668 11396
rect 10724 11340 13692 11396
rect 13748 11340 14476 11396
rect 14532 11340 14542 11396
rect 2930 11228 2940 11284
rect 2996 11228 6188 11284
rect 6244 11228 6254 11284
rect 8754 11228 8764 11284
rect 8820 11228 10892 11284
rect 10948 11228 12012 11284
rect 12068 11228 12078 11284
rect 12338 11228 12348 11284
rect 12404 11228 14028 11284
rect 14084 11228 14094 11284
rect 3042 11116 3052 11172
rect 3108 11116 5852 11172
rect 5908 11116 5918 11172
rect 6290 11116 6300 11172
rect 6356 11116 6860 11172
rect 6916 11116 6926 11172
rect 10994 11116 11004 11172
rect 11060 11116 11564 11172
rect 11620 11116 11630 11172
rect 17238 11116 17276 11172
rect 17332 11116 17342 11172
rect 22054 11116 22092 11172
rect 22148 11116 22158 11172
rect 0 11060 800 11088
rect 0 11004 1708 11060
rect 1764 11004 1774 11060
rect 0 10976 800 11004
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 7186 10892 7196 10948
rect 7252 10892 7756 10948
rect 7812 10892 7822 10948
rect 21186 10892 21196 10948
rect 21252 10892 22092 10948
rect 22148 10892 22158 10948
rect 6738 10780 6748 10836
rect 6804 10780 9996 10836
rect 10052 10780 10062 10836
rect 15362 10780 15372 10836
rect 15428 10780 16940 10836
rect 16996 10780 17006 10836
rect 17378 10780 17388 10836
rect 17444 10780 18172 10836
rect 18228 10780 18238 10836
rect 22194 10780 22204 10836
rect 22260 10780 23996 10836
rect 24052 10780 24062 10836
rect 24210 10780 24220 10836
rect 24276 10780 30156 10836
rect 30212 10780 30222 10836
rect 5842 10668 5852 10724
rect 5908 10668 8764 10724
rect 8820 10668 8830 10724
rect 13682 10668 13692 10724
rect 13748 10668 15260 10724
rect 15316 10668 15326 10724
rect 19730 10668 19740 10724
rect 19796 10668 20524 10724
rect 20580 10668 22316 10724
rect 22372 10668 22382 10724
rect 2258 10556 2268 10612
rect 2324 10556 4844 10612
rect 4900 10556 4910 10612
rect 6300 10388 6356 10668
rect 6514 10556 6524 10612
rect 6580 10556 6972 10612
rect 7028 10556 7038 10612
rect 17602 10556 17612 10612
rect 17668 10556 19404 10612
rect 19460 10556 19470 10612
rect 21858 10556 21868 10612
rect 21924 10556 23100 10612
rect 23156 10556 23166 10612
rect 15474 10444 15484 10500
rect 15540 10444 20748 10500
rect 20804 10444 21644 10500
rect 21700 10444 21710 10500
rect 22978 10444 22988 10500
rect 23044 10444 29148 10500
rect 29204 10444 29214 10500
rect 6300 10332 6524 10388
rect 6580 10332 6590 10388
rect 21942 10220 21980 10276
rect 22036 10220 22046 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19170 10108 19180 10164
rect 19236 10108 20132 10164
rect 20076 10052 20132 10108
rect 20076 9996 22652 10052
rect 22708 9996 22718 10052
rect 23314 9996 23324 10052
rect 23380 9996 25340 10052
rect 25396 9996 27244 10052
rect 27300 9996 27310 10052
rect 2258 9884 2268 9940
rect 2324 9884 4284 9940
rect 4340 9884 4350 9940
rect 6962 9884 6972 9940
rect 7028 9884 7420 9940
rect 7476 9884 8092 9940
rect 8148 9884 9548 9940
rect 9604 9884 9614 9940
rect 13010 9884 13020 9940
rect 13076 9884 13580 9940
rect 13636 9884 18508 9940
rect 18564 9884 18574 9940
rect 21980 9884 25116 9940
rect 25172 9884 25182 9940
rect 29698 9884 29708 9940
rect 29764 9884 30604 9940
rect 30660 9884 30670 9940
rect 7746 9772 7756 9828
rect 7812 9772 15148 9828
rect 15204 9772 15214 9828
rect 0 9716 800 9744
rect 21980 9716 22036 9884
rect 23202 9772 23212 9828
rect 23268 9772 29260 9828
rect 29316 9772 29326 9828
rect 28140 9716 28196 9772
rect 0 9660 1708 9716
rect 1764 9660 1774 9716
rect 20934 9660 20972 9716
rect 21028 9660 21038 9716
rect 21410 9660 21420 9716
rect 21476 9660 21868 9716
rect 21924 9660 22036 9716
rect 22754 9660 22764 9716
rect 22820 9660 23996 9716
rect 24052 9660 24062 9716
rect 28130 9660 28140 9716
rect 28196 9660 28206 9716
rect 0 9632 800 9660
rect 5954 9548 5964 9604
rect 6020 9548 6412 9604
rect 6468 9548 6478 9604
rect 9986 9548 9996 9604
rect 10052 9548 15708 9604
rect 15764 9548 15774 9604
rect 19730 9548 19740 9604
rect 19796 9548 20636 9604
rect 20692 9548 24332 9604
rect 24388 9548 24398 9604
rect 29586 9548 29596 9604
rect 29652 9548 30268 9604
rect 30324 9548 31388 9604
rect 31444 9548 31454 9604
rect 11778 9436 11788 9492
rect 11844 9436 13356 9492
rect 13412 9436 13422 9492
rect 20738 9436 20748 9492
rect 20804 9436 21196 9492
rect 21252 9436 21262 9492
rect 22306 9436 22316 9492
rect 22372 9436 23100 9492
rect 23156 9436 23166 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 2034 9324 2044 9380
rect 2100 9324 14700 9380
rect 14756 9324 15820 9380
rect 15876 9324 15886 9380
rect 20850 9324 20860 9380
rect 20916 9324 21308 9380
rect 21364 9324 21374 9380
rect 15362 9212 15372 9268
rect 15428 9212 16156 9268
rect 16212 9212 16222 9268
rect 22642 9212 22652 9268
rect 22708 9212 23996 9268
rect 24052 9212 24062 9268
rect 14690 9100 14700 9156
rect 14756 9100 15148 9156
rect 15810 9100 15820 9156
rect 15876 9100 16716 9156
rect 16772 9100 16782 9156
rect 22418 9100 22428 9156
rect 22484 9100 23436 9156
rect 23492 9100 23502 9156
rect 15092 9044 15148 9100
rect 15092 8988 21196 9044
rect 21252 8988 29596 9044
rect 29652 8988 29662 9044
rect 15026 8876 15036 8932
rect 15092 8876 21420 8932
rect 21476 8876 21486 8932
rect 23090 8876 23100 8932
rect 23156 8876 26012 8932
rect 26068 8876 26078 8932
rect 10546 8764 10556 8820
rect 10612 8764 12012 8820
rect 12068 8764 22092 8820
rect 22148 8764 22988 8820
rect 23044 8764 23054 8820
rect 10892 8652 11116 8708
rect 11172 8652 11182 8708
rect 15810 8652 15820 8708
rect 15876 8652 16716 8708
rect 16772 8652 17276 8708
rect 17332 8652 20748 8708
rect 20804 8652 20814 8708
rect 20962 8652 20972 8708
rect 21028 8652 21980 8708
rect 22036 8652 22046 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 0 8372 800 8400
rect 10892 8372 10948 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 18498 8540 18508 8596
rect 18564 8540 19180 8596
rect 19236 8540 19246 8596
rect 12684 8428 14420 8484
rect 19058 8428 19068 8484
rect 19124 8428 19516 8484
rect 19572 8428 19582 8484
rect 12684 8372 12740 8428
rect 14364 8372 14420 8428
rect 0 8316 1708 8372
rect 1764 8316 2492 8372
rect 2548 8316 2558 8372
rect 9874 8316 9884 8372
rect 9940 8316 10668 8372
rect 10724 8316 10734 8372
rect 10892 8316 12740 8372
rect 13010 8316 13020 8372
rect 13076 8316 13356 8372
rect 13412 8316 14140 8372
rect 14196 8316 14206 8372
rect 14364 8316 16268 8372
rect 16324 8316 16334 8372
rect 16594 8316 16604 8372
rect 16660 8316 18732 8372
rect 18788 8316 19292 8372
rect 19348 8316 19852 8372
rect 19908 8316 19918 8372
rect 20514 8316 20524 8372
rect 20580 8316 21644 8372
rect 21700 8316 22316 8372
rect 22372 8316 22382 8372
rect 22530 8316 22540 8372
rect 22596 8316 23548 8372
rect 23604 8316 26124 8372
rect 26180 8316 26190 8372
rect 0 8288 800 8316
rect 16268 8260 16324 8316
rect 10770 8204 10780 8260
rect 10836 8204 11564 8260
rect 11620 8204 12908 8260
rect 12964 8204 13468 8260
rect 13524 8204 13534 8260
rect 16268 8204 18508 8260
rect 18564 8204 19964 8260
rect 20020 8204 20030 8260
rect 20178 8204 20188 8260
rect 20244 8204 21756 8260
rect 21812 8204 21822 8260
rect 19964 8148 20020 8204
rect 9426 8092 9436 8148
rect 9492 8092 12348 8148
rect 12404 8092 12414 8148
rect 12786 8092 12796 8148
rect 12852 8092 14364 8148
rect 14420 8092 15036 8148
rect 15092 8092 15102 8148
rect 15922 8092 15932 8148
rect 15988 8092 16604 8148
rect 16660 8092 16828 8148
rect 16884 8092 16894 8148
rect 19964 8092 20356 8148
rect 20738 8092 20748 8148
rect 20804 8092 21868 8148
rect 21924 8092 22204 8148
rect 22260 8092 22270 8148
rect 12348 8036 12404 8092
rect 20300 8036 20356 8092
rect 7858 7980 7868 8036
rect 7924 7980 9884 8036
rect 9940 7980 9950 8036
rect 10322 7980 10332 8036
rect 10388 7980 11004 8036
rect 11060 7980 12012 8036
rect 12068 7980 12078 8036
rect 12348 7980 13580 8036
rect 13636 7980 15484 8036
rect 15540 7980 15550 8036
rect 16930 7980 16940 8036
rect 16996 7980 18620 8036
rect 18676 7980 18686 8036
rect 19506 7980 19516 8036
rect 19572 7980 19964 8036
rect 20020 7980 20030 8036
rect 20300 7980 22876 8036
rect 22932 7980 22942 8036
rect 10770 7868 10780 7924
rect 10836 7868 10948 7924
rect 10892 7812 10948 7868
rect 14700 7868 17388 7924
rect 17444 7868 19572 7924
rect 14700 7812 14756 7868
rect 10892 7756 14756 7812
rect 17826 7756 17836 7812
rect 17892 7756 19292 7812
rect 19348 7756 19358 7812
rect 19516 7700 19572 7868
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 9762 7644 9772 7700
rect 9828 7644 10220 7700
rect 10276 7644 10286 7700
rect 10434 7644 10444 7700
rect 10500 7644 11788 7700
rect 11844 7644 11854 7700
rect 15362 7644 15372 7700
rect 15428 7644 15820 7700
rect 15876 7644 18172 7700
rect 18228 7644 18238 7700
rect 18386 7644 18396 7700
rect 18452 7644 18956 7700
rect 19012 7644 19022 7700
rect 19516 7644 20300 7700
rect 20356 7644 20366 7700
rect 21410 7644 21420 7700
rect 21476 7644 21756 7700
rect 21812 7644 21822 7700
rect 10444 7476 10500 7644
rect 17154 7532 17164 7588
rect 17220 7532 17724 7588
rect 17780 7532 17790 7588
rect 19954 7532 19964 7588
rect 20020 7532 20636 7588
rect 20692 7532 21980 7588
rect 22036 7532 35084 7588
rect 35140 7532 35150 7588
rect 9986 7420 9996 7476
rect 10052 7420 10500 7476
rect 14130 7420 14140 7476
rect 14196 7420 16828 7476
rect 16884 7420 16894 7476
rect 10994 7308 11004 7364
rect 11060 7308 11508 7364
rect 11666 7308 11676 7364
rect 11732 7308 12460 7364
rect 12516 7308 12526 7364
rect 16594 7308 16604 7364
rect 16660 7308 18956 7364
rect 19012 7308 19022 7364
rect 11452 7252 11508 7308
rect 11442 7196 11452 7252
rect 11508 7196 19516 7252
rect 19572 7196 19582 7252
rect 13346 7084 13356 7140
rect 13412 7084 13916 7140
rect 13972 7084 13982 7140
rect 0 7028 800 7056
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 0 6972 1708 7028
rect 1764 6972 2492 7028
rect 2548 6972 2558 7028
rect 0 6944 800 6972
rect 11890 6860 11900 6916
rect 11956 6860 13244 6916
rect 13300 6860 13310 6916
rect 17938 6748 17948 6804
rect 18004 6748 18284 6804
rect 18340 6748 18350 6804
rect 7074 6636 7084 6692
rect 7140 6636 8092 6692
rect 8148 6636 10220 6692
rect 10276 6636 10286 6692
rect 11442 6636 11452 6692
rect 11508 6636 12684 6692
rect 12740 6636 12750 6692
rect 15138 6636 15148 6692
rect 15204 6636 17836 6692
rect 17892 6636 18844 6692
rect 18900 6636 21308 6692
rect 21364 6636 21374 6692
rect 37762 6636 37772 6692
rect 37828 6636 42812 6692
rect 42868 6636 42878 6692
rect 12786 6524 12796 6580
rect 12852 6524 13692 6580
rect 13748 6524 13758 6580
rect 8866 6412 8876 6468
rect 8932 6412 10668 6468
rect 10724 6412 10734 6468
rect 11330 6412 11340 6468
rect 11396 6412 11900 6468
rect 11956 6412 11966 6468
rect 13794 6412 13804 6468
rect 13860 6412 15596 6468
rect 15652 6412 15662 6468
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 2146 6076 2156 6132
rect 2212 6076 3276 6132
rect 3332 6076 3342 6132
rect 10210 5852 10220 5908
rect 10276 5852 10556 5908
rect 10612 5852 10892 5908
rect 10948 5852 10958 5908
rect 0 5684 800 5712
rect 0 5628 1708 5684
rect 1764 5628 2492 5684
rect 2548 5628 2558 5684
rect 17042 5628 17052 5684
rect 17108 5628 18396 5684
rect 18452 5628 18462 5684
rect 0 5600 800 5628
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 10210 5180 10220 5236
rect 10276 5180 11004 5236
rect 11060 5180 11070 5236
rect 11778 5180 11788 5236
rect 11844 5180 12684 5236
rect 12740 5180 24220 5236
rect 24276 5180 24286 5236
rect 16370 5068 16380 5124
rect 16436 5068 17500 5124
rect 17556 5068 17566 5124
rect 42578 5068 42588 5124
rect 42644 5068 43148 5124
rect 43204 5068 43214 5124
rect 1698 4844 1708 4900
rect 1764 4844 2492 4900
rect 2548 4844 2558 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 44200 4564 45000 4592
rect 8372 4508 10108 4564
rect 10164 4508 10174 4564
rect 23492 4508 23884 4564
rect 23940 4508 23950 4564
rect 43138 4508 43148 4564
rect 43204 4508 45000 4564
rect 0 4340 800 4368
rect 8372 4340 8428 4508
rect 23492 4340 23548 4508
rect 44200 4480 45000 4508
rect 0 4284 1708 4340
rect 1764 4284 1774 4340
rect 6066 4284 6076 4340
rect 6132 4284 8428 4340
rect 20962 4284 20972 4340
rect 21028 4284 22988 4340
rect 23044 4284 23548 4340
rect 28802 4284 28812 4340
rect 28868 4284 30380 4340
rect 30436 4284 30446 4340
rect 35074 4284 35084 4340
rect 35140 4284 42812 4340
rect 42868 4284 42878 4340
rect 0 4256 800 4284
rect 6290 4060 6300 4116
rect 6356 4060 7420 4116
rect 7476 4060 7486 4116
rect 13458 4060 13468 4116
rect 13524 4060 14700 4116
rect 14756 4060 14766 4116
rect 29586 4060 29596 4116
rect 29652 4060 30828 4116
rect 30884 4060 30894 4116
rect 36754 4060 36764 4116
rect 36820 4060 37996 4116
rect 38052 4060 38062 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 27794 3612 27804 3668
rect 27860 3612 29372 3668
rect 29428 3612 29438 3668
rect 34962 3612 34972 3668
rect 35028 3612 36988 3668
rect 37044 3612 37054 3668
rect 38546 3612 38556 3668
rect 38612 3612 40796 3668
rect 40852 3612 40862 3668
rect 8754 3500 8764 3556
rect 8820 3500 14028 3556
rect 14084 3500 14094 3556
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 0 2996 800 3024
rect 0 2940 1820 2996
rect 1876 2940 1886 2996
rect 0 2912 800 2940
<< via3 >>
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 8204 37884 8260 37940
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 7756 36876 7812 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 8092 36764 8148 36820
rect 6972 36316 7028 36372
rect 8204 36316 8260 36372
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 7756 35868 7812 35924
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 11340 33740 11396 33796
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 17388 32508 17444 32564
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 8092 31612 8148 31668
rect 11452 31500 11508 31556
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 11004 30604 11060 30660
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 16156 30268 16212 30324
rect 17724 30268 17780 30324
rect 11452 30044 11508 30100
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 16156 29708 16212 29764
rect 16604 29372 16660 29428
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 11340 28812 11396 28868
rect 27356 28700 27412 28756
rect 15820 28588 15876 28644
rect 16268 28476 16324 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 27356 28140 27412 28196
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 11452 27132 11508 27188
rect 11004 27020 11060 27076
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 16268 26460 16324 26516
rect 15820 26348 15876 26404
rect 16604 26124 16660 26180
rect 11452 25900 11508 25956
rect 17388 25900 17444 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 33852 25788 33908 25844
rect 17724 25228 17780 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 15036 24892 15092 24948
rect 15148 24444 15204 24500
rect 10108 24332 10164 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 33852 23436 33908 23492
rect 13244 23100 13300 23156
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 5852 22540 5908 22596
rect 10108 22316 10164 22372
rect 11228 22092 11284 22148
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 17388 21868 17444 21924
rect 15708 21756 15764 21812
rect 16828 21420 16884 21476
rect 22316 21308 22372 21364
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 17388 21084 17444 21140
rect 15820 20860 15876 20916
rect 21868 20860 21924 20916
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 22428 19292 22484 19348
rect 13580 19068 13636 19124
rect 22316 18844 22372 18900
rect 13244 18732 13300 18788
rect 18732 18732 18788 18788
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 21868 17724 21924 17780
rect 13580 17388 13636 17444
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 14700 16828 14756 16884
rect 22428 16828 22484 16884
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 17612 16380 17668 16436
rect 10108 16268 10164 16324
rect 18732 15708 18788 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 16828 15372 16884 15428
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 11228 14588 11284 14644
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 6972 13020 7028 13076
rect 5852 12796 5908 12852
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 17612 12460 17668 12516
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 17276 11116 17332 11172
rect 22092 11116 22148 11172
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 21980 10220 22036 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 20972 9660 21028 9716
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 14700 9100 14756 9156
rect 22092 8764 22148 8820
rect 17276 8652 17332 8708
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 21980 7532 22036 7588
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 20972 4284 21028 4340
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 41580 4768 41612
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 19808 40796 20128 41612
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 8204 37940 8260 37950
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 7756 36932 7812 36942
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 6972 36372 7028 36382
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 5852 22596 5908 22606
rect 5852 12852 5908 22540
rect 6972 13076 7028 36316
rect 7756 35924 7812 36876
rect 7756 35858 7812 35868
rect 8092 36820 8148 36830
rect 8092 31668 8148 36764
rect 8204 36372 8260 37884
rect 8204 36306 8260 36316
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 8092 31602 8148 31612
rect 11340 33796 11396 33806
rect 11004 30660 11060 30670
rect 11004 27076 11060 30604
rect 11340 28868 11396 33740
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 17388 32564 17444 32574
rect 11452 31556 11508 31566
rect 11452 30100 11508 31500
rect 11452 30034 11508 30044
rect 16156 30324 16212 30334
rect 16156 29764 16212 30268
rect 16156 29698 16212 29708
rect 11340 28802 11396 28812
rect 16604 29428 16660 29438
rect 15820 28644 15876 28654
rect 11004 27010 11060 27020
rect 11452 27188 11508 27198
rect 11452 25956 11508 27132
rect 15820 26404 15876 28588
rect 16268 28532 16324 28542
rect 16268 26516 16324 28476
rect 16268 26450 16324 26460
rect 15820 26338 15876 26348
rect 16604 26180 16660 29372
rect 16604 26114 16660 26124
rect 11452 25890 11508 25900
rect 17388 25956 17444 32508
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 17388 25890 17444 25900
rect 17724 30324 17780 30334
rect 17724 25284 17780 30268
rect 17724 25218 17780 25228
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 35168 41580 35488 41612
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 27356 28756 27412 28766
rect 27356 28196 27412 28700
rect 27356 28130 27412 28140
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 15036 24948 15204 24958
rect 15092 24902 15204 24948
rect 15036 24882 15092 24892
rect 15148 24500 15204 24902
rect 15148 24434 15204 24444
rect 10108 24388 10164 24398
rect 10108 22372 10164 24332
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 10108 16324 10164 22316
rect 13244 23156 13300 23166
rect 10108 16258 10164 16268
rect 11228 22148 11284 22158
rect 11228 14644 11284 22092
rect 13244 18788 13300 23100
rect 19808 21980 20128 23492
rect 33852 25844 33908 25854
rect 33852 23492 33908 25788
rect 33852 23426 33908 23436
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 17388 21924 17444 21934
rect 15708 21812 15764 21822
rect 15708 20998 15764 21756
rect 16828 21476 16884 21486
rect 15708 20942 15876 20998
rect 15820 20916 15876 20942
rect 15820 20850 15876 20860
rect 13244 18722 13300 18732
rect 13580 19124 13636 19134
rect 13580 17444 13636 19068
rect 13580 17378 13636 17388
rect 11228 14578 11284 14588
rect 14700 16884 14756 16894
rect 6972 13010 7028 13020
rect 5852 12786 5908 12796
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 14700 9156 14756 16828
rect 16828 15428 16884 21420
rect 17388 21140 17444 21868
rect 17388 21074 17444 21084
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 22316 21364 22372 21374
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 18732 18788 18788 18798
rect 16828 15362 16884 15372
rect 17612 16436 17668 16446
rect 17612 12516 17668 16380
rect 18732 15764 18788 18732
rect 18732 15698 18788 15708
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 21868 20916 21924 20926
rect 21868 17780 21924 20860
rect 22316 18900 22372 21308
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 22316 18834 22372 18844
rect 22428 19348 22484 19358
rect 21868 17714 21924 17724
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 22428 16884 22484 19292
rect 22428 16818 22484 16828
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 17612 12450 17668 12460
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 14700 9090 14756 9100
rect 17276 11172 17332 11182
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 17276 8708 17332 11116
rect 17276 8642 17332 8652
rect 19808 11004 20128 12516
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 22092 11172 22148 11182
rect 21980 10276 22036 10286
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 20972 9716 21028 9726
rect 20972 4340 21028 9660
rect 21980 7588 22036 10220
rect 22092 8820 22148 11116
rect 22092 8754 22148 8764
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 21980 7522 22036 7532
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 20972 4274 21028 4284
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _397_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _398_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15120 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _399_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19936 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _400_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _401_
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _402_
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _403_
timestamp 1698431365
transform 1 0 16128 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _404_
timestamp 1698431365
transform 1 0 22288 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _405_
timestamp 1698431365
transform -1 0 25872 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _406_
timestamp 1698431365
transform 1 0 24192 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _407_
timestamp 1698431365
transform 1 0 28000 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _408_
timestamp 1698431365
transform 1 0 26992 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _409_
timestamp 1698431365
transform 1 0 27104 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _410_
timestamp 1698431365
transform 1 0 27440 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _411_
timestamp 1698431365
transform 1 0 30576 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _412_
timestamp 1698431365
transform 1 0 30352 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _413_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _414_
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _415_
timestamp 1698431365
transform 1 0 27664 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _416_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11648 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _417_
timestamp 1698431365
transform -1 0 14448 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _418_
timestamp 1698431365
transform 1 0 11200 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _419_
timestamp 1698431365
transform -1 0 14672 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _420_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _421_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6496 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _422_
timestamp 1698431365
transform 1 0 3584 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _423_
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _424_
timestamp 1698431365
transform 1 0 21952 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _425_
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _426_
timestamp 1698431365
transform -1 0 30352 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _427_
timestamp 1698431365
transform 1 0 31024 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _428_
timestamp 1698431365
transform 1 0 23184 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _429_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _430_
timestamp 1698431365
transform 1 0 31696 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _431_
timestamp 1698431365
transform 1 0 22960 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _432_
timestamp 1698431365
transform 1 0 24416 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _433_
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _434_
timestamp 1698431365
transform 1 0 26880 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _435_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _436_
timestamp 1698431365
transform 1 0 31024 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _437_
timestamp 1698431365
transform 1 0 29008 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _438_
timestamp 1698431365
transform 1 0 31136 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _439_
timestamp 1698431365
transform 1 0 34832 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _440_
timestamp 1698431365
transform 1 0 31472 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _441_
timestamp 1698431365
transform 1 0 34048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _442_
timestamp 1698431365
transform 1 0 35840 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _443_
timestamp 1698431365
transform 1 0 32592 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _444_
timestamp 1698431365
transform 1 0 34272 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _445_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _446_
timestamp 1698431365
transform 1 0 18256 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _447_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6048 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _448_
timestamp 1698431365
transform 1 0 6048 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _449_
timestamp 1698431365
transform 1 0 15120 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _450_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18592 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _451_
timestamp 1698431365
transform -1 0 22176 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _452_
timestamp 1698431365
transform 1 0 21952 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _453_
timestamp 1698431365
transform -1 0 26096 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _454_
timestamp 1698431365
transform -1 0 28112 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _455_
timestamp 1698431365
transform 1 0 28000 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _456_
timestamp 1698431365
transform 1 0 29456 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _457_
timestamp 1698431365
transform 1 0 25872 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _458_
timestamp 1698431365
transform 1 0 38192 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _459_
timestamp 1698431365
transform 1 0 23968 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _460_
timestamp 1698431365
transform 1 0 38976 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _461_
timestamp 1698431365
transform -1 0 19824 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _462_
timestamp 1698431365
transform -1 0 18144 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _463_
timestamp 1698431365
transform 1 0 29568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _464_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _465_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35280 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _466_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _467_
timestamp 1698431365
transform -1 0 15008 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _468_
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _469_
timestamp 1698431365
transform 1 0 11088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _470_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1792 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _471_
timestamp 1698431365
transform 1 0 2912 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _472_
timestamp 1698431365
transform 1 0 2912 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _473_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3696 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _474_
timestamp 1698431365
transform 1 0 2800 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _475_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15344 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _476_
timestamp 1698431365
transform -1 0 2352 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _477_
timestamp 1698431365
transform 1 0 5712 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _478_
timestamp 1698431365
transform 1 0 3360 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _479_
timestamp 1698431365
transform -1 0 2800 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _480_
timestamp 1698431365
transform 1 0 3808 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _481_
timestamp 1698431365
transform -1 0 2800 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _482_
timestamp 1698431365
transform 1 0 1680 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _483_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6160 0 1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _484_
timestamp 1698431365
transform 1 0 15792 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _485_
timestamp 1698431365
transform 1 0 3472 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _486_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6048 0 -1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _487_
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _488_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14448 0 1 20384
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _489_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _490_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10976 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _491_
timestamp 1698431365
transform 1 0 10640 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _492_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5264 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _493_
timestamp 1698431365
transform 1 0 16464 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _494_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15680 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _495_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6160 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _496_
timestamp 1698431365
transform -1 0 8848 0 -1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _497_
timestamp 1698431365
transform 1 0 6384 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _498_
timestamp 1698431365
transform 1 0 4368 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _499_
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _500_
timestamp 1698431365
transform 1 0 15120 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _501_
timestamp 1698431365
transform -1 0 7952 0 -1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _502_
timestamp 1698431365
transform -1 0 11088 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _503_
timestamp 1698431365
transform -1 0 12880 0 -1 32928
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _504_
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _505_
timestamp 1698431365
transform 1 0 16016 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _506_
timestamp 1698431365
transform 1 0 4368 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _507_
timestamp 1698431365
transform 1 0 11200 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _508_
timestamp 1698431365
transform 1 0 15344 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _509_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11536 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _510_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12880 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _511_
timestamp 1698431365
transform -1 0 18816 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _512_
timestamp 1698431365
transform -1 0 11760 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _513_
timestamp 1698431365
transform 1 0 4928 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _514_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4368 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _515_
timestamp 1698431365
transform 1 0 11312 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _516_
timestamp 1698431365
transform 1 0 10976 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _517_
timestamp 1698431365
transform -1 0 11200 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _518_
timestamp 1698431365
transform 1 0 14672 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _519_
timestamp 1698431365
transform -1 0 14224 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _520_
timestamp 1698431365
transform -1 0 14896 0 -1 36064
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _521_
timestamp 1698431365
transform -1 0 8288 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _522_
timestamp 1698431365
transform 1 0 7280 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _523_
timestamp 1698431365
transform -1 0 17248 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _524_
timestamp 1698431365
transform -1 0 18256 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _525_
timestamp 1698431365
transform 1 0 9744 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _526_
timestamp 1698431365
transform -1 0 11088 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _527_
timestamp 1698431365
transform 1 0 8176 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _528_
timestamp 1698431365
transform -1 0 17024 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _529_
timestamp 1698431365
transform 1 0 9520 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _530_
timestamp 1698431365
transform -1 0 11872 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _531_
timestamp 1698431365
transform 1 0 5712 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _532_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10416 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _533_
timestamp 1698431365
transform 1 0 11200 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _534_
timestamp 1698431365
transform -1 0 10528 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _535_
timestamp 1698431365
transform -1 0 17360 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _536_
timestamp 1698431365
transform -1 0 10976 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _537_
timestamp 1698431365
transform -1 0 8064 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _538_
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _539_
timestamp 1698431365
transform 1 0 12768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _540_
timestamp 1698431365
transform 1 0 13664 0 -1 17248
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _541_
timestamp 1698431365
transform 1 0 14224 0 -1 32928
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _542_
timestamp 1698431365
transform 1 0 15792 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _543_
timestamp 1698431365
transform 1 0 8176 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _544_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6720 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _545_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7952 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _546_
timestamp 1698431365
transform -1 0 7840 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _547_
timestamp 1698431365
transform 1 0 5600 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _548_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _549_
timestamp 1698431365
transform 1 0 12096 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _550_
timestamp 1698431365
transform -1 0 11312 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _551_
timestamp 1698431365
transform -1 0 12432 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _552_
timestamp 1698431365
transform 1 0 15344 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _553_
timestamp 1698431365
transform -1 0 12432 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _554_
timestamp 1698431365
transform -1 0 8176 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _555_
timestamp 1698431365
transform 1 0 6608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _556_
timestamp 1698431365
transform 1 0 13664 0 1 15680
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _557_
timestamp 1698431365
transform 1 0 14000 0 1 32928
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _558_
timestamp 1698431365
transform 1 0 9408 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _559_
timestamp 1698431365
transform -1 0 7616 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _560_
timestamp 1698431365
transform -1 0 8176 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _561_
timestamp 1698431365
transform -1 0 8176 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _562_
timestamp 1698431365
transform -1 0 12656 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _563_
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _564_
timestamp 1698431365
transform -1 0 14896 0 -1 37632
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _565_
timestamp 1698431365
transform -1 0 17360 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _566_
timestamp 1698431365
transform -1 0 17024 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _567_
timestamp 1698431365
transform -1 0 16128 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _568_
timestamp 1698431365
transform -1 0 12208 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _569_
timestamp 1698431365
transform 1 0 10192 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _570_
timestamp 1698431365
transform -1 0 19824 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _571_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5600 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _572_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _573_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11984 0 -1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _574_
timestamp 1698431365
transform -1 0 10416 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _575_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _576_
timestamp 1698431365
transform 1 0 16576 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _577_
timestamp 1698431365
transform -1 0 14448 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _578_
timestamp 1698431365
transform -1 0 11984 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _579_
timestamp 1698431365
transform 1 0 15680 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _580_
timestamp 1698431365
transform 1 0 15456 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _581_
timestamp 1698431365
transform 1 0 16352 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _582_
timestamp 1698431365
transform -1 0 17136 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _583_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29680 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _584_
timestamp 1698431365
transform 1 0 14784 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _585_
timestamp 1698431365
transform 1 0 32032 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _586_
timestamp 1698431365
transform 1 0 31360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _587_
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _588_
timestamp 1698431365
transform 1 0 27440 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _589_
timestamp 1698431365
transform 1 0 29232 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _590_
timestamp 1698431365
transform 1 0 17360 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _591_
timestamp 1698431365
transform 1 0 34496 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _592_
timestamp 1698431365
transform 1 0 33488 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _593_
timestamp 1698431365
transform -1 0 33600 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _594_
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _595_
timestamp 1698431365
transform 1 0 9856 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _596_
timestamp 1698431365
transform 1 0 29680 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _597_
timestamp 1698431365
transform -1 0 36624 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _598_
timestamp 1698431365
transform 1 0 33824 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _599_
timestamp 1698431365
transform 1 0 35280 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _600_
timestamp 1698431365
transform 1 0 14560 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _601_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3696 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _602_
timestamp 1698431365
transform -1 0 15008 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _603_
timestamp 1698431365
transform -1 0 8960 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _604_
timestamp 1698431365
transform 1 0 8288 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _605_
timestamp 1698431365
transform -1 0 7392 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _606_
timestamp 1698431365
transform -1 0 16128 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _607_
timestamp 1698431365
transform -1 0 6384 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _608_
timestamp 1698431365
transform -1 0 4704 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _609_
timestamp 1698431365
transform -1 0 3584 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _610_
timestamp 1698431365
transform 1 0 4480 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _611_
timestamp 1698431365
transform -1 0 10752 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _612_
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _613_
timestamp 1698431365
transform 1 0 2464 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _614_
timestamp 1698431365
transform -1 0 5152 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _615_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2912 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _616_
timestamp 1698431365
transform -1 0 7392 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _617_
timestamp 1698431365
transform -1 0 7056 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _618_
timestamp 1698431365
transform 1 0 4592 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _619_
timestamp 1698431365
transform 1 0 4816 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _620_
timestamp 1698431365
transform 1 0 5600 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _621_
timestamp 1698431365
transform -1 0 4928 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _622_
timestamp 1698431365
transform -1 0 2912 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _623_
timestamp 1698431365
transform 1 0 21392 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _624_
timestamp 1698431365
transform -1 0 21168 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _625_
timestamp 1698431365
transform 1 0 1904 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _626_
timestamp 1698431365
transform 1 0 10192 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _627_
timestamp 1698431365
transform 1 0 9296 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _628_
timestamp 1698431365
transform 1 0 8176 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _629_
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _630_
timestamp 1698431365
transform 1 0 1904 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _631_
timestamp 1698431365
transform 1 0 4704 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _632_
timestamp 1698431365
transform 1 0 2352 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _633_
timestamp 1698431365
transform 1 0 22064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _634_
timestamp 1698431365
transform 1 0 10304 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _635_
timestamp 1698431365
transform 1 0 7168 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _636_
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _637_
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _638_
timestamp 1698431365
transform -1 0 8288 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _639_
timestamp 1698431365
transform -1 0 7952 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _640_
timestamp 1698431365
transform -1 0 20832 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _641_
timestamp 1698431365
transform -1 0 10304 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _642_
timestamp 1698431365
transform 1 0 7280 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _643_
timestamp 1698431365
transform -1 0 16800 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _644_
timestamp 1698431365
transform -1 0 12880 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _645_
timestamp 1698431365
transform 1 0 11424 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _646_
timestamp 1698431365
transform -1 0 7504 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _647_
timestamp 1698431365
transform -1 0 12096 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _648_
timestamp 1698431365
transform -1 0 11424 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _649_
timestamp 1698431365
transform -1 0 6720 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _650_
timestamp 1698431365
transform 1 0 6048 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _651_
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _652_
timestamp 1698431365
transform -1 0 10864 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _653_
timestamp 1698431365
transform 1 0 8624 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _654_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _655_
timestamp 1698431365
transform -1 0 7392 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _656_
timestamp 1698431365
transform -1 0 6048 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _657_
timestamp 1698431365
transform 1 0 5600 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _658_
timestamp 1698431365
transform 1 0 17920 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _659_
timestamp 1698431365
transform 1 0 12544 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _660_
timestamp 1698431365
transform 1 0 12096 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _661_
timestamp 1698431365
transform 1 0 10528 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _662_
timestamp 1698431365
transform -1 0 12544 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _663_
timestamp 1698431365
transform -1 0 11648 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _664_
timestamp 1698431365
transform -1 0 11760 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _665_
timestamp 1698431365
transform -1 0 11760 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _666_
timestamp 1698431365
transform -1 0 11648 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _667_
timestamp 1698431365
transform -1 0 11088 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _668_
timestamp 1698431365
transform 1 0 26208 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _669_
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _670_
timestamp 1698431365
transform 1 0 12768 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _671_
timestamp 1698431365
transform -1 0 12768 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _672_
timestamp 1698431365
transform -1 0 10864 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _673_
timestamp 1698431365
transform -1 0 10752 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _674_
timestamp 1698431365
transform 1 0 9632 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _675_
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _676_
timestamp 1698431365
transform 1 0 12544 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _677_
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _678_
timestamp 1698431365
transform 1 0 13440 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _679_
timestamp 1698431365
transform 1 0 6048 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _680_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _681_
timestamp 1698431365
transform 1 0 18256 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _682_
timestamp 1698431365
transform -1 0 16464 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _683_
timestamp 1698431365
transform 1 0 17024 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _684_
timestamp 1698431365
transform -1 0 17920 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _685_
timestamp 1698431365
transform -1 0 16128 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _686_
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _687_
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _688_
timestamp 1698431365
transform 1 0 17248 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _689_
timestamp 1698431365
transform -1 0 18368 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _690_
timestamp 1698431365
transform 1 0 16464 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _691_
timestamp 1698431365
transform 1 0 18816 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _692_
timestamp 1698431365
transform -1 0 17920 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _693_
timestamp 1698431365
transform -1 0 19488 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _694_
timestamp 1698431365
transform 1 0 16464 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _695_
timestamp 1698431365
transform -1 0 18816 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _696_
timestamp 1698431365
transform 1 0 19712 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _697_
timestamp 1698431365
transform 1 0 19264 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _698_
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _699_
timestamp 1698431365
transform 1 0 20272 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _700_
timestamp 1698431365
transform 1 0 21280 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _701_
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _702_
timestamp 1698431365
transform 1 0 22176 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _703_
timestamp 1698431365
transform -1 0 23072 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _704_
timestamp 1698431365
transform 1 0 22736 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _705_
timestamp 1698431365
transform 1 0 22176 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _706_
timestamp 1698431365
transform 1 0 22848 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _707_
timestamp 1698431365
transform 1 0 21392 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _708_
timestamp 1698431365
transform 1 0 21504 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _709_
timestamp 1698431365
transform 1 0 22736 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _710_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _711_
timestamp 1698431365
transform -1 0 18256 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _712_
timestamp 1698431365
transform -1 0 15680 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _713_
timestamp 1698431365
transform 1 0 15568 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _714_
timestamp 1698431365
transform -1 0 17024 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _715_
timestamp 1698431365
transform -1 0 14224 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _716_
timestamp 1698431365
transform -1 0 25872 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _717_
timestamp 1698431365
transform -1 0 20832 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _718_
timestamp 1698431365
transform 1 0 14224 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _719_
timestamp 1698431365
transform 1 0 17808 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _720_
timestamp 1698431365
transform 1 0 17136 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _721_
timestamp 1698431365
transform 1 0 17920 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _722_
timestamp 1698431365
transform 1 0 15008 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _723_
timestamp 1698431365
transform -1 0 16576 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _724_
timestamp 1698431365
transform -1 0 16128 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _725_
timestamp 1698431365
transform 1 0 18032 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _726_
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _727_
timestamp 1698431365
transform 1 0 18368 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _728_
timestamp 1698431365
transform 1 0 20048 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _729_
timestamp 1698431365
transform 1 0 22176 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _730_
timestamp 1698431365
transform 1 0 21056 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _731_
timestamp 1698431365
transform 1 0 22848 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _732_
timestamp 1698431365
transform -1 0 24864 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _733_
timestamp 1698431365
transform 1 0 23856 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _734_
timestamp 1698431365
transform 1 0 23632 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _735_
timestamp 1698431365
transform 1 0 23632 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _736_
timestamp 1698431365
transform -1 0 25984 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _737_
timestamp 1698431365
transform 1 0 22288 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _738_
timestamp 1698431365
transform 1 0 23408 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _739_
timestamp 1698431365
transform 1 0 23968 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _740_
timestamp 1698431365
transform 1 0 21728 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _741_
timestamp 1698431365
transform 1 0 22400 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _742_
timestamp 1698431365
transform 1 0 22960 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _743_
timestamp 1698431365
transform 1 0 17584 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _744_
timestamp 1698431365
transform -1 0 20832 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _745_
timestamp 1698431365
transform 1 0 20384 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _746_
timestamp 1698431365
transform 1 0 16464 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _747_
timestamp 1698431365
transform 1 0 20272 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _748_
timestamp 1698431365
transform 1 0 20384 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _749_
timestamp 1698431365
transform 1 0 21504 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _750_
timestamp 1698431365
transform 1 0 22736 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _751_
timestamp 1698431365
transform 1 0 20384 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _752_
timestamp 1698431365
transform 1 0 22176 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _753_
timestamp 1698431365
transform -1 0 22736 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _754_
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _755_
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _756_
timestamp 1698431365
transform 1 0 21504 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _757_
timestamp 1698431365
transform -1 0 20384 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _758_
timestamp 1698431365
transform -1 0 20608 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _759_
timestamp 1698431365
transform 1 0 20608 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _760_
timestamp 1698431365
transform 1 0 25872 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _761_
timestamp 1698431365
transform 1 0 27104 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _762_
timestamp 1698431365
transform 1 0 26096 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _763_
timestamp 1698431365
transform 1 0 27664 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _764_
timestamp 1698431365
transform 1 0 26656 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _765_
timestamp 1698431365
transform -1 0 28112 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _766_
timestamp 1698431365
transform 1 0 27440 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _767_
timestamp 1698431365
transform 1 0 27888 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _768_
timestamp 1698431365
transform 1 0 28448 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _769_
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _770_
timestamp 1698431365
transform 1 0 30576 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _771_
timestamp 1698431365
transform -1 0 30576 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _772_
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _773_
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _774_
timestamp 1698431365
transform 1 0 29680 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _775_
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _776_
timestamp 1698431365
transform -1 0 18480 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _777_
timestamp 1698431365
transform 1 0 18368 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _778_
timestamp 1698431365
transform -1 0 16576 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _779_
timestamp 1698431365
transform -1 0 16576 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _780_
timestamp 1698431365
transform 1 0 17584 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _781_
timestamp 1698431365
transform -1 0 26208 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _782_
timestamp 1698431365
transform -1 0 21840 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _783_
timestamp 1698431365
transform 1 0 19152 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _784_
timestamp 1698431365
transform -1 0 22624 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _785_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _786_
timestamp 1698431365
transform 1 0 19152 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _787_
timestamp 1698431365
transform -1 0 21168 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _788_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _789_
timestamp 1698431365
transform 1 0 22400 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _790_
timestamp 1698431365
transform 1 0 20048 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _791_
timestamp 1698431365
transform -1 0 24416 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _792_
timestamp 1698431365
transform -1 0 23856 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _793_
timestamp 1698431365
transform 1 0 25872 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _794_
timestamp 1698431365
transform 1 0 26208 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _795_
timestamp 1698431365
transform 1 0 27104 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _796_
timestamp 1698431365
transform 1 0 26432 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _797_
timestamp 1698431365
transform -1 0 28448 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _798_
timestamp 1698431365
transform -1 0 27888 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _799_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _800_
timestamp 1698431365
transform 1 0 28448 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _801_
timestamp 1698431365
transform 1 0 29568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _802_
timestamp 1698431365
transform 1 0 16576 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _803_
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _804_
timestamp 1698431365
transform 1 0 17360 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _805_
timestamp 1698431365
transform -1 0 24304 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _806_
timestamp 1698431365
transform -1 0 22512 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _807_
timestamp 1698431365
transform -1 0 23632 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _808_
timestamp 1698431365
transform -1 0 22288 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _809_
timestamp 1698431365
transform -1 0 24080 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _810_
timestamp 1698431365
transform -1 0 21840 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _811_
timestamp 1698431365
transform -1 0 22512 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _812_
timestamp 1698431365
transform 1 0 24304 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _813_
timestamp 1698431365
transform 1 0 22624 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _814_
timestamp 1698431365
transform 1 0 22512 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _815_
timestamp 1698431365
transform -1 0 24304 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _816_
timestamp 1698431365
transform 1 0 22512 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _817_
timestamp 1698431365
transform 1 0 27216 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _818_
timestamp 1698431365
transform 1 0 26544 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _819_
timestamp 1698431365
transform -1 0 28224 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _820_
timestamp 1698431365
transform -1 0 27552 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _821_
timestamp 1698431365
transform -1 0 28560 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _822_
timestamp 1698431365
transform -1 0 28112 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _823_
timestamp 1698431365
transform 1 0 28224 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _824_
timestamp 1698431365
transform -1 0 30016 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _825_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _826_
timestamp 1698431365
transform 1 0 30016 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _827_
timestamp 1698431365
transform -1 0 32032 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _828_
timestamp 1698431365
transform 1 0 33936 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _829_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33040 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _830_
timestamp 1698431365
transform -1 0 9184 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _831_
timestamp 1698431365
transform -1 0 4816 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _832_
timestamp 1698431365
transform -1 0 6720 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _833_
timestamp 1698431365
transform -1 0 4816 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _834_
timestamp 1698431365
transform -1 0 4816 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _835_
timestamp 1698431365
transform -1 0 6832 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _836_
timestamp 1698431365
transform -1 0 13104 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _837_
timestamp 1698431365
transform -1 0 9408 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _838_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31920 0 1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _839_
timestamp 1698431365
transform 1 0 33152 0 1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _840_
timestamp 1698431365
transform 1 0 35168 0 -1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _841_
timestamp 1698431365
transform -1 0 6720 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _842_
timestamp 1698431365
transform -1 0 5040 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _843_
timestamp 1698431365
transform 1 0 1680 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _844_
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _845_
timestamp 1698431365
transform -1 0 11536 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _846_
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _847_
timestamp 1698431365
transform 1 0 8512 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _848_
timestamp 1698431365
transform 1 0 4928 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _849_
timestamp 1698431365
transform 1 0 2016 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _850_
timestamp 1698431365
transform 1 0 7392 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _851_
timestamp 1698431365
transform 1 0 2016 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _852_
timestamp 1698431365
transform 1 0 10976 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _853_
timestamp 1698431365
transform 1 0 7952 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _854_
timestamp 1698431365
transform 1 0 10752 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _855_
timestamp 1698431365
transform 1 0 6944 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _856_
timestamp 1698431365
transform -1 0 16576 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _857_
timestamp 1698431365
transform 1 0 14896 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _858_
timestamp 1698431365
transform -1 0 19040 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _859_
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _860_
timestamp 1698431365
transform 1 0 17696 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _861_
timestamp 1698431365
transform 1 0 21168 0 -1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _862_
timestamp 1698431365
transform 1 0 23072 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _863_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _864_
timestamp 1698431365
transform 1 0 28336 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _865_
timestamp 1698431365
transform -1 0 15232 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _866_
timestamp 1698431365
transform 1 0 17584 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _867_
timestamp 1698431365
transform -1 0 16576 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _868_
timestamp 1698431365
transform 1 0 17696 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _869_
timestamp 1698431365
transform 1 0 25536 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _870_
timestamp 1698431365
transform 1 0 25424 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _871_
timestamp 1698431365
transform 1 0 28672 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _872_
timestamp 1698431365
transform 1 0 22736 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _873_
timestamp 1698431365
transform -1 0 22736 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _874_
timestamp 1698431365
transform 1 0 23408 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _875_
timestamp 1698431365
transform 1 0 21728 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _876_
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _877_
timestamp 1698431365
transform -1 0 28784 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _878_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _879_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _880_
timestamp 1698431365
transform 1 0 31024 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _881_
timestamp 1698431365
transform 1 0 12544 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _882_
timestamp 1698431365
transform -1 0 22288 0 -1 14112
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _883_
timestamp 1698431365
transform -1 0 20048 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _884_
timestamp 1698431365
transform 1 0 22400 0 1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _885_
timestamp 1698431365
transform 1 0 26992 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _886_
timestamp 1698431365
transform 1 0 26768 0 -1 14112
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _887_
timestamp 1698431365
transform 1 0 29232 0 -1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _888_
timestamp 1698431365
transform -1 0 20496 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _889_
timestamp 1698431365
transform -1 0 22400 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _890_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _891_
timestamp 1698431365
transform 1 0 22512 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _892_
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _893_
timestamp 1698431365
transform -1 0 28672 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _894_
timestamp 1698431365
transform -1 0 31808 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _895_
timestamp 1698431365
transform 1 0 29232 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _896_
timestamp 1698431365
transform 1 0 30576 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _897_
timestamp 1698431365
transform 1 0 30688 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _898_
timestamp 1698431365
transform 1 0 33600 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A1 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__I1
timestamp 1698431365
transform -1 0 18816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__S
timestamp 1698431365
transform 1 0 19040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__A1
timestamp 1698431365
transform -1 0 17696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__I1
timestamp 1698431365
transform 1 0 26544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__S
timestamp 1698431365
transform 1 0 26096 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__I0
timestamp 1698431365
transform 1 0 29904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__I1
timestamp 1698431365
transform 1 0 30128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__S
timestamp 1698431365
transform 1 0 30352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__I1
timestamp 1698431365
transform 1 0 29232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__S
timestamp 1698431365
transform 1 0 26880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__I0
timestamp 1698431365
transform 1 0 32480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__S
timestamp 1698431365
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__I
timestamp 1698431365
transform 1 0 18592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__A1
timestamp 1698431365
transform -1 0 23968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__A1
timestamp 1698431365
transform 1 0 11872 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__A1
timestamp 1698431365
transform 1 0 14672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__A1
timestamp 1698431365
transform -1 0 12768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__A2
timestamp 1698431365
transform -1 0 10192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A1
timestamp 1698431365
transform -1 0 15120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__A1
timestamp 1698431365
transform -1 0 14672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A1
timestamp 1698431365
transform 1 0 6720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A2
timestamp 1698431365
transform 1 0 5376 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__I
timestamp 1698431365
transform -1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__I0
timestamp 1698431365
transform -1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__S
timestamp 1698431365
transform 1 0 28336 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__I
timestamp 1698431365
transform 1 0 23856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__I
timestamp 1698431365
transform 1 0 31472 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__431__I
timestamp 1698431365
transform 1 0 23632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__A1
timestamp 1698431365
transform 1 0 24192 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__A2
timestamp 1698431365
transform 1 0 28784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__A1
timestamp 1698431365
transform -1 0 31136 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__A2
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__I
timestamp 1698431365
transform 1 0 32144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A1
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A2
timestamp 1698431365
transform 1 0 35168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__I
timestamp 1698431365
transform 1 0 33712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__A1
timestamp 1698431365
transform 1 0 34048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__A1
timestamp 1698431365
transform -1 0 19824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__A1
timestamp 1698431365
transform -1 0 5488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__A2
timestamp 1698431365
transform -1 0 5040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A1
timestamp 1698431365
transform -1 0 7840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A2
timestamp 1698431365
transform 1 0 5824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__A1
timestamp 1698431365
transform -1 0 15120 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__A2
timestamp 1698431365
transform 1 0 18816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__A2
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__A1
timestamp 1698431365
transform -1 0 24080 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__A2
timestamp 1698431365
transform 1 0 21168 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__453__A2
timestamp 1698431365
transform 1 0 25200 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__A1
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__A2
timestamp 1698431365
transform 1 0 26880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__A1
timestamp 1698431365
transform -1 0 28000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__A2
timestamp 1698431365
transform 1 0 29232 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__456__A1
timestamp 1698431365
transform 1 0 30688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__456__A2
timestamp 1698431365
transform 1 0 30240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A1
timestamp 1698431365
transform 1 0 26208 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A2
timestamp 1698431365
transform 1 0 26656 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__A1
timestamp 1698431365
transform 1 0 26208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__I
timestamp 1698431365
transform 1 0 20048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__I
timestamp 1698431365
transform 1 0 29344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A1
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A2
timestamp 1698431365
transform -1 0 12656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__A2
timestamp 1698431365
transform -1 0 34608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__I
timestamp 1698431365
transform 1 0 15232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__I
timestamp 1698431365
transform 1 0 15120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__B2
timestamp 1698431365
transform 1 0 17472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__C2
timestamp 1698431365
transform 1 0 14224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__493__I
timestamp 1698431365
transform 1 0 15568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__A1
timestamp 1698431365
transform -1 0 14672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__I
timestamp 1698431365
transform 1 0 14448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__I
timestamp 1698431365
transform 1 0 9184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__I
timestamp 1698431365
transform 1 0 14896 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__A1
timestamp 1698431365
transform 1 0 12992 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__B2
timestamp 1698431365
transform 1 0 11312 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__C
timestamp 1698431365
transform 1 0 11984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A1
timestamp 1698431365
transform 1 0 10080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__I
timestamp 1698431365
transform -1 0 14672 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__I
timestamp 1698431365
transform 1 0 13104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__A2
timestamp 1698431365
transform 1 0 11872 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__C1
timestamp 1698431365
transform -1 0 15344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__I
timestamp 1698431365
transform -1 0 16576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__A1
timestamp 1698431365
transform 1 0 18480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__B2
timestamp 1698431365
transform -1 0 19152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__526__C
timestamp 1698431365
transform 1 0 11760 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__A1
timestamp 1698431365
transform 1 0 17472 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A1
timestamp 1698431365
transform -1 0 10752 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__B2
timestamp 1698431365
transform 1 0 9296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__A1
timestamp 1698431365
transform -1 0 12432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__B2
timestamp 1698431365
transform -1 0 11200 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__A1
timestamp 1698431365
transform -1 0 16912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__B2
timestamp 1698431365
transform -1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__A2
timestamp 1698431365
transform 1 0 14000 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__C1
timestamp 1698431365
transform 1 0 17024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__542__I
timestamp 1698431365
transform 1 0 15120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__A1
timestamp 1698431365
transform -1 0 8400 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__A1
timestamp 1698431365
transform -1 0 10640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__549__A1
timestamp 1698431365
transform -1 0 13552 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__549__B2
timestamp 1698431365
transform 1 0 11872 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__B2
timestamp 1698431365
transform 1 0 13552 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__C1
timestamp 1698431365
transform -1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__556__B2
timestamp 1698431365
transform -1 0 16688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__A2
timestamp 1698431365
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__B1
timestamp 1698431365
transform 1 0 13776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__C1
timestamp 1698431365
transform -1 0 17024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__A1
timestamp 1698431365
transform 1 0 11312 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__560__A1
timestamp 1698431365
transform 1 0 6720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__563__A1
timestamp 1698431365
transform 1 0 14672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__563__C2
timestamp 1698431365
transform 1 0 14224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__B2
timestamp 1698431365
transform 1 0 14896 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__C1
timestamp 1698431365
transform -1 0 16016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__565__A1
timestamp 1698431365
transform -1 0 17808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__566__A1
timestamp 1698431365
transform -1 0 18144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__566__B2
timestamp 1698431365
transform 1 0 17472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__C
timestamp 1698431365
transform 1 0 12880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__572__A1
timestamp 1698431365
transform -1 0 14224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__572__B
timestamp 1698431365
transform 1 0 10864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__572__C
timestamp 1698431365
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__573__A1
timestamp 1698431365
transform 1 0 14560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__573__B2
timestamp 1698431365
transform 1 0 14784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__574__B2
timestamp 1698431365
transform -1 0 10640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__575__A1
timestamp 1698431365
transform 1 0 15008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__576__A1
timestamp 1698431365
transform 1 0 18368 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__C
timestamp 1698431365
transform 1 0 12208 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A1
timestamp 1698431365
transform 1 0 15232 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A2
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__583__A1
timestamp 1698431365
transform 1 0 28000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__583__A3
timestamp 1698431365
transform 1 0 28448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__A2
timestamp 1698431365
transform 1 0 14560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__A2
timestamp 1698431365
transform 1 0 31808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__586__A1
timestamp 1698431365
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__I
timestamp 1698431365
transform -1 0 27440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__A3
timestamp 1698431365
transform -1 0 29456 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__A2
timestamp 1698431365
transform 1 0 16464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__591__A2
timestamp 1698431365
transform -1 0 34496 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__592__A1
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__A1
timestamp 1698431365
transform 1 0 30688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__A3
timestamp 1698431365
transform 1 0 30240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__597__A2
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__598__A1
timestamp 1698431365
transform -1 0 35168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__A1
timestamp 1698431365
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__A1
timestamp 1698431365
transform 1 0 15008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__A2
timestamp 1698431365
transform 1 0 15232 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__I
timestamp 1698431365
transform 1 0 8960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__605__A1
timestamp 1698431365
transform -1 0 6832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__607__A2
timestamp 1698431365
transform 1 0 6608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__611__I
timestamp 1698431365
transform -1 0 10976 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__614__A1
timestamp 1698431365
transform 1 0 4704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__615__C
timestamp 1698431365
transform -1 0 4704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__616__I
timestamp 1698431365
transform 1 0 7056 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__617__A1
timestamp 1698431365
transform -1 0 6608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__622__A1
timestamp 1698431365
transform -1 0 2464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__I
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__625__C
timestamp 1698431365
transform 1 0 3248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__626__I
timestamp 1698431365
transform 1 0 9968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__A1
timestamp 1698431365
transform -1 0 10304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__631__A1
timestamp 1698431365
transform 1 0 5600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__C
timestamp 1698431365
transform 1 0 3696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__633__I
timestamp 1698431365
transform 1 0 21840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__634__A1
timestamp 1698431365
transform 1 0 11088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__638__A1
timestamp 1698431365
transform 1 0 8512 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__638__A2
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__640__I
timestamp 1698431365
transform 1 0 19936 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__642__B
timestamp 1698431365
transform -1 0 7616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__644__A2
timestamp 1698431365
transform 1 0 13104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__A1
timestamp 1698431365
transform 1 0 7728 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__A2
timestamp 1698431365
transform 1 0 12320 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__649__A1
timestamp 1698431365
transform -1 0 6160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__650__B
timestamp 1698431365
transform 1 0 7392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__651__I
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__652__A1
timestamp 1698431365
transform -1 0 11312 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__654__B
timestamp 1698431365
transform 1 0 10304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__655__A1
timestamp 1698431365
transform 1 0 6608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__A1
timestamp 1698431365
transform -1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__657__B
timestamp 1698431365
transform 1 0 6944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__658__I
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__659__A1
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__664__A1
timestamp 1698431365
transform 1 0 10976 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__666__A1
timestamp 1698431365
transform 1 0 11872 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__668__I
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__669__A1
timestamp 1698431365
transform 1 0 14112 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__672__A1
timestamp 1698431365
transform 1 0 11984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__A1
timestamp 1698431365
transform 1 0 12320 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__681__I
timestamp 1698431365
transform 1 0 16240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__682__A1
timestamp 1698431365
transform -1 0 15456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__685__A1
timestamp 1698431365
transform 1 0 15344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__688__A1
timestamp 1698431365
transform 1 0 17024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__C
timestamp 1698431365
transform 1 0 18592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__690__A1
timestamp 1698431365
transform -1 0 15904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__691__A1
timestamp 1698431365
transform 1 0 19936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__693__A1
timestamp 1698431365
transform -1 0 18928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__694__A1
timestamp 1698431365
transform 1 0 15792 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__696__A1
timestamp 1698431365
transform -1 0 19712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__A1
timestamp 1698431365
transform 1 0 19712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__701__A1
timestamp 1698431365
transform 1 0 21392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__701__A2
timestamp 1698431365
transform 1 0 20160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__702__A1
timestamp 1698431365
transform 1 0 23520 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__704__A1
timestamp 1698431365
transform -1 0 22736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__704__A2
timestamp 1698431365
transform 1 0 22960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__705__A1
timestamp 1698431365
transform 1 0 22960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__707__A1
timestamp 1698431365
transform 1 0 20720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__707__A2
timestamp 1698431365
transform 1 0 20272 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__A1
timestamp 1698431365
transform -1 0 21504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__710__A1
timestamp 1698431365
transform -1 0 17472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__710__A2
timestamp 1698431365
transform 1 0 17696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__712__A1
timestamp 1698431365
transform -1 0 16128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__A2
timestamp 1698431365
transform -1 0 16352 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__I
timestamp 1698431365
transform -1 0 26992 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__719__A1
timestamp 1698431365
transform 1 0 19488 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__722__A1
timestamp 1698431365
transform 1 0 16240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__725__A1
timestamp 1698431365
transform -1 0 19040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__729__A1
timestamp 1698431365
transform 1 0 21952 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__731__A1
timestamp 1698431365
transform 1 0 23408 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__734__A1
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__A1
timestamp 1698431365
transform 1 0 22960 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__738__A1
timestamp 1698431365
transform 1 0 24976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__740__A1
timestamp 1698431365
transform 1 0 20832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__743__A1
timestamp 1698431365
transform 1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__743__A2
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__745__A1
timestamp 1698431365
transform -1 0 19936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__746__A1
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__746__A2
timestamp 1698431365
transform 1 0 15120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__751__A1
timestamp 1698431365
transform 1 0 21168 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__752__A1
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__754__A1
timestamp 1698431365
transform -1 0 20384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__757__A1
timestamp 1698431365
transform 1 0 19600 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__761__A1
timestamp 1698431365
transform -1 0 27216 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__763__A1
timestamp 1698431365
transform -1 0 28672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__766__A1
timestamp 1698431365
transform 1 0 28224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__767__A1
timestamp 1698431365
transform 1 0 27664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__770__A1
timestamp 1698431365
transform -1 0 31584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__772__A1
timestamp 1698431365
transform -1 0 29008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__775__A1
timestamp 1698431365
transform 1 0 18480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__778__A1
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__779__A1
timestamp 1698431365
transform 1 0 15232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__779__C
timestamp 1698431365
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__780__A1
timestamp 1698431365
transform 1 0 17360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__780__A2
timestamp 1698431365
transform 1 0 18032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__782__A1
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__783__A1
timestamp 1698431365
transform 1 0 18928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__786__A1
timestamp 1698431365
transform 1 0 19712 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__788__A1
timestamp 1698431365
transform 1 0 19264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__789__A1
timestamp 1698431365
transform 1 0 22512 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__791__A1
timestamp 1698431365
transform 1 0 24640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__793__A1
timestamp 1698431365
transform 1 0 25648 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__794__A1
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__796__A1
timestamp 1698431365
transform 1 0 25200 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__797__A1
timestamp 1698431365
transform 1 0 29232 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__800__A1
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__802__A1
timestamp 1698431365
transform 1 0 15680 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__803__A1
timestamp 1698431365
transform 1 0 18704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__804__A1
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__804__A2
timestamp 1698431365
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__807__A1
timestamp 1698431365
transform 1 0 23520 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__809__I
timestamp 1698431365
transform 1 0 24752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__810__A1
timestamp 1698431365
transform 1 0 20272 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__812__A1
timestamp 1698431365
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__815__A1
timestamp 1698431365
transform 1 0 22736 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__816__A1
timestamp 1698431365
transform 1 0 24304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__819__A1
timestamp 1698431365
transform 1 0 27328 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__821__A1
timestamp 1698431365
transform 1 0 28784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__822__A1
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__824__A1
timestamp 1698431365
transform 1 0 30352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__824__C
timestamp 1698431365
transform 1 0 28000 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__825__A1
timestamp 1698431365
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__826__A1
timestamp 1698431365
transform 1 0 31360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__826__C
timestamp 1698431365
transform 1 0 29904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__827__A1
timestamp 1698431365
transform 1 0 30912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__827__A2
timestamp 1698431365
transform -1 0 31360 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__828__A1
timestamp 1698431365
transform 1 0 33600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__828__A2
timestamp 1698431365
transform -1 0 33936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__829__CLK
timestamp 1698431365
transform 1 0 32928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__831__CLK
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__838__CLK
timestamp 1698431365
transform 1 0 35616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__839__CLK
timestamp 1698431365
transform 1 0 32928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__840__CLK
timestamp 1698431365
transform 1 0 34944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__841__CLK
timestamp 1698431365
transform -1 0 7392 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__843__CLK
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__844__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__845__CLK
timestamp 1698431365
transform 1 0 11760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__846__CLK
timestamp 1698431365
transform 1 0 5712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__847__CLK
timestamp 1698431365
transform 1 0 11984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__848__CLK
timestamp 1698431365
transform 1 0 7616 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__849__CLK
timestamp 1698431365
transform 1 0 4368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__850__CLK
timestamp 1698431365
transform 1 0 10640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__851__CLK
timestamp 1698431365
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__852__CLK
timestamp 1698431365
transform 1 0 14448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__853__CLK
timestamp 1698431365
transform -1 0 10640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__854__CLK
timestamp 1698431365
transform 1 0 14224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__855__CLK
timestamp 1698431365
transform 1 0 10192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__865__CLK
timestamp 1698431365
transform -1 0 15456 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__866__CLK
timestamp 1698431365
transform 1 0 17360 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__867__CLK
timestamp 1698431365
transform 1 0 12880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__868__CLK
timestamp 1698431365
transform 1 0 16912 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__873__CLK
timestamp 1698431365
transform 1 0 23072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__875__CLK
timestamp 1698431365
transform 1 0 25200 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__877__CLK
timestamp 1698431365
transform 1 0 29232 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__879__CLK
timestamp 1698431365
transform 1 0 33264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__880__CLK
timestamp 1698431365
transform 1 0 30800 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__888__CLK
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__889__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__890__CLK
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__891__CLK
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__892__CLK
timestamp 1698431365
transform 1 0 25536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__893__CLK
timestamp 1698431365
transform 1 0 28896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__894__CLK
timestamp 1698431365
transform 1 0 32032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__895__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__896__CLK
timestamp 1698431365
transform 1 0 34272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__897__CLK
timestamp 1698431365
transform 1 0 34160 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__898__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 25648 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 23968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 19152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 26320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 16576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 26880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 1792 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 1792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 2464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 33376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 1792 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 3136 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 2688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 1792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 2688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 3136 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 4704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 7168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 15120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 17360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 18480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 19600 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 21280 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 5600 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 6944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 9632 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 9408 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 11536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 11312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 13104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 14000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 42672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 42672 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 43120 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 42224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 42672 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 42672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output48_I
timestamp 1698431365
transform 1 0 23856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output50_I
timestamp 1698431365
transform 1 0 27552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output79_I
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output80_I
timestamp 1698431365
transform 1 0 36624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output81_I
timestamp 1698431365
transform -1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24528 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1698431365
transform -1 0 22848 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1698431365
transform 1 0 26544 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1698431365
transform -1 0 16128 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1698431365
transform 1 0 11200 0 -1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1698431365
transform 1 0 27104 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_6
timestamp 1698431365
transform 1 0 2016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_40
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_74
timestamp 1698431365
transform 1 0 9632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_108
timestamp 1698431365
transform 1 0 13440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142
timestamp 1698431365
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698431365
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_232
timestamp 1698431365
transform 1 0 27328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698431365
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_266
timestamp 1698431365
transform 1 0 31136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_282
timestamp 1698431365
transform 1 0 32928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_284 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33152 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_291 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_299
timestamp 1698431365
transform 1 0 34832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_334
timestamp 1698431365
transform 1 0 38752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_368
timestamp 1698431365
transform 1 0 42560 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_372
timestamp 1698431365
transform 1 0 43008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_374
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_10
timestamp 1698431365
transform 1 0 2464 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_76
timestamp 1698431365
transform 1 0 9856 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_79
timestamp 1698431365
transform 1 0 10192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_135
timestamp 1698431365
transform 1 0 16464 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_171
timestamp 1698431365
transform 1 0 20496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_199
timestamp 1698431365
transform 1 0 23632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698431365
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698431365
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_247
timestamp 1698431365
transform 1 0 29008 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_251
timestamp 1698431365
transform 1 0 29456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_286 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_302
timestamp 1698431365
transform 1 0 35168 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_310
timestamp 1698431365
transform 1 0 36064 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_343
timestamp 1698431365
transform 1 0 39760 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_347
timestamp 1698431365
transform 1 0 40208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_360
timestamp 1698431365
transform 1 0 41664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_362
timestamp 1698431365
transform 1 0 41888 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_373
timestamp 1698431365
transform 1 0 43120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_8
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_12
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_28
timestamp 1698431365
transform 1 0 4480 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_32
timestamp 1698431365
transform 1 0 4928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_53
timestamp 1698431365
transform 1 0 7280 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_57
timestamp 1698431365
transform 1 0 7728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_98
timestamp 1698431365
transform 1 0 12320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_102
timestamp 1698431365
transform 1 0 12768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_136
timestamp 1698431365
transform 1 0 16576 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_144
timestamp 1698431365
transform 1 0 17472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_349
timestamp 1698431365
transform 1 0 40432 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_365
timestamp 1698431365
transform 1 0 42224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_8
timestamp 1698431365
transform 1 0 2240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_12
timestamp 1698431365
transform 1 0 2688 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_44
timestamp 1698431365
transform 1 0 6272 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_60
timestamp 1698431365
transform 1 0 8064 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_68
timestamp 1698431365
transform 1 0 8960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_76
timestamp 1698431365
transform 1 0 9856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_78
timestamp 1698431365
transform 1 0 10080 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_81
timestamp 1698431365
transform 1 0 10416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_83
timestamp 1698431365
transform 1 0 10640 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_113
timestamp 1698431365
transform 1 0 14000 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_117
timestamp 1698431365
transform 1 0 14448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_133
timestamp 1698431365
transform 1 0 16240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_137
timestamp 1698431365
transform 1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_168
timestamp 1698431365
transform 1 0 20160 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_176
timestamp 1698431365
transform 1 0 21056 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_208
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_368
timestamp 1698431365
transform 1 0 42560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_372
timestamp 1698431365
transform 1 0 43008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_374
timestamp 1698431365
transform 1 0 43232 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_45
timestamp 1698431365
transform 1 0 6384 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_49
timestamp 1698431365
transform 1 0 6832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_92
timestamp 1698431365
transform 1 0 11648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_96
timestamp 1698431365
transform 1 0 12096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_116
timestamp 1698431365
transform 1 0 14336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_120
timestamp 1698431365
transform 1 0 14784 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_150
timestamp 1698431365
transform 1 0 18144 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_154
timestamp 1698431365
transform 1 0 18592 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_157
timestamp 1698431365
transform 1 0 18928 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_161
timestamp 1698431365
transform 1 0 19376 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_164
timestamp 1698431365
transform 1 0 19712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_168
timestamp 1698431365
transform 1 0 20160 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_349
timestamp 1698431365
transform 1 0 40432 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_365
timestamp 1698431365
transform 1 0 42224 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_373
timestamp 1698431365
transform 1 0 43120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_8
timestamp 1698431365
transform 1 0 2240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_12
timestamp 1698431365
transform 1 0 2688 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_44
timestamp 1698431365
transform 1 0 6272 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_60
timestamp 1698431365
transform 1 0 8064 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_76
timestamp 1698431365
transform 1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_78
timestamp 1698431365
transform 1 0 10080 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_84
timestamp 1698431365
transform 1 0 10752 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_88
timestamp 1698431365
transform 1 0 11200 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_92
timestamp 1698431365
transform 1 0 11648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_107
timestamp 1698431365
transform 1 0 13328 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_123
timestamp 1698431365
transform 1 0 15120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_161
timestamp 1698431365
transform 1 0 19376 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_165
timestamp 1698431365
transform 1 0 19824 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_174
timestamp 1698431365
transform 1 0 20832 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_185
timestamp 1698431365
transform 1 0 22064 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_191
timestamp 1698431365
transform 1 0 22736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_195
timestamp 1698431365
transform 1 0 23184 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_203
timestamp 1698431365
transform 1 0 24080 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_207
timestamp 1698431365
transform 1 0 24528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_368
timestamp 1698431365
transform 1 0 42560 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_372
timestamp 1698431365
transform 1 0 43008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_374
timestamp 1698431365
transform 1 0 43232 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_73
timestamp 1698431365
transform 1 0 9520 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_93
timestamp 1698431365
transform 1 0 11760 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_97
timestamp 1698431365
transform 1 0 12208 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_112
timestamp 1698431365
transform 1 0 13888 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_116
timestamp 1698431365
transform 1 0 14336 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_124
timestamp 1698431365
transform 1 0 15232 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_128
timestamp 1698431365
transform 1 0 15680 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_131
timestamp 1698431365
transform 1 0 16016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_148
timestamp 1698431365
transform 1 0 17920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_150
timestamp 1698431365
transform 1 0 18144 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_162
timestamp 1698431365
transform 1 0 19488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_196
timestamp 1698431365
transform 1 0 23296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_200
timestamp 1698431365
transform 1 0 23744 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_232
timestamp 1698431365
transform 1 0 27328 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_240
timestamp 1698431365
transform 1 0 28224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_349
timestamp 1698431365
transform 1 0 40432 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_365
timestamp 1698431365
transform 1 0 42224 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_373
timestamp 1698431365
transform 1 0 43120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_8
timestamp 1698431365
transform 1 0 2240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_12
timestamp 1698431365
transform 1 0 2688 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_28
timestamp 1698431365
transform 1 0 4480 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_36
timestamp 1698431365
transform 1 0 5376 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_40
timestamp 1698431365
transform 1 0 5824 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_43
timestamp 1698431365
transform 1 0 6160 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_59
timestamp 1698431365
transform 1 0 7952 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_85
timestamp 1698431365
transform 1 0 10864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_93
timestamp 1698431365
transform 1 0 11760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_97
timestamp 1698431365
transform 1 0 12208 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_113
timestamp 1698431365
transform 1 0 14000 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_121
timestamp 1698431365
transform 1 0 14896 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_123
timestamp 1698431365
transform 1 0 15120 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_126
timestamp 1698431365
transform 1 0 15456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_200
timestamp 1698431365
transform 1 0 23744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_204
timestamp 1698431365
transform 1 0 24192 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_208
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_270
timestamp 1698431365
transform 1 0 31584 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_368
timestamp 1698431365
transform 1 0 42560 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_372
timestamp 1698431365
transform 1 0 43008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_374
timestamp 1698431365
transform 1 0 43232 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_10
timestamp 1698431365
transform 1 0 2464 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_26
timestamp 1698431365
transform 1 0 4256 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_30
timestamp 1698431365
transform 1 0 4704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_32
timestamp 1698431365
transform 1 0 4928 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_41
timestamp 1698431365
transform 1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_48
timestamp 1698431365
transform 1 0 6720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_52
timestamp 1698431365
transform 1 0 7168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_56
timestamp 1698431365
transform 1 0 7616 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_72
timestamp 1698431365
transform 1 0 9408 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_80
timestamp 1698431365
transform 1 0 10304 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_84
timestamp 1698431365
transform 1 0 10752 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_111
timestamp 1698431365
transform 1 0 13776 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_115
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_117
timestamp 1698431365
transform 1 0 14448 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_126
timestamp 1698431365
transform 1 0 15456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_128
timestamp 1698431365
transform 1 0 15680 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_158
timestamp 1698431365
transform 1 0 19040 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_162
timestamp 1698431365
transform 1 0 19488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_166
timestamp 1698431365
transform 1 0 19936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_223
timestamp 1698431365
transform 1 0 26320 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_231
timestamp 1698431365
transform 1 0 27216 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_235
timestamp 1698431365
transform 1 0 27664 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_243
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_256
timestamp 1698431365
transform 1 0 30016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_260
timestamp 1698431365
transform 1 0 30464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_264
timestamp 1698431365
transform 1 0 30912 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_296
timestamp 1698431365
transform 1 0 34496 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_312
timestamp 1698431365
transform 1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_349
timestamp 1698431365
transform 1 0 40432 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_365
timestamp 1698431365
transform 1 0 42224 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_373
timestamp 1698431365
transform 1 0 43120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_35
timestamp 1698431365
transform 1 0 5264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_55
timestamp 1698431365
transform 1 0 7504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_59
timestamp 1698431365
transform 1 0 7952 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_67
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_82
timestamp 1698431365
transform 1 0 10528 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_85
timestamp 1698431365
transform 1 0 10864 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_115
timestamp 1698431365
transform 1 0 14224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_119
timestamp 1698431365
transform 1 0 14672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_148
timestamp 1698431365
transform 1 0 17920 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_156
timestamp 1698431365
transform 1 0 18816 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_166
timestamp 1698431365
transform 1 0 19936 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_168
timestamp 1698431365
transform 1 0 20160 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_171
timestamp 1698431365
transform 1 0 20496 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_175
timestamp 1698431365
transform 1 0 20944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_189
timestamp 1698431365
transform 1 0 22512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_199
timestamp 1698431365
transform 1 0 23632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_203
timestamp 1698431365
transform 1 0 24080 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_228
timestamp 1698431365
transform 1 0 26880 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_260
timestamp 1698431365
transform 1 0 30464 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_368
timestamp 1698431365
transform 1 0 42560 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_372
timestamp 1698431365
transform 1 0 43008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_374
timestamp 1698431365
transform 1 0 43232 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_83
timestamp 1698431365
transform 1 0 10640 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_157
timestamp 1698431365
transform 1 0 18928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_161
timestamp 1698431365
transform 1 0 19376 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_169
timestamp 1698431365
transform 1 0 20272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_191
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_195
timestamp 1698431365
transform 1 0 23184 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_227
timestamp 1698431365
transform 1 0 26768 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_349
timestamp 1698431365
transform 1 0 40432 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_365
timestamp 1698431365
transform 1 0 42224 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_373
timestamp 1698431365
transform 1 0 43120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_10
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_14
timestamp 1698431365
transform 1 0 2912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_18
timestamp 1698431365
transform 1 0 3360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_26
timestamp 1698431365
transform 1 0 4256 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_29
timestamp 1698431365
transform 1 0 4592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_33
timestamp 1698431365
transform 1 0 5040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_47
timestamp 1698431365
transform 1 0 6608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_54
timestamp 1698431365
transform 1 0 7392 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_58
timestamp 1698431365
transform 1 0 7840 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_62
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_64
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_85
timestamp 1698431365
transform 1 0 10864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_89
timestamp 1698431365
transform 1 0 11312 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_105
timestamp 1698431365
transform 1 0 13104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_117
timestamp 1698431365
transform 1 0 14448 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_121
timestamp 1698431365
transform 1 0 14896 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_129
timestamp 1698431365
transform 1 0 15792 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_133
timestamp 1698431365
transform 1 0 16240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_135
timestamp 1698431365
transform 1 0 16464 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_152
timestamp 1698431365
transform 1 0 18368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_156
timestamp 1698431365
transform 1 0 18816 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_188
timestamp 1698431365
transform 1 0 22400 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_204
timestamp 1698431365
transform 1 0 24192 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_222
timestamp 1698431365
transform 1 0 26208 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_275
timestamp 1698431365
transform 1 0 32144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698431365
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_368
timestamp 1698431365
transform 1 0 42560 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_372
timestamp 1698431365
transform 1 0 43008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_374
timestamp 1698431365
transform 1 0 43232 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_24
timestamp 1698431365
transform 1 0 4032 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_39
timestamp 1698431365
transform 1 0 5712 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_42
timestamp 1698431365
transform 1 0 6048 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_46
timestamp 1698431365
transform 1 0 6496 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_49
timestamp 1698431365
transform 1 0 6832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_53
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_69
timestamp 1698431365
transform 1 0 9072 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_77
timestamp 1698431365
transform 1 0 9968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_79
timestamp 1698431365
transform 1 0 10192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_82
timestamp 1698431365
transform 1 0 10528 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_98
timestamp 1698431365
transform 1 0 12320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_119
timestamp 1698431365
transform 1 0 14672 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_123
timestamp 1698431365
transform 1 0 15120 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_148
timestamp 1698431365
transform 1 0 17920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_150
timestamp 1698431365
transform 1 0 18144 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_161
timestamp 1698431365
transform 1 0 19376 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_165
timestamp 1698431365
transform 1 0 19824 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_219
timestamp 1698431365
transform 1 0 25872 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_227
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_229
timestamp 1698431365
transform 1 0 26992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698431365
transform 1 0 28000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698431365
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_349
timestamp 1698431365
transform 1 0 40432 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_365
timestamp 1698431365
transform 1 0 42224 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_373
timestamp 1698431365
transform 1 0 43120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_10
timestamp 1698431365
transform 1 0 2464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_28
timestamp 1698431365
transform 1 0 4480 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_36
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_40
timestamp 1698431365
transform 1 0 5824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_58
timestamp 1698431365
transform 1 0 7840 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_92
timestamp 1698431365
transform 1 0 11648 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_96
timestamp 1698431365
transform 1 0 12096 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_112
timestamp 1698431365
transform 1 0 13888 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_116
timestamp 1698431365
transform 1 0 14336 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_119
timestamp 1698431365
transform 1 0 14672 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_123
timestamp 1698431365
transform 1 0 15120 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_126
timestamp 1698431365
transform 1 0 15456 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_134
timestamp 1698431365
transform 1 0 16352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_187
timestamp 1698431365
transform 1 0 22288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_191
timestamp 1698431365
transform 1 0 22736 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698431365
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_258
timestamp 1698431365
transform 1 0 30240 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698431365
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_360
timestamp 1698431365
transform 1 0 41664 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_364
timestamp 1698431365
transform 1 0 42112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_366
timestamp 1698431365
transform 1 0 42336 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_12
timestamp 1698431365
transform 1 0 2688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_22
timestamp 1698431365
transform 1 0 3808 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_63
timestamp 1698431365
transform 1 0 8400 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_71
timestamp 1698431365
transform 1 0 9296 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_75
timestamp 1698431365
transform 1 0 9744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_87
timestamp 1698431365
transform 1 0 11088 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_96
timestamp 1698431365
transform 1 0 12096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_100
timestamp 1698431365
transform 1 0 12544 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_122
timestamp 1698431365
transform 1 0 15008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_145
timestamp 1698431365
transform 1 0 17584 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_161
timestamp 1698431365
transform 1 0 19376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_169
timestamp 1698431365
transform 1 0 20272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_187
timestamp 1698431365
transform 1 0 22288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_206
timestamp 1698431365
transform 1 0 24416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_210
timestamp 1698431365
transform 1 0 24864 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_212
timestamp 1698431365
transform 1 0 25088 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_215
timestamp 1698431365
transform 1 0 25424 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698431365
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_251
timestamp 1698431365
transform 1 0 29456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_287
timestamp 1698431365
transform 1 0 33488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_303
timestamp 1698431365
transform 1 0 35280 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_349
timestamp 1698431365
transform 1 0 40432 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_365
timestamp 1698431365
transform 1 0 42224 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_373
timestamp 1698431365
transform 1 0 43120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_11
timestamp 1698431365
transform 1 0 2576 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_59
timestamp 1698431365
transform 1 0 7952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_61
timestamp 1698431365
transform 1 0 8176 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_82
timestamp 1698431365
transform 1 0 10528 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_103
timestamp 1698431365
transform 1 0 12880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_107
timestamp 1698431365
transform 1 0 13328 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_115
timestamp 1698431365
transform 1 0 14224 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_119
timestamp 1698431365
transform 1 0 14672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_121
timestamp 1698431365
transform 1 0 14896 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_124
timestamp 1698431365
transform 1 0 15232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_147
timestamp 1698431365
transform 1 0 17808 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_151
timestamp 1698431365
transform 1 0 18256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_155
timestamp 1698431365
transform 1 0 18704 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_163
timestamp 1698431365
transform 1 0 19600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_173
timestamp 1698431365
transform 1 0 20720 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_177
timestamp 1698431365
transform 1 0 21168 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_183
timestamp 1698431365
transform 1 0 21840 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_190
timestamp 1698431365
transform 1 0 22624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_194
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_239
timestamp 1698431365
transform 1 0 28112 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_241
timestamp 1698431365
transform 1 0 28336 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_247
timestamp 1698431365
transform 1 0 29008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698431365
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_368
timestamp 1698431365
transform 1 0 42560 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_372
timestamp 1698431365
transform 1 0 43008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_374
timestamp 1698431365
transform 1 0 43232 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_4
timestamp 1698431365
transform 1 0 1792 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_21
timestamp 1698431365
transform 1 0 3696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_25
timestamp 1698431365
transform 1 0 4144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_74
timestamp 1698431365
transform 1 0 9632 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_82
timestamp 1698431365
transform 1 0 10528 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_97
timestamp 1698431365
transform 1 0 12208 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_109
timestamp 1698431365
transform 1 0 13552 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_141
timestamp 1698431365
transform 1 0 17136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_153
timestamp 1698431365
transform 1 0 18480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_164
timestamp 1698431365
transform 1 0 19712 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_187
timestamp 1698431365
transform 1 0 22288 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_219
timestamp 1698431365
transform 1 0 25872 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_227
timestamp 1698431365
transform 1 0 26768 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_230
timestamp 1698431365
transform 1 0 27104 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_238
timestamp 1698431365
transform 1 0 28000 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_260
timestamp 1698431365
transform 1 0 30464 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_268
timestamp 1698431365
transform 1 0 31360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_272
timestamp 1698431365
transform 1 0 31808 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_304
timestamp 1698431365
transform 1 0 35392 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_308
timestamp 1698431365
transform 1 0 35840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_349
timestamp 1698431365
transform 1 0 40432 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_365
timestamp 1698431365
transform 1 0 42224 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_373
timestamp 1698431365
transform 1 0 43120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_4
timestamp 1698431365
transform 1 0 1792 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_67
timestamp 1698431365
transform 1 0 8848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_86
timestamp 1698431365
transform 1 0 10976 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_135
timestamp 1698431365
transform 1 0 16464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_153
timestamp 1698431365
transform 1 0 18480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_157
timestamp 1698431365
transform 1 0 18928 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_165
timestamp 1698431365
transform 1 0 19824 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_177
timestamp 1698431365
transform 1 0 21168 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_193
timestamp 1698431365
transform 1 0 22960 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_228
timestamp 1698431365
transform 1 0 26880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_230
timestamp 1698431365
transform 1 0 27104 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_239
timestamp 1698431365
transform 1 0 28112 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_251
timestamp 1698431365
transform 1 0 29456 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_267
timestamp 1698431365
transform 1 0 31248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698431365
transform 1 0 32144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_288
timestamp 1698431365
transform 1 0 33600 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_320
timestamp 1698431365
transform 1 0 37184 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_336
timestamp 1698431365
transform 1 0 38976 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_344
timestamp 1698431365
transform 1 0 39872 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_348
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_368
timestamp 1698431365
transform 1 0 42560 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_372
timestamp 1698431365
transform 1 0 43008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_374
timestamp 1698431365
transform 1 0 43232 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_80
timestamp 1698431365
transform 1 0 10304 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_94
timestamp 1698431365
transform 1 0 11872 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_102
timestamp 1698431365
transform 1 0 12768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_115
timestamp 1698431365
transform 1 0 14224 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_131
timestamp 1698431365
transform 1 0 16016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_137
timestamp 1698431365
transform 1 0 16688 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_141
timestamp 1698431365
transform 1 0 17136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_158
timestamp 1698431365
transform 1 0 19040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_162
timestamp 1698431365
transform 1 0 19488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_166
timestamp 1698431365
transform 1 0 19936 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_181
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_214
timestamp 1698431365
transform 1 0 25312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_218
timestamp 1698431365
transform 1 0 25760 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_234
timestamp 1698431365
transform 1 0 27552 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_242
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_255
timestamp 1698431365
transform 1 0 29904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_259
timestamp 1698431365
transform 1 0 30352 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_261
timestamp 1698431365
transform 1 0 30576 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_291
timestamp 1698431365
transform 1 0 33936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_295
timestamp 1698431365
transform 1 0 34384 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_349
timestamp 1698431365
transform 1 0 40432 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_365
timestamp 1698431365
transform 1 0 42224 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_373
timestamp 1698431365
transform 1 0 43120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_14
timestamp 1698431365
transform 1 0 2912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698431365
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698431365
transform 1 0 10304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_84
timestamp 1698431365
transform 1 0 10752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_87
timestamp 1698431365
transform 1 0 11088 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_113
timestamp 1698431365
transform 1 0 14000 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_117
timestamp 1698431365
transform 1 0 14448 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_121
timestamp 1698431365
transform 1 0 14896 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_129
timestamp 1698431365
transform 1 0 15792 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_133
timestamp 1698431365
transform 1 0 16240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_135
timestamp 1698431365
transform 1 0 16464 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_165
timestamp 1698431365
transform 1 0 19824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_189
timestamp 1698431365
transform 1 0 22512 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_196
timestamp 1698431365
transform 1 0 23296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_200
timestamp 1698431365
transform 1 0 23744 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_272
timestamp 1698431365
transform 1 0 31808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_290
timestamp 1698431365
transform 1 0 33824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_294
timestamp 1698431365
transform 1 0 34272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_297
timestamp 1698431365
transform 1 0 34608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_299
timestamp 1698431365
transform 1 0 34832 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_333
timestamp 1698431365
transform 1 0 38640 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_368
timestamp 1698431365
transform 1 0 42560 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_372
timestamp 1698431365
transform 1 0 43008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_374
timestamp 1698431365
transform 1 0 43232 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_28
timestamp 1698431365
transform 1 0 4480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_54
timestamp 1698431365
transform 1 0 7392 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_70
timestamp 1698431365
transform 1 0 9184 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_74
timestamp 1698431365
transform 1 0 9632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_84
timestamp 1698431365
transform 1 0 10752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_86
timestamp 1698431365
transform 1 0 10976 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_116
timestamp 1698431365
transform 1 0 14336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_120
timestamp 1698431365
transform 1 0 14784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_124
timestamp 1698431365
transform 1 0 15232 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_203
timestamp 1698431365
transform 1 0 24080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_207
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_211
timestamp 1698431365
transform 1 0 24976 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_321
timestamp 1698431365
transform 1 0 37296 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_353
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_369
timestamp 1698431365
transform 1 0 42672 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_373
timestamp 1698431365
transform 1 0 43120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_28
timestamp 1698431365
transform 1 0 4480 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_36
timestamp 1698431365
transform 1 0 5376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_38
timestamp 1698431365
transform 1 0 5600 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_47
timestamp 1698431365
transform 1 0 6608 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_63
timestamp 1698431365
transform 1 0 8400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_92
timestamp 1698431365
transform 1 0 11648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_94
timestamp 1698431365
transform 1 0 11872 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_118
timestamp 1698431365
transform 1 0 14560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_122
timestamp 1698431365
transform 1 0 15008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_146
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_154
timestamp 1698431365
transform 1 0 18592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_158
timestamp 1698431365
transform 1 0 19040 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_188
timestamp 1698431365
transform 1 0 22400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_190
timestamp 1698431365
transform 1 0 22624 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_205
timestamp 1698431365
transform 1 0 24304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_216
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_232
timestamp 1698431365
transform 1 0 27328 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_236
timestamp 1698431365
transform 1 0 27776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_240
timestamp 1698431365
transform 1 0 28224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_244
timestamp 1698431365
transform 1 0 28672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_260
timestamp 1698431365
transform 1 0 30464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_264
timestamp 1698431365
transform 1 0 30912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_312
timestamp 1698431365
transform 1 0 36288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_316
timestamp 1698431365
transform 1 0 36736 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_348
timestamp 1698431365
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_368
timestamp 1698431365
transform 1 0 42560 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_372
timestamp 1698431365
transform 1 0 43008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_374
timestamp 1698431365
transform 1 0 43232 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_31
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_53
timestamp 1698431365
transform 1 0 7280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_55
timestamp 1698431365
transform 1 0 7504 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_62
timestamp 1698431365
transform 1 0 8288 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_80
timestamp 1698431365
transform 1 0 10304 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_96
timestamp 1698431365
transform 1 0 12096 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_98
timestamp 1698431365
transform 1 0 12320 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_112
timestamp 1698431365
transform 1 0 13888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_114
timestamp 1698431365
transform 1 0 14112 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_142
timestamp 1698431365
transform 1 0 17248 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_144
timestamp 1698431365
transform 1 0 17472 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_154
timestamp 1698431365
transform 1 0 18592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_158
timestamp 1698431365
transform 1 0 19040 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_187
timestamp 1698431365
transform 1 0 22288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_211
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_215
timestamp 1698431365
transform 1 0 25424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_219
timestamp 1698431365
transform 1 0 25872 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_227
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_239
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_256
timestamp 1698431365
transform 1 0 30016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_260
timestamp 1698431365
transform 1 0 30464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_266
timestamp 1698431365
transform 1 0 31136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_280
timestamp 1698431365
transform 1 0 32704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_284
timestamp 1698431365
transform 1 0 33152 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_288
timestamp 1698431365
transform 1 0 33600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_298
timestamp 1698431365
transform 1 0 34720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_302
timestamp 1698431365
transform 1 0 35168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_310
timestamp 1698431365
transform 1 0 36064 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_349
timestamp 1698431365
transform 1 0 40432 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_365
timestamp 1698431365
transform 1 0 42224 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_373
timestamp 1698431365
transform 1 0 43120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_28
timestamp 1698431365
transform 1 0 4480 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_36
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_40
timestamp 1698431365
transform 1 0 5824 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_91
timestamp 1698431365
transform 1 0 11536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_95
timestamp 1698431365
transform 1 0 11984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_99
timestamp 1698431365
transform 1 0 12432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_135
timestamp 1698431365
transform 1 0 16464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_137
timestamp 1698431365
transform 1 0 16688 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_148
timestamp 1698431365
transform 1 0 17920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_152
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_156
timestamp 1698431365
transform 1 0 18816 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698431365
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_221
timestamp 1698431365
transform 1 0 26096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_243
timestamp 1698431365
transform 1 0 28560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_247
timestamp 1698431365
transform 1 0 29008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_251
timestamp 1698431365
transform 1 0 29456 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_267
timestamp 1698431365
transform 1 0 31248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_271
timestamp 1698431365
transform 1 0 31696 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698431365
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698431365
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_290
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_296
timestamp 1698431365
transform 1 0 34496 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_328
timestamp 1698431365
transform 1 0 38080 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_344
timestamp 1698431365
transform 1 0 39872 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_348
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_368
timestamp 1698431365
transform 1 0 42560 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_372
timestamp 1698431365
transform 1 0 43008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_374
timestamp 1698431365
transform 1 0 43232 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698431365
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_69
timestamp 1698431365
transform 1 0 9072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_93
timestamp 1698431365
transform 1 0 11760 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_97
timestamp 1698431365
transform 1 0 12208 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_117
timestamp 1698431365
transform 1 0 14448 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_125
timestamp 1698431365
transform 1 0 15344 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_157
timestamp 1698431365
transform 1 0 18928 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_186
timestamp 1698431365
transform 1 0 22176 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_188
timestamp 1698431365
transform 1 0 22400 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_218
timestamp 1698431365
transform 1 0 25760 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_222
timestamp 1698431365
transform 1 0 26208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_240
timestamp 1698431365
transform 1 0 28224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_242
timestamp 1698431365
transform 1 0 28448 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_253
timestamp 1698431365
transform 1 0 29680 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_257
timestamp 1698431365
transform 1 0 30128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_261
timestamp 1698431365
transform 1 0 30576 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_277
timestamp 1698431365
transform 1 0 32368 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_285
timestamp 1698431365
transform 1 0 33264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_295
timestamp 1698431365
transform 1 0 34384 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_302
timestamp 1698431365
transform 1 0 35168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_306
timestamp 1698431365
transform 1 0 35616 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_349
timestamp 1698431365
transform 1 0 40432 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_365
timestamp 1698431365
transform 1 0 42224 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_373
timestamp 1698431365
transform 1 0 43120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_18
timestamp 1698431365
transform 1 0 3360 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_48
timestamp 1698431365
transform 1 0 6720 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_56
timestamp 1698431365
transform 1 0 7616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_65
timestamp 1698431365
transform 1 0 8624 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_80
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_84
timestamp 1698431365
transform 1 0 10752 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_116
timestamp 1698431365
transform 1 0 14336 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_132
timestamp 1698431365
transform 1 0 16128 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_158
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_170
timestamp 1698431365
transform 1 0 20384 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_202
timestamp 1698431365
transform 1 0 23968 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_228
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_234
timestamp 1698431365
transform 1 0 27552 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_266
timestamp 1698431365
transform 1 0 31136 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_270
timestamp 1698431365
transform 1 0 31584 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_317
timestamp 1698431365
transform 1 0 36848 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_360
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_364
timestamp 1698431365
transform 1 0 42112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_366
timestamp 1698431365
transform 1 0 42336 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_73
timestamp 1698431365
transform 1 0 9520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_94
timestamp 1698431365
transform 1 0 11872 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_102
timestamp 1698431365
transform 1 0 12768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_133
timestamp 1698431365
transform 1 0 16240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_148
timestamp 1698431365
transform 1 0 17920 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_156
timestamp 1698431365
transform 1 0 18816 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_249
timestamp 1698431365
transform 1 0 29232 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_258
timestamp 1698431365
transform 1 0 30240 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_274
timestamp 1698431365
transform 1 0 32032 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_349
timestamp 1698431365
transform 1 0 40432 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_365
timestamp 1698431365
transform 1 0 42224 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_373
timestamp 1698431365
transform 1 0 43120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_28
timestamp 1698431365
transform 1 0 4480 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_44
timestamp 1698431365
transform 1 0 6272 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_46
timestamp 1698431365
transform 1 0 6496 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_58
timestamp 1698431365
transform 1 0 7840 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_89
timestamp 1698431365
transform 1 0 11312 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_93
timestamp 1698431365
transform 1 0 11760 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_105
timestamp 1698431365
transform 1 0 13104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_109
timestamp 1698431365
transform 1 0 13552 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_128
timestamp 1698431365
transform 1 0 15680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_130
timestamp 1698431365
transform 1 0 15904 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_158
timestamp 1698431365
transform 1 0 19040 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_165
timestamp 1698431365
transform 1 0 19824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_169
timestamp 1698431365
transform 1 0 20272 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_185
timestamp 1698431365
transform 1 0 22064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_193
timestamp 1698431365
transform 1 0 22960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_199
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_203
timestamp 1698431365
transform 1 0 24080 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698431365
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_214
timestamp 1698431365
transform 1 0 25312 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_244
timestamp 1698431365
transform 1 0 28672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_248
timestamp 1698431365
transform 1 0 29120 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_286
timestamp 1698431365
transform 1 0 33376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_297
timestamp 1698431365
transform 1 0 34608 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_329
timestamp 1698431365
transform 1 0 38192 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_345
timestamp 1698431365
transform 1 0 39984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_368
timestamp 1698431365
transform 1 0 42560 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_372
timestamp 1698431365
transform 1 0 43008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_374
timestamp 1698431365
transform 1 0 43232 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_31
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_42
timestamp 1698431365
transform 1 0 6048 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_61
timestamp 1698431365
transform 1 0 8176 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_77
timestamp 1698431365
transform 1 0 9968 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_83
timestamp 1698431365
transform 1 0 10640 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_91
timestamp 1698431365
transform 1 0 11536 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_103
timestamp 1698431365
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_123
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_130
timestamp 1698431365
transform 1 0 15904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_142
timestamp 1698431365
transform 1 0 17248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_146
timestamp 1698431365
transform 1 0 17696 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_162
timestamp 1698431365
transform 1 0 19488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_166
timestamp 1698431365
transform 1 0 19936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_182
timestamp 1698431365
transform 1 0 21728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_192
timestamp 1698431365
transform 1 0 22848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_196
timestamp 1698431365
transform 1 0 23296 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_232
timestamp 1698431365
transform 1 0 27328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698431365
transform 1 0 28224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_263
timestamp 1698431365
transform 1 0 30800 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_267
timestamp 1698431365
transform 1 0 31248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_273
timestamp 1698431365
transform 1 0 31920 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_277
timestamp 1698431365
transform 1 0 32368 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_285
timestamp 1698431365
transform 1 0 33264 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_291
timestamp 1698431365
transform 1 0 33936 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_307
timestamp 1698431365
transform 1 0 35728 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_349
timestamp 1698431365
transform 1 0 40432 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_365
timestamp 1698431365
transform 1 0 42224 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_373
timestamp 1698431365
transform 1 0 43120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_18
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_49
timestamp 1698431365
transform 1 0 6832 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_61
timestamp 1698431365
transform 1 0 8176 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_88
timestamp 1698431365
transform 1 0 11200 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_102
timestamp 1698431365
transform 1 0 12768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_106
timestamp 1698431365
transform 1 0 13216 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_122
timestamp 1698431365
transform 1 0 15008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_124
timestamp 1698431365
transform 1 0 15232 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_150
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_158
timestamp 1698431365
transform 1 0 19040 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_199
timestamp 1698431365
transform 1 0 23632 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_228
timestamp 1698431365
transform 1 0 26880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_230
timestamp 1698431365
transform 1 0 27104 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_239
timestamp 1698431365
transform 1 0 28112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_243
timestamp 1698431365
transform 1 0 28560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_247
timestamp 1698431365
transform 1 0 29008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_251
timestamp 1698431365
transform 1 0 29456 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_267
timestamp 1698431365
transform 1 0 31248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_275
timestamp 1698431365
transform 1 0 32144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_292
timestamp 1698431365
transform 1 0 34048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_296
timestamp 1698431365
transform 1 0 34496 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_328
timestamp 1698431365
transform 1 0 38080 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_344
timestamp 1698431365
transform 1 0 39872 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_368
timestamp 1698431365
transform 1 0 42560 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_372
timestamp 1698431365
transform 1 0 43008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_374
timestamp 1698431365
transform 1 0 43232 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698431365
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_51
timestamp 1698431365
transform 1 0 7056 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_60
timestamp 1698431365
transform 1 0 8064 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_115
timestamp 1698431365
transform 1 0 14224 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_143
timestamp 1698431365
transform 1 0 17360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_147
timestamp 1698431365
transform 1 0 17808 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_163
timestamp 1698431365
transform 1 0 19600 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_167
timestamp 1698431365
transform 1 0 20048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_169
timestamp 1698431365
transform 1 0 20272 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_211
timestamp 1698431365
transform 1 0 24976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_215
timestamp 1698431365
transform 1 0 25424 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_260
timestamp 1698431365
transform 1 0 30464 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_290
timestamp 1698431365
transform 1 0 33824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_300
timestamp 1698431365
transform 1 0 34944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_304
timestamp 1698431365
transform 1 0 35392 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_349
timestamp 1698431365
transform 1 0 40432 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_365
timestamp 1698431365
transform 1 0 42224 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_373
timestamp 1698431365
transform 1 0 43120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_28
timestamp 1698431365
transform 1 0 4480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_32
timestamp 1698431365
transform 1 0 4928 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_64
timestamp 1698431365
transform 1 0 8512 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_101
timestamp 1698431365
transform 1 0 12656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_105
timestamp 1698431365
transform 1 0 13104 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_121
timestamp 1698431365
transform 1 0 14896 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_129
timestamp 1698431365
transform 1 0 15792 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_135
timestamp 1698431365
transform 1 0 16464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_178
timestamp 1698431365
transform 1 0 21280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_188
timestamp 1698431365
transform 1 0 22400 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698431365
transform 1 0 24192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_311
timestamp 1698431365
transform 1 0 36176 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_343
timestamp 1698431365
transform 1 0 39760 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_347
timestamp 1698431365
transform 1 0 40208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_368
timestamp 1698431365
transform 1 0 42560 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_372
timestamp 1698431365
transform 1 0 43008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_374
timestamp 1698431365
transform 1 0 43232 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_72
timestamp 1698431365
transform 1 0 9408 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_76
timestamp 1698431365
transform 1 0 9856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_78
timestamp 1698431365
transform 1 0 10080 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_83
timestamp 1698431365
transform 1 0 10640 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_95
timestamp 1698431365
transform 1 0 11984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_99
timestamp 1698431365
transform 1 0 12432 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_103
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_117
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_121
timestamp 1698431365
transform 1 0 14896 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_125
timestamp 1698431365
transform 1 0 15344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_141
timestamp 1698431365
transform 1 0 17136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_153
timestamp 1698431365
transform 1 0 18480 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_161
timestamp 1698431365
transform 1 0 19376 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_165
timestamp 1698431365
transform 1 0 19824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_167
timestamp 1698431365
transform 1 0 20048 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_209
timestamp 1698431365
transform 1 0 24752 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_225
timestamp 1698431365
transform 1 0 26544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_229
timestamp 1698431365
transform 1 0 26992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_240
timestamp 1698431365
transform 1 0 28224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_252
timestamp 1698431365
transform 1 0 29568 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_266
timestamp 1698431365
transform 1 0 31136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_270
timestamp 1698431365
transform 1 0 31584 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_278
timestamp 1698431365
transform 1 0 32480 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_283
timestamp 1698431365
transform 1 0 33040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_287
timestamp 1698431365
transform 1 0 33488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_291
timestamp 1698431365
transform 1 0 33936 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_307
timestamp 1698431365
transform 1 0 35728 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_349
timestamp 1698431365
transform 1 0 40432 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_365
timestamp 1698431365
transform 1 0 42224 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_373
timestamp 1698431365
transform 1 0 43120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_36
timestamp 1698431365
transform 1 0 5376 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_45
timestamp 1698431365
transform 1 0 6384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_49
timestamp 1698431365
transform 1 0 6832 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_65
timestamp 1698431365
transform 1 0 8624 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_69
timestamp 1698431365
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_132
timestamp 1698431365
transform 1 0 16128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_134
timestamp 1698431365
transform 1 0 16352 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_151
timestamp 1698431365
transform 1 0 18256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_155
timestamp 1698431365
transform 1 0 18704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_159
timestamp 1698431365
transform 1 0 19152 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_167
timestamp 1698431365
transform 1 0 20048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_175
timestamp 1698431365
transform 1 0 20944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_179
timestamp 1698431365
transform 1 0 21392 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_195
timestamp 1698431365
transform 1 0 23184 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_203
timestamp 1698431365
transform 1 0 24080 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_207
timestamp 1698431365
transform 1 0 24528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_227
timestamp 1698431365
transform 1 0 26768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_231
timestamp 1698431365
transform 1 0 27216 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_239
timestamp 1698431365
transform 1 0 28112 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_243
timestamp 1698431365
transform 1 0 28560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_247
timestamp 1698431365
transform 1 0 29008 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_290
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_294
timestamp 1698431365
transform 1 0 34272 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_326
timestamp 1698431365
transform 1 0 37856 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_342
timestamp 1698431365
transform 1 0 39648 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_368
timestamp 1698431365
transform 1 0 42560 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_372
timestamp 1698431365
transform 1 0 43008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_374
timestamp 1698431365
transform 1 0 43232 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_33
timestamp 1698431365
transform 1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_46
timestamp 1698431365
transform 1 0 6496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_50
timestamp 1698431365
transform 1 0 6944 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_82
timestamp 1698431365
transform 1 0 10528 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_99
timestamp 1698431365
transform 1 0 12432 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_150
timestamp 1698431365
transform 1 0 18144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_154
timestamp 1698431365
transform 1 0 18592 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_162
timestamp 1698431365
transform 1 0 19488 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_179
timestamp 1698431365
transform 1 0 21392 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_191
timestamp 1698431365
transform 1 0 22736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_195
timestamp 1698431365
transform 1 0 23184 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_232
timestamp 1698431365
transform 1 0 27328 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_238
timestamp 1698431365
transform 1 0 28000 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_252
timestamp 1698431365
transform 1 0 29568 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_261
timestamp 1698431365
transform 1 0 30576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_302
timestamp 1698431365
transform 1 0 35168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_310
timestamp 1698431365
transform 1 0 36064 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_349
timestamp 1698431365
transform 1 0 40432 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_365
timestamp 1698431365
transform 1 0 42224 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_373
timestamp 1698431365
transform 1 0 43120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_6
timestamp 1698431365
transform 1 0 2016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_26
timestamp 1698431365
transform 1 0 4256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_30
timestamp 1698431365
transform 1 0 4704 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_34
timestamp 1698431365
transform 1 0 5152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_38
timestamp 1698431365
transform 1 0 5600 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_74
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_85
timestamp 1698431365
transform 1 0 10864 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_89
timestamp 1698431365
transform 1 0 11312 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_99
timestamp 1698431365
transform 1 0 12432 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_107
timestamp 1698431365
transform 1 0 13328 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_111
timestamp 1698431365
transform 1 0 13776 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_118
timestamp 1698431365
transform 1 0 14560 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_126
timestamp 1698431365
transform 1 0 15456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_130
timestamp 1698431365
transform 1 0 15904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_134
timestamp 1698431365
transform 1 0 16352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_138
timestamp 1698431365
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_158
timestamp 1698431365
transform 1 0 19040 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_166
timestamp 1698431365
transform 1 0 19936 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_180
timestamp 1698431365
transform 1 0 21504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_182
timestamp 1698431365
transform 1 0 21728 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_191
timestamp 1698431365
transform 1 0 22736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_197
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_201
timestamp 1698431365
transform 1 0 23856 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_203
timestamp 1698431365
transform 1 0 24080 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_228
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_232
timestamp 1698431365
transform 1 0 27328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_234
timestamp 1698431365
transform 1 0 27552 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_250
timestamp 1698431365
transform 1 0 29344 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_258
timestamp 1698431365
transform 1 0 30240 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_262
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_274
timestamp 1698431365
transform 1 0 32032 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_278
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698431365
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_368
timestamp 1698431365
transform 1 0 42560 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_372
timestamp 1698431365
transform 1 0 43008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_374
timestamp 1698431365
transform 1 0 43232 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_28
timestamp 1698431365
transform 1 0 4480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_32
timestamp 1698431365
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_64
timestamp 1698431365
transform 1 0 8512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_68
timestamp 1698431365
transform 1 0 8960 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_87
timestamp 1698431365
transform 1 0 11088 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_91
timestamp 1698431365
transform 1 0 11536 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_99
timestamp 1698431365
transform 1 0 12432 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_103
timestamp 1698431365
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_111
timestamp 1698431365
transform 1 0 13776 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_115
timestamp 1698431365
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_119
timestamp 1698431365
transform 1 0 14672 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_137
timestamp 1698431365
transform 1 0 16688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_139
timestamp 1698431365
transform 1 0 16912 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_142
timestamp 1698431365
transform 1 0 17248 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_214
timestamp 1698431365
transform 1 0 25312 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_230
timestamp 1698431365
transform 1 0 27104 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_238
timestamp 1698431365
transform 1 0 28000 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_242
timestamp 1698431365
transform 1 0 28448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_276
timestamp 1698431365
transform 1 0 32256 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_308
timestamp 1698431365
transform 1 0 35840 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_323
timestamp 1698431365
transform 1 0 37520 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_355
timestamp 1698431365
transform 1 0 41104 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_363
timestamp 1698431365
transform 1 0 42000 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_4
timestamp 1698431365
transform 1 0 1792 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_15
timestamp 1698431365
transform 1 0 3024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_19
timestamp 1698431365
transform 1 0 3472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_23
timestamp 1698431365
transform 1 0 3920 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_31
timestamp 1698431365
transform 1 0 4816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_33
timestamp 1698431365
transform 1 0 5040 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_48
timestamp 1698431365
transform 1 0 6720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_76
timestamp 1698431365
transform 1 0 9856 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_103
timestamp 1698431365
transform 1 0 12880 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_152
timestamp 1698431365
transform 1 0 18368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_156
timestamp 1698431365
transform 1 0 18816 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_188
timestamp 1698431365
transform 1 0 22400 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_204
timestamp 1698431365
transform 1 0 24192 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_262
timestamp 1698431365
transform 1 0 30688 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_278
timestamp 1698431365
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_368
timestamp 1698431365
transform 1 0 42560 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_372
timestamp 1698431365
transform 1 0 43008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_374
timestamp 1698431365
transform 1 0 43232 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_33
timestamp 1698431365
transform 1 0 5040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_47
timestamp 1698431365
transform 1 0 6608 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_50
timestamp 1698431365
transform 1 0 6944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_54
timestamp 1698431365
transform 1 0 7392 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_62
timestamp 1698431365
transform 1 0 8288 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_70
timestamp 1698431365
transform 1 0 9184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_95
timestamp 1698431365
transform 1 0 11984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_99
timestamp 1698431365
transform 1 0 12432 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_167
timestamp 1698431365
transform 1 0 20048 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_193
timestamp 1698431365
transform 1 0 22960 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_201
timestamp 1698431365
transform 1 0 23856 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_203
timestamp 1698431365
transform 1 0 24080 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_219
timestamp 1698431365
transform 1 0 25872 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_223
timestamp 1698431365
transform 1 0 26320 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_227
timestamp 1698431365
transform 1 0 26768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_229
timestamp 1698431365
transform 1 0 26992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_255
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_259
timestamp 1698431365
transform 1 0 30352 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_291
timestamp 1698431365
transform 1 0 33936 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_307
timestamp 1698431365
transform 1 0 35728 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_349
timestamp 1698431365
transform 1 0 40432 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_365
timestamp 1698431365
transform 1 0 42224 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_373
timestamp 1698431365
transform 1 0 43120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_4
timestamp 1698431365
transform 1 0 1792 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_59
timestamp 1698431365
transform 1 0 7952 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_63
timestamp 1698431365
transform 1 0 8400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_67
timestamp 1698431365
transform 1 0 8848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_80
timestamp 1698431365
transform 1 0 10304 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_83
timestamp 1698431365
transform 1 0 10640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_87
timestamp 1698431365
transform 1 0 11088 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_138
timestamp 1698431365
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_150
timestamp 1698431365
transform 1 0 18144 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_156
timestamp 1698431365
transform 1 0 18816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_175
timestamp 1698431365
transform 1 0 20944 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_191
timestamp 1698431365
transform 1 0 22736 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_204
timestamp 1698431365
transform 1 0 24192 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_230
timestamp 1698431365
transform 1 0 27104 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_253
timestamp 1698431365
transform 1 0 29680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_257
timestamp 1698431365
transform 1 0 30128 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_286
timestamp 1698431365
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_368
timestamp 1698431365
transform 1 0 42560 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_372
timestamp 1698431365
transform 1 0 43008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_374
timestamp 1698431365
transform 1 0 43232 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_47
timestamp 1698431365
transform 1 0 6608 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_56
timestamp 1698431365
transform 1 0 7616 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_72
timestamp 1698431365
transform 1 0 9408 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_76
timestamp 1698431365
transform 1 0 9856 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_84
timestamp 1698431365
transform 1 0 10752 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_99
timestamp 1698431365
transform 1 0 12432 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_103
timestamp 1698431365
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_111
timestamp 1698431365
transform 1 0 13776 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_115
timestamp 1698431365
transform 1 0 14224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_132
timestamp 1698431365
transform 1 0 16128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_136
timestamp 1698431365
transform 1 0 16576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_140
timestamp 1698431365
transform 1 0 17024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_144
timestamp 1698431365
transform 1 0 17472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_148
timestamp 1698431365
transform 1 0 17920 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_164
timestamp 1698431365
transform 1 0 19712 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_166
timestamp 1698431365
transform 1 0 19936 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_181
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_183
timestamp 1698431365
transform 1 0 21840 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_191
timestamp 1698431365
transform 1 0 22736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_195
timestamp 1698431365
transform 1 0 23184 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_210
timestamp 1698431365
transform 1 0 24864 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_214
timestamp 1698431365
transform 1 0 25312 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_349
timestamp 1698431365
transform 1 0 40432 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_365
timestamp 1698431365
transform 1 0 42224 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_373
timestamp 1698431365
transform 1 0 43120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_36
timestamp 1698431365
transform 1 0 5376 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_40
timestamp 1698431365
transform 1 0 5824 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_44
timestamp 1698431365
transform 1 0 6272 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_46
timestamp 1698431365
transform 1 0 6496 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_59
timestamp 1698431365
transform 1 0 7952 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_63
timestamp 1698431365
transform 1 0 8400 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_86
timestamp 1698431365
transform 1 0 10976 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_121
timestamp 1698431365
transform 1 0 14896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_125
timestamp 1698431365
transform 1 0 15344 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_129
timestamp 1698431365
transform 1 0 15792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_131
timestamp 1698431365
transform 1 0 16016 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_134
timestamp 1698431365
transform 1 0 16352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1698431365
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_144
timestamp 1698431365
transform 1 0 17472 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_151
timestamp 1698431365
transform 1 0 18256 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_167
timestamp 1698431365
transform 1 0 20048 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_171
timestamp 1698431365
transform 1 0 20496 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_173
timestamp 1698431365
transform 1 0 20720 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_220
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_236
timestamp 1698431365
transform 1 0 27776 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_273
timestamp 1698431365
transform 1 0 31920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_277
timestamp 1698431365
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_368
timestamp 1698431365
transform 1 0 42560 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_372
timestamp 1698431365
transform 1 0 43008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_374
timestamp 1698431365
transform 1 0 43232 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_28
timestamp 1698431365
transform 1 0 4480 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_51
timestamp 1698431365
transform 1 0 7056 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_68
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_70
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_76
timestamp 1698431365
transform 1 0 9856 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_80
timestamp 1698431365
transform 1 0 10304 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_96
timestamp 1698431365
transform 1 0 12096 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_115
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_119
timestamp 1698431365
transform 1 0 14672 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_128
timestamp 1698431365
transform 1 0 15680 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_132
timestamp 1698431365
transform 1 0 16128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_140
timestamp 1698431365
transform 1 0 17024 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_148
timestamp 1698431365
transform 1 0 17920 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_154
timestamp 1698431365
transform 1 0 18592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_158
timestamp 1698431365
transform 1 0 19040 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_166
timestamp 1698431365
transform 1 0 19936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_187
timestamp 1698431365
transform 1 0 22288 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_209
timestamp 1698431365
transform 1 0 24752 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_213
timestamp 1698431365
transform 1 0 25200 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_215
timestamp 1698431365
transform 1 0 25424 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_28
timestamp 1698431365
transform 1 0 4480 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_44
timestamp 1698431365
transform 1 0 6272 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_85
timestamp 1698431365
transform 1 0 10864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_89
timestamp 1698431365
transform 1 0 11312 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_93
timestamp 1698431365
transform 1 0 11760 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_95
timestamp 1698431365
transform 1 0 11984 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_121
timestamp 1698431365
transform 1 0 14896 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_127
timestamp 1698431365
transform 1 0 15568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_131
timestamp 1698431365
transform 1 0 16016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_135
timestamp 1698431365
transform 1 0 16464 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_160
timestamp 1698431365
transform 1 0 19264 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_164
timestamp 1698431365
transform 1 0 19712 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_196
timestamp 1698431365
transform 1 0 23296 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_204
timestamp 1698431365
transform 1 0 24192 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_368
timestamp 1698431365
transform 1 0 42560 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_372
timestamp 1698431365
transform 1 0 43008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_374
timestamp 1698431365
transform 1 0 43232 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_28
timestamp 1698431365
transform 1 0 4480 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_41
timestamp 1698431365
transform 1 0 5936 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_49
timestamp 1698431365
transform 1 0 6832 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_53
timestamp 1698431365
transform 1 0 7280 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_91
timestamp 1698431365
transform 1 0 11536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_95
timestamp 1698431365
transform 1 0 11984 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_109
timestamp 1698431365
transform 1 0 13552 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_136
timestamp 1698431365
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698431365
transform 1 0 16800 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_185
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_189
timestamp 1698431365
transform 1 0 22512 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_220
timestamp 1698431365
transform 1 0 25984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_224
timestamp 1698431365
transform 1 0 26432 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_240
timestamp 1698431365
transform 1 0 28224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_242
timestamp 1698431365
transform 1 0 28448 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_253
timestamp 1698431365
transform 1 0 29680 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_271
timestamp 1698431365
transform 1 0 31696 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_303
timestamp 1698431365
transform 1 0 35280 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_333
timestamp 1698431365
transform 1 0 38640 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_341
timestamp 1698431365
transform 1 0 39536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_369
timestamp 1698431365
transform 1 0 42672 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_373
timestamp 1698431365
transform 1 0 43120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_80
timestamp 1698431365
transform 1 0 10304 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_88
timestamp 1698431365
transform 1 0 11200 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_92
timestamp 1698431365
transform 1 0 11648 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_94
timestamp 1698431365
transform 1 0 11872 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_146
timestamp 1698431365
transform 1 0 17696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_156
timestamp 1698431365
transform 1 0 18816 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_160
timestamp 1698431365
transform 1 0 19264 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_165
timestamp 1698431365
transform 1 0 19824 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_172
timestamp 1698431365
transform 1 0 20608 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_188
timestamp 1698431365
transform 1 0 22400 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_196
timestamp 1698431365
transform 1 0 23296 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_220
timestamp 1698431365
transform 1 0 25984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_224
timestamp 1698431365
transform 1 0 26432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_228
timestamp 1698431365
transform 1 0 26880 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_232
timestamp 1698431365
transform 1 0 27328 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_239
timestamp 1698431365
transform 1 0 28112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_243
timestamp 1698431365
transform 1 0 28560 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_277
timestamp 1698431365
transform 1 0 32368 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_279
timestamp 1698431365
transform 1 0 32592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_288
timestamp 1698431365
transform 1 0 33600 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_296
timestamp 1698431365
transform 1 0 34496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_300
timestamp 1698431365
transform 1 0 34944 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_302
timestamp 1698431365
transform 1 0 35168 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_335
timestamp 1698431365
transform 1 0 38864 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_342
timestamp 1698431365
transform 1 0 39648 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_368
timestamp 1698431365
transform 1 0 42560 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_372
timestamp 1698431365
transform 1 0 43008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_374
timestamp 1698431365
transform 1 0 43232 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_31
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_41
timestamp 1698431365
transform 1 0 5936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_45
timestamp 1698431365
transform 1 0 6384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_47
timestamp 1698431365
transform 1 0 6608 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_50
timestamp 1698431365
transform 1 0 6944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_54
timestamp 1698431365
transform 1 0 7392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_93
timestamp 1698431365
transform 1 0 11760 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_97
timestamp 1698431365
transform 1 0 12208 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_136
timestamp 1698431365
transform 1 0 16576 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_140
timestamp 1698431365
transform 1 0 17024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_142
timestamp 1698431365
transform 1 0 17248 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698431365
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_183
timestamp 1698431365
transform 1 0 21840 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_227
timestamp 1698431365
transform 1 0 26768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_305
timestamp 1698431365
transform 1 0 35504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_307
timestamp 1698431365
transform 1 0 35728 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698431365
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_369
timestamp 1698431365
transform 1 0 42672 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_373
timestamp 1698431365
transform 1 0 43120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_60
timestamp 1698431365
transform 1 0 8064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_68
timestamp 1698431365
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_84
timestamp 1698431365
transform 1 0 10752 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_88
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_103
timestamp 1698431365
transform 1 0 12880 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_107
timestamp 1698431365
transform 1 0 13328 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_113
timestamp 1698431365
transform 1 0 14000 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_121
timestamp 1698431365
transform 1 0 14896 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_123
timestamp 1698431365
transform 1 0 15120 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_126
timestamp 1698431365
transform 1 0 15456 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_134
timestamp 1698431365
transform 1 0 16352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_138
timestamp 1698431365
transform 1 0 16800 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_174
timestamp 1698431365
transform 1 0 20832 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_180
timestamp 1698431365
transform 1 0 21504 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_196
timestamp 1698431365
transform 1 0 23296 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_271
timestamp 1698431365
transform 1 0 31696 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_334
timestamp 1698431365
transform 1 0 38752 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_368
timestamp 1698431365
transform 1 0 42560 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_372
timestamp 1698431365
transform 1 0 43008 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_36
timestamp 1698431365
transform 1 0 5376 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_40
timestamp 1698431365
transform 1 0 5824 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_48
timestamp 1698431365
transform 1 0 6720 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_52
timestamp 1698431365
transform 1 0 7168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_54
timestamp 1698431365
transform 1 0 7392 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_61
timestamp 1698431365
transform 1 0 8176 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_70
timestamp 1698431365
transform 1 0 9184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_74
timestamp 1698431365
transform 1 0 9632 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_82
timestamp 1698431365
transform 1 0 10528 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_86
timestamp 1698431365
transform 1 0 10976 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_110
timestamp 1698431365
transform 1 0 13664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_112
timestamp 1698431365
transform 1 0 13888 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_119
timestamp 1698431365
transform 1 0 14672 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_129
timestamp 1698431365
transform 1 0 15792 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_138
timestamp 1698431365
transform 1 0 16800 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_140
timestamp 1698431365
transform 1 0 17024 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_149
timestamp 1698431365
transform 1 0 18032 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_159
timestamp 1698431365
transform 1 0 19152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_169
timestamp 1698431365
transform 1 0 20272 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_232
timestamp 1698431365
transform 1 0 27328 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_236
timestamp 1698431365
transform 1 0 27776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_266
timestamp 1698431365
transform 1 0 31136 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_270
timestamp 1698431365
transform 1 0 31584 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_300
timestamp 1698431365
transform 1 0 34944 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_304
timestamp 1698431365
transform 1 0 35392 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_334
timestamp 1698431365
transform 1 0 38752 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_338
timestamp 1698431365
transform 1 0 39200 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_368
timestamp 1698431365
transform 1 0 42560 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold1
timestamp 1698431365
transform -1 0 11984 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold2
timestamp 1698431365
transform -1 0 7280 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold3
timestamp 1698431365
transform -1 0 5824 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold4
timestamp 1698431365
transform -1 0 8288 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold5
timestamp 1698431365
transform -1 0 8512 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold6
timestamp 1698431365
transform -1 0 8176 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold7
timestamp 1698431365
transform -1 0 8288 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold8
timestamp 1698431365
transform -1 0 12208 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input6
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 33936 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input9
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input12
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input13
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input16
timestamp 1698431365
transform 1 0 8176 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 15120 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 15904 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 18032 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 19152 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 20272 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 21280 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 4592 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 4480 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 7392 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 8288 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 8288 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 12208 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input29
timestamp 1698431365
transform 1 0 11984 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 14672 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 43344 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 43344 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 43344 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input35
timestamp 1698431365
transform 1 0 42224 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input36
timestamp 1698431365
transform -1 0 43344 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform -1 0 43344 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output38 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4480 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output39
timestamp 1698431365
transform -1 0 4480 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output40
timestamp 1698431365
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output41
timestamp 1698431365
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output42
timestamp 1698431365
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output43
timestamp 1698431365
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output44
timestamp 1698431365
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output45
timestamp 1698431365
transform -1 0 4480 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output46
timestamp 1698431365
transform -1 0 4480 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output47
timestamp 1698431365
transform -1 0 5152 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output48
timestamp 1698431365
transform -1 0 23632 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output49
timestamp 1698431365
transform 1 0 21280 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output50
timestamp 1698431365
transform -1 0 27328 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51
timestamp 1698431365
transform -1 0 29008 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output52
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53
timestamp 1698431365
transform 1 0 29680 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698431365
transform -1 0 6272 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698431365
transform 1 0 6272 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output57
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output58
timestamp 1698431365
transform -1 0 13552 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output59
timestamp 1698431365
transform 1 0 13552 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output60
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output61
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output62
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output63
timestamp 1698431365
transform 1 0 21280 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output64
timestamp 1698431365
transform 1 0 35840 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output65
timestamp 1698431365
transform 1 0 35840 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output66
timestamp 1698431365
transform 1 0 35280 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output67
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output68
timestamp 1698431365
transform 1 0 39648 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output69
timestamp 1698431365
transform 1 0 39760 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output70
timestamp 1698431365
transform 1 0 22960 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output71
timestamp 1698431365
transform 1 0 24416 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output72
timestamp 1698431365
transform 1 0 25200 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output73
timestamp 1698431365
transform 1 0 28224 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output74
timestamp 1698431365
transform 1 0 28112 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output75
timestamp 1698431365
transform -1 0 31920 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output76
timestamp 1698431365
transform 1 0 32032 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output77
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output78
timestamp 1698431365
transform 1 0 31920 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output79
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output80
timestamp 1698431365
transform 1 0 36848 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output81
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output82
timestamp 1698431365
transform -1 0 4480 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output83
timestamp 1698431365
transform -1 0 4480 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output84
timestamp 1698431365
transform -1 0 4480 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output85
timestamp 1698431365
transform -1 0 4480 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output86
timestamp 1698431365
transform -1 0 4480 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output87
timestamp 1698431365
transform -1 0 4480 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output88
timestamp 1698431365
transform -1 0 4480 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output89
timestamp 1698431365
transform -1 0 7392 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output90
timestamp 1698431365
transform 1 0 39760 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output91
timestamp 1698431365
transform 1 0 40432 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_49 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 43568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 43568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 43568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 43568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 43568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 43568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 43568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 43568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 43568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 43568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 43568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 43568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 43568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 43568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 43568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 43568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 43568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 43568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 43568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 43568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 43568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 43568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 43568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 43568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 43568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 43568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 43568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 43568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 43568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 43568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 43568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 43568 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 43568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 43568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 43568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 43568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 43568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 43568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 43568 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 43568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 43568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 43568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 43568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 43568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 43568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 43568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 43568 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 43568 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 43568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_108
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_109
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_110
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_111
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_112
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_113
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_114
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_115
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_117
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_118
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_119
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_120
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_121
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_122
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_123
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_124
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_125
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_126
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_127
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_128
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_129
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_130
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_131
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_132
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_133
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_134
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_135
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_136
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_137
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_138
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_139
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_140
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_141
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_142
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_143
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_144
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_145
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_146
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_147
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_148
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_149
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_150
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_151
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_152
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_153
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_154
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_155
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_156
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_157
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_158
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_159
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_160
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_161
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_162
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_163
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_164
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_165
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_166
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_167
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_168
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_169
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_170
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_171
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_172
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_173
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_174
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_175
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_176
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_177
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_178
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_179
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_180
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_181
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_182
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_183
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_184
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_185
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_186
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_187
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_188
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_189
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_190
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_191
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_192
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_193
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_194
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_195
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_196
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_197
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_198
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_199
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_200
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_201
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_202
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_203
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_204
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_205
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_208
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_209
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_210
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_212
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_213
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_214
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_215
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_216
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_217
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_218
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_219
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_220
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_221
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_222
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_223
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_224
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_225
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_226
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_227
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_228
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_229
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_230
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_231
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_232
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_233
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_234
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_235
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_236
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_237
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_238
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_239
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_240
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_241
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_242
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_243
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_244
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_245
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_246
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_247
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_248
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_249
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_250
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_251
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_252
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_253
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_254
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_255
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_256
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_257
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_258
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_259
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_260
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_261
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_262
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_263
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_264
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_265
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_266
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_267
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_268
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_269
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_270
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_271
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_272
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_273
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_274
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_275
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_276
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_277
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_278
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_279
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_280
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_281
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_282
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_283
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_284
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_285
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_286
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_287
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_288
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_289
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_290
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_291
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_292
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_293
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_294
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_295
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_296
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_297
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_298
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_299
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_300
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_301
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_302
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_303
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_304
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_305
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_306
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_307
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_308
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_309
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_310
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_311
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_312
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_313
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_314
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_315
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_316
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_317
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_318
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_319
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_320
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_321
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_322
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_323
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_324
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_325
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_326
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_327
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_328
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_329
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_330
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_331
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_332
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_333
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_334
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_335
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_336
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_337
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_338
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_339
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_340
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_341
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_342
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_343
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_344
timestamp 1698431365
transform 1 0 8960 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_345
timestamp 1698431365
transform 1 0 12768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_346
timestamp 1698431365
transform 1 0 16576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_347
timestamp 1698431365
transform 1 0 20384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_348
timestamp 1698431365
transform 1 0 24192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_349
timestamp 1698431365
transform 1 0 28000 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_350
timestamp 1698431365
transform 1 0 31808 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_351
timestamp 1698431365
transform 1 0 35616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_352
timestamp 1698431365
transform 1 0 39424 0 1 40768
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 31136 800 31248 0 FreeSans 448 0 0 0 RXD
port 0 nsew signal tristate
flabel metal3 s 0 29792 800 29904 0 FreeSans 448 0 0 0 TXD
port 1 nsew signal input
flabel metal3 s 0 2912 800 3024 0 FreeSans 448 0 0 0 addr[0]
port 2 nsew signal input
flabel metal3 s 0 4256 800 4368 0 FreeSans 448 0 0 0 addr[1]
port 3 nsew signal input
flabel metal3 s 0 5600 800 5712 0 FreeSans 448 0 0 0 addr[2]
port 4 nsew signal input
flabel metal3 s 0 6944 800 7056 0 FreeSans 448 0 0 0 addr[3]
port 5 nsew signal input
flabel metal2 s 31360 0 31472 800 0 FreeSans 448 90 0 0 bus_cyc
port 6 nsew signal input
flabel metal2 s 33152 0 33264 800 0 FreeSans 448 90 0 0 bus_we
port 7 nsew signal input
flabel metal3 s 0 8288 800 8400 0 FreeSans 448 0 0 0 data_in[0]
port 8 nsew signal input
flabel metal3 s 0 9632 800 9744 0 FreeSans 448 0 0 0 data_in[1]
port 9 nsew signal input
flabel metal3 s 0 10976 800 11088 0 FreeSans 448 0 0 0 data_in[2]
port 10 nsew signal input
flabel metal3 s 0 12320 800 12432 0 FreeSans 448 0 0 0 data_in[3]
port 11 nsew signal input
flabel metal3 s 0 13664 800 13776 0 FreeSans 448 0 0 0 data_in[4]
port 12 nsew signal input
flabel metal3 s 0 15008 800 15120 0 FreeSans 448 0 0 0 data_in[5]
port 13 nsew signal input
flabel metal3 s 0 16352 800 16464 0 FreeSans 448 0 0 0 data_in[6]
port 14 nsew signal input
flabel metal3 s 0 17696 800 17808 0 FreeSans 448 0 0 0 data_in[7]
port 15 nsew signal input
flabel metal3 s 0 19040 800 19152 0 FreeSans 448 0 0 0 data_out[0]
port 16 nsew signal tristate
flabel metal3 s 0 20384 800 20496 0 FreeSans 448 0 0 0 data_out[1]
port 17 nsew signal tristate
flabel metal3 s 0 21728 800 21840 0 FreeSans 448 0 0 0 data_out[2]
port 18 nsew signal tristate
flabel metal3 s 0 23072 800 23184 0 FreeSans 448 0 0 0 data_out[3]
port 19 nsew signal tristate
flabel metal3 s 0 24416 800 24528 0 FreeSans 448 0 0 0 data_out[4]
port 20 nsew signal tristate
flabel metal3 s 0 25760 800 25872 0 FreeSans 448 0 0 0 data_out[5]
port 21 nsew signal tristate
flabel metal3 s 0 27104 800 27216 0 FreeSans 448 0 0 0 data_out[6]
port 22 nsew signal tristate
flabel metal3 s 0 28448 800 28560 0 FreeSans 448 0 0 0 data_out[7]
port 23 nsew signal tristate
flabel metal2 s 3808 44200 3920 45000 0 FreeSans 448 90 0 0 io_in[0]
port 24 nsew signal input
flabel metal2 s 15008 44200 15120 45000 0 FreeSans 448 90 0 0 io_in[10]
port 25 nsew signal input
flabel metal2 s 16128 44200 16240 45000 0 FreeSans 448 90 0 0 io_in[11]
port 26 nsew signal input
flabel metal2 s 17248 44200 17360 45000 0 FreeSans 448 90 0 0 io_in[12]
port 27 nsew signal input
flabel metal2 s 18368 44200 18480 45000 0 FreeSans 448 90 0 0 io_in[13]
port 28 nsew signal input
flabel metal2 s 19488 44200 19600 45000 0 FreeSans 448 90 0 0 io_in[14]
port 29 nsew signal input
flabel metal2 s 20608 44200 20720 45000 0 FreeSans 448 90 0 0 io_in[15]
port 30 nsew signal input
flabel metal2 s 4928 44200 5040 45000 0 FreeSans 448 90 0 0 io_in[1]
port 31 nsew signal input
flabel metal2 s 6048 44200 6160 45000 0 FreeSans 448 90 0 0 io_in[2]
port 32 nsew signal input
flabel metal2 s 7168 44200 7280 45000 0 FreeSans 448 90 0 0 io_in[3]
port 33 nsew signal input
flabel metal2 s 8288 44200 8400 45000 0 FreeSans 448 90 0 0 io_in[4]
port 34 nsew signal input
flabel metal2 s 9408 44200 9520 45000 0 FreeSans 448 90 0 0 io_in[5]
port 35 nsew signal input
flabel metal2 s 10528 44200 10640 45000 0 FreeSans 448 90 0 0 io_in[6]
port 36 nsew signal input
flabel metal2 s 11648 44200 11760 45000 0 FreeSans 448 90 0 0 io_in[7]
port 37 nsew signal input
flabel metal2 s 12768 44200 12880 45000 0 FreeSans 448 90 0 0 io_in[8]
port 38 nsew signal input
flabel metal2 s 13888 44200 14000 45000 0 FreeSans 448 90 0 0 io_in[9]
port 39 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 40 nsew signal tristate
flabel metal2 s 20608 0 20720 800 0 FreeSans 448 90 0 0 io_oeb[10]
port 41 nsew signal tristate
flabel metal2 s 22400 0 22512 800 0 FreeSans 448 90 0 0 io_oeb[11]
port 42 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 io_oeb[12]
port 43 nsew signal tristate
flabel metal2 s 25984 0 26096 800 0 FreeSans 448 90 0 0 io_oeb[13]
port 44 nsew signal tristate
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 io_oeb[14]
port 45 nsew signal tristate
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 io_oeb[15]
port 46 nsew signal tristate
flabel metal2 s 4480 0 4592 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 47 nsew signal tristate
flabel metal2 s 6272 0 6384 800 0 FreeSans 448 90 0 0 io_oeb[2]
port 48 nsew signal tristate
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 49 nsew signal tristate
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 io_oeb[4]
port 50 nsew signal tristate
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 io_oeb[5]
port 51 nsew signal tristate
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 io_oeb[6]
port 52 nsew signal tristate
flabel metal2 s 15232 0 15344 800 0 FreeSans 448 90 0 0 io_oeb[7]
port 53 nsew signal tristate
flabel metal2 s 17024 0 17136 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 54 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 55 nsew signal tristate
flabel metal2 s 21728 44200 21840 45000 0 FreeSans 448 90 0 0 io_out[0]
port 56 nsew signal tristate
flabel metal2 s 32928 44200 33040 45000 0 FreeSans 448 90 0 0 io_out[10]
port 57 nsew signal tristate
flabel metal2 s 34048 44200 34160 45000 0 FreeSans 448 90 0 0 io_out[11]
port 58 nsew signal tristate
flabel metal2 s 35168 44200 35280 45000 0 FreeSans 448 90 0 0 io_out[12]
port 59 nsew signal tristate
flabel metal2 s 36288 44200 36400 45000 0 FreeSans 448 90 0 0 io_out[13]
port 60 nsew signal tristate
flabel metal2 s 37408 44200 37520 45000 0 FreeSans 448 90 0 0 io_out[14]
port 61 nsew signal tristate
flabel metal2 s 38528 44200 38640 45000 0 FreeSans 448 90 0 0 io_out[15]
port 62 nsew signal tristate
flabel metal2 s 22848 44200 22960 45000 0 FreeSans 448 90 0 0 io_out[1]
port 63 nsew signal tristate
flabel metal2 s 23968 44200 24080 45000 0 FreeSans 448 90 0 0 io_out[2]
port 64 nsew signal tristate
flabel metal2 s 25088 44200 25200 45000 0 FreeSans 448 90 0 0 io_out[3]
port 65 nsew signal tristate
flabel metal2 s 26208 44200 26320 45000 0 FreeSans 448 90 0 0 io_out[4]
port 66 nsew signal tristate
flabel metal2 s 27328 44200 27440 45000 0 FreeSans 448 90 0 0 io_out[5]
port 67 nsew signal tristate
flabel metal2 s 28448 44200 28560 45000 0 FreeSans 448 90 0 0 io_out[6]
port 68 nsew signal tristate
flabel metal2 s 29568 44200 29680 45000 0 FreeSans 448 90 0 0 io_out[7]
port 69 nsew signal tristate
flabel metal2 s 30688 44200 30800 45000 0 FreeSans 448 90 0 0 io_out[8]
port 70 nsew signal tristate
flabel metal2 s 31808 44200 31920 45000 0 FreeSans 448 90 0 0 io_out[9]
port 71 nsew signal tristate
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 irq0
port 72 nsew signal tristate
flabel metal2 s 36736 0 36848 800 0 FreeSans 448 90 0 0 irq6
port 73 nsew signal tristate
flabel metal2 s 38528 0 38640 800 0 FreeSans 448 90 0 0 irq7
port 74 nsew signal tristate
flabel metal3 s 0 32480 800 32592 0 FreeSans 448 0 0 0 la_data_out[0]
port 75 nsew signal tristate
flabel metal3 s 0 33824 800 33936 0 FreeSans 448 0 0 0 la_data_out[1]
port 76 nsew signal tristate
flabel metal3 s 0 35168 800 35280 0 FreeSans 448 0 0 0 la_data_out[2]
port 77 nsew signal tristate
flabel metal3 s 0 36512 800 36624 0 FreeSans 448 0 0 0 la_data_out[3]
port 78 nsew signal tristate
flabel metal3 s 0 37856 800 37968 0 FreeSans 448 0 0 0 la_data_out[4]
port 79 nsew signal tristate
flabel metal3 s 0 39200 800 39312 0 FreeSans 448 0 0 0 la_data_out[5]
port 80 nsew signal tristate
flabel metal3 s 0 40544 800 40656 0 FreeSans 448 0 0 0 la_data_out[6]
port 81 nsew signal tristate
flabel metal3 s 0 41888 800 42000 0 FreeSans 448 0 0 0 la_data_out[7]
port 82 nsew signal tristate
flabel metal3 s 44200 22400 45000 22512 0 FreeSans 448 0 0 0 pwm0
port 83 nsew signal input
flabel metal3 s 44200 31360 45000 31472 0 FreeSans 448 0 0 0 pwm1
port 84 nsew signal input
flabel metal3 s 44200 40320 45000 40432 0 FreeSans 448 0 0 0 pwm2
port 85 nsew signal input
flabel metal2 s 42112 0 42224 800 0 FreeSans 448 90 0 0 rst
port 86 nsew signal input
flabel metal2 s 39648 44200 39760 45000 0 FreeSans 448 90 0 0 tmr0_clk
port 87 nsew signal tristate
flabel metal3 s 44200 4480 45000 4592 0 FreeSans 448 0 0 0 tmr0_o
port 88 nsew signal input
flabel metal2 s 40768 44200 40880 45000 0 FreeSans 448 90 0 0 tmr1_clk
port 89 nsew signal tristate
flabel metal3 s 44200 13440 45000 13552 0 FreeSans 448 0 0 0 tmr1_o
port 90 nsew signal input
flabel metal4 s 4448 3076 4768 41612 0 FreeSans 1280 90 0 0 vdd
port 91 nsew power bidirectional
flabel metal4 s 35168 3076 35488 41612 0 FreeSans 1280 90 0 0 vdd
port 91 nsew power bidirectional
flabel metal4 s 19808 3076 20128 41612 0 FreeSans 1280 90 0 0 vss
port 92 nsew ground bidirectional
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 wb_clk_i
port 93 nsew signal input
rlabel metal1 22456 41552 22456 41552 0 vdd
rlabel metal1 22456 40768 22456 40768 0 vss
rlabel metal2 5096 11592 5096 11592 0 DDRA\[0\]
rlabel metal2 10472 11704 10472 11704 0 DDRA\[1\]
rlabel metal3 3584 13048 3584 13048 0 DDRA\[2\]
rlabel metal2 13720 12320 13720 12320 0 DDRA\[3\]
rlabel metal2 11928 6776 11928 6776 0 DDRA\[4\]
rlabel metal2 13048 8008 13048 8008 0 DDRA\[5\]
rlabel metal3 11144 7672 11144 7672 0 DDRA\[6\]
rlabel metal3 13272 6552 13272 6552 0 DDRA\[7\]
rlabel metal2 17864 21224 17864 21224 0 DDRB\[0\]
rlabel metal2 16744 12656 16744 12656 0 DDRB\[1\]
rlabel metal2 20776 22568 20776 22568 0 DDRB\[2\]
rlabel metal2 21224 9968 21224 9968 0 DDRB\[3\]
rlabel metal2 25368 21616 25368 21616 0 DDRB\[4\]
rlabel metal2 16632 16968 16632 16968 0 DDRB\[5\]
rlabel metal3 28168 9744 28168 9744 0 DDRB\[6\]
rlabel metal2 29624 9352 29624 9352 0 DDRB\[7\]
rlabel metal3 15512 37912 15512 37912 0 PORTA\[0\]
rlabel metal3 17192 37800 17192 37800 0 PORTA\[1\]
rlabel metal3 12880 39704 12880 39704 0 PORTA\[2\]
rlabel metal3 22736 38136 22736 38136 0 PORTA\[3\]
rlabel metal2 28616 36232 28616 36232 0 PORTA\[4\]
rlabel metal2 28504 34832 28504 34832 0 PORTA\[5\]
rlabel metal2 31752 35896 31752 35896 0 PORTA\[6\]
rlabel metal3 22456 36344 22456 36344 0 PORTA\[7\]
rlabel metal2 19656 25760 19656 25760 0 PORTB\[0\]
rlabel metal2 29176 37968 29176 37968 0 PORTB\[1\]
rlabel metal3 25144 27160 25144 27160 0 PORTB\[2\]
rlabel metal2 20328 31696 20328 31696 0 PORTB\[3\]
rlabel metal2 27944 27832 27944 27832 0 PORTB\[4\]
rlabel metal2 27720 31360 27720 31360 0 PORTB\[5\]
rlabel metal2 30856 28280 30856 28280 0 PORTB\[6\]
rlabel metal2 29288 29792 29288 29792 0 PORTB\[7\]
rlabel metal3 1358 31192 1358 31192 0 RXD
rlabel metal2 15064 22064 15064 22064 0 SPA\[0\]
rlabel metal2 11928 14000 11928 14000 0 SPA\[1\]
rlabel metal2 16968 33320 16968 33320 0 SPA\[2\]
rlabel metal2 14728 12824 14728 12824 0 SPA\[3\]
rlabel metal2 29512 27496 29512 27496 0 SPA\[4\]
rlabel metal2 28336 30184 28336 30184 0 SPA\[5\]
rlabel metal2 29736 14672 29736 14672 0 SPA\[6\]
rlabel metal2 10248 33040 10248 33040 0 SPA\[7\]
rlabel metal2 17640 23464 17640 23464 0 SPB\[0\]
rlabel metal2 28000 30744 28000 30744 0 SPB\[1\]
rlabel metal2 23912 24976 23912 24976 0 SPB\[2\]
rlabel metal3 24640 38696 24640 38696 0 SPB\[3\]
rlabel metal2 25592 25704 25592 25704 0 SPB\[4\]
rlabel metal2 16240 16072 16240 16072 0 SPB\[5\]
rlabel metal2 31640 25536 31640 25536 0 SPB\[6\]
rlabel metal2 32760 29288 32760 29288 0 SPB\[7\]
rlabel metal2 1848 30128 1848 30128 0 TXD
rlabel metal2 34776 19656 34776 19656 0 _000_
rlabel metal2 8288 21448 8288 21448 0 _001_
rlabel metal3 7112 20888 7112 20888 0 _002_
rlabel metal2 5768 23464 5768 23464 0 _003_
rlabel metal3 5376 24024 5376 24024 0 _004_
rlabel metal2 3864 25312 3864 25312 0 _005_
rlabel metal2 5880 26432 5880 26432 0 _006_
rlabel metal2 12096 27160 12096 27160 0 _007_
rlabel metal2 8456 28504 8456 28504 0 _008_
rlabel metal2 32872 16240 32872 16240 0 _009_
rlabel metal2 33320 23464 33320 23464 0 _010_
rlabel metal2 36064 18536 36064 18536 0 _011_
rlabel metal2 5768 34440 5768 34440 0 _012_
rlabel metal2 3864 29848 3864 29848 0 _013_
rlabel metal2 2968 37632 2968 37632 0 _014_
rlabel metal2 2464 35560 2464 35560 0 _015_
rlabel metal2 9800 37688 9800 37688 0 _016_
rlabel metal2 2520 38192 2520 38192 0 _017_
rlabel metal2 9688 39256 9688 39256 0 _018_
rlabel metal3 6720 37464 6720 37464 0 _019_
rlabel metal2 6272 10808 6272 10808 0 _020_
rlabel metal2 8344 11760 8344 11760 0 _021_
rlabel metal2 3024 10696 3024 10696 0 _022_
rlabel metal2 12264 10192 12264 10192 0 _023_
rlabel metal2 8904 5824 8904 5824 0 _024_
rlabel metal2 11704 6664 11704 6664 0 _025_
rlabel metal2 7896 7336 7896 7336 0 _026_
rlabel metal2 15624 5824 15624 5824 0 _027_
rlabel metal2 15848 6832 15848 6832 0 _028_
rlabel metal2 18088 10976 18088 10976 0 _029_
rlabel metal2 18200 5712 18200 5712 0 _030_
rlabel metal2 18592 5208 18592 5208 0 _031_
rlabel metal2 22120 6328 22120 6328 0 _032_
rlabel metal3 23408 9688 23408 9688 0 _033_
rlabel metal3 24584 8904 24584 8904 0 _034_
rlabel metal2 29232 9128 29232 9128 0 _035_
rlabel metal2 14392 38696 14392 38696 0 _036_
rlabel metal2 18312 39256 18312 39256 0 _037_
rlabel metal2 15736 39256 15736 39256 0 _038_
rlabel metal2 18648 37688 18648 37688 0 _039_
rlabel metal2 24248 36288 24248 36288 0 _040_
rlabel metal2 26376 35056 26376 35056 0 _041_
rlabel metal3 26936 35560 26936 35560 0 _042_
rlabel metal2 23240 37240 23240 37240 0 _043_
rlabel metal3 22400 26152 22400 26152 0 _044_
rlabel metal3 23408 30184 23408 30184 0 _045_
rlabel metal2 22680 27440 22680 27440 0 _046_
rlabel metal2 21000 31416 21000 31416 0 _047_
rlabel metal2 27832 26712 27832 26712 0 _048_
rlabel metal2 28728 31416 28728 31416 0 _049_
rlabel metal2 33880 28168 33880 28168 0 _050_
rlabel metal3 30968 30072 30968 30072 0 _051_
rlabel metal2 15624 20552 15624 20552 0 _052_
rlabel metal2 21392 13832 21392 13832 0 _053_
rlabel metal2 21392 22008 21392 22008 0 _054_
rlabel metal2 23408 13048 23408 13048 0 _055_
rlabel metal2 27944 11144 27944 11144 0 _056_
rlabel metal2 27664 13832 27664 13832 0 _057_
rlabel metal2 30128 15400 30128 15400 0 _058_
rlabel metal2 18200 18256 18200 18256 0 _059_
rlabel metal2 21448 20328 21448 20328 0 _060_
rlabel metal3 23968 18424 23968 18424 0 _061_
rlabel metal2 23464 21392 23464 21392 0 _062_
rlabel metal2 23016 18368 23016 18368 0 _063_
rlabel metal2 27048 23352 27048 23352 0 _064_
rlabel metal2 30856 18480 30856 18480 0 _065_
rlabel metal2 29512 23576 29512 23576 0 _066_
rlabel metal2 31248 23352 31248 23352 0 _067_
rlabel metal2 31528 17528 31528 17528 0 _068_
rlabel metal2 34496 23240 34496 23240 0 _069_
rlabel metal2 5768 12880 5768 12880 0 _070_
rlabel metal3 18032 38248 18032 38248 0 _071_
rlabel metal2 21112 39480 21112 39480 0 _072_
rlabel metal3 7056 12376 7056 12376 0 _073_
rlabel metal2 16856 39256 16856 39256 0 _074_
rlabel metal2 24528 40376 24528 40376 0 _075_
rlabel metal2 28280 35560 28280 35560 0 _076_
rlabel metal2 27384 36176 27384 36176 0 _077_
rlabel metal2 30856 36568 30856 36568 0 _078_
rlabel metal2 23912 39200 23912 39200 0 _079_
rlabel metal2 25816 39256 25816 39256 0 _080_
rlabel metal2 5768 30072 5768 30072 0 _081_
rlabel metal2 20216 23408 20216 23408 0 _082_
rlabel metal2 29288 37968 29288 37968 0 _083_
rlabel metal3 30632 38808 30632 38808 0 _084_
rlabel metal2 23464 25088 23464 25088 0 _085_
rlabel metal2 31528 34860 31528 34860 0 _086_
rlabel metal2 22904 22064 22904 22064 0 _087_
rlabel metal2 33096 35280 33096 35280 0 _088_
rlabel metal2 25928 21952 25928 21952 0 _089_
rlabel metal2 29736 28168 29736 28168 0 _090_
rlabel metal2 31192 30856 31192 30856 0 _091_
rlabel metal2 31864 34944 31864 34944 0 _092_
rlabel metal2 28000 9912 28000 9912 0 _093_
rlabel metal3 35336 27272 35336 27272 0 _094_
rlabel metal2 30688 9912 30688 9912 0 _095_
rlabel metal2 35000 30856 35000 30856 0 _096_
rlabel metal2 38360 39144 38360 39144 0 _097_
rlabel metal2 24696 39088 24696 39088 0 _098_
rlabel metal3 17920 23912 17920 23912 0 _099_
rlabel metal2 17640 26320 17640 26320 0 _100_
rlabel metal2 33096 23240 33096 23240 0 _101_
rlabel metal2 13832 20384 13832 20384 0 _102_
rlabel metal2 15512 26824 15512 26824 0 _103_
rlabel metal2 10584 27664 10584 27664 0 _104_
rlabel metal2 9800 23912 9800 23912 0 _105_
rlabel metal2 11368 21896 11368 21896 0 _106_
rlabel metal2 2632 14616 2632 14616 0 _107_
rlabel metal2 3696 13832 3696 13832 0 _108_
rlabel metal2 5824 18424 5824 18424 0 _109_
rlabel metal2 3192 16464 3192 16464 0 _110_
rlabel metal2 15400 23800 15400 23800 0 _111_
rlabel metal2 16128 24696 16128 24696 0 _112_
rlabel metal2 6104 18480 6104 18480 0 _113_
rlabel metal2 10136 17192 10136 17192 0 _114_
rlabel metal2 5656 14784 5656 14784 0 _115_
rlabel metal2 7168 13720 7168 13720 0 _116_
rlabel metal2 2632 16520 2632 16520 0 _117_
rlabel metal2 7392 13832 7392 13832 0 _118_
rlabel metal2 2296 16072 2296 16072 0 _119_
rlabel metal2 16408 25480 16408 25480 0 _120_
rlabel metal2 15960 20888 15960 20888 0 _121_
rlabel metal2 7224 17640 7224 17640 0 _122_
rlabel metal2 8120 19600 8120 19600 0 _123_
rlabel metal3 10024 19992 10024 19992 0 _124_
rlabel metal2 11424 22232 11424 22232 0 _125_
rlabel metal2 6664 14756 6664 14756 0 _126_
rlabel metal2 17304 15512 17304 15512 0 _127_
rlabel metal2 10136 24528 10136 24528 0 _128_
rlabel metal2 3136 17752 3136 17752 0 _129_
rlabel metal3 16912 24920 16912 24920 0 _130_
rlabel metal2 15176 24976 15176 24976 0 _131_
rlabel metal2 5880 17192 5880 17192 0 _132_
rlabel metal2 6496 21336 6496 21336 0 _133_
rlabel metal3 11984 35336 11984 35336 0 _134_
rlabel metal3 4704 14616 4704 14616 0 _135_
rlabel metal2 17416 34384 17416 34384 0 _136_
rlabel metal2 15848 30968 15848 30968 0 _137_
rlabel metal2 17416 16296 17416 16296 0 _138_
rlabel metal2 12600 32872 12600 32872 0 _139_
rlabel metal2 12488 25536 12488 25536 0 _140_
rlabel metal2 16296 32088 16296 32088 0 _141_
rlabel metal2 11592 32368 11592 32368 0 _142_
rlabel metal3 8288 15960 8288 15960 0 _143_
rlabel metal2 11592 18200 11592 18200 0 _144_
rlabel metal2 7896 31080 7896 31080 0 _145_
rlabel metal2 12376 25592 12376 25592 0 _146_
rlabel metal2 11704 23016 11704 23016 0 _147_
rlabel metal2 18312 23352 18312 23352 0 _148_
rlabel metal3 7728 21448 7728 21448 0 _149_
rlabel metal3 8848 20664 8848 20664 0 _150_
rlabel metal2 11928 15736 11928 15736 0 _151_
rlabel metal2 11368 15512 11368 15512 0 _152_
rlabel metal2 10584 20216 10584 20216 0 _153_
rlabel metal2 15848 33600 15848 33600 0 _154_
rlabel metal2 14616 36568 14616 36568 0 _155_
rlabel metal2 9912 31024 9912 31024 0 _156_
rlabel metal2 9800 24416 9800 24416 0 _157_
rlabel metal3 9184 31080 9184 31080 0 _158_
rlabel metal2 16520 26936 16520 26936 0 _159_
rlabel metal2 17752 29736 17752 29736 0 _160_
rlabel metal2 10528 23576 10528 23576 0 _161_
rlabel metal2 8456 23632 8456 23632 0 _162_
rlabel metal2 11704 24304 11704 24304 0 _163_
rlabel metal2 10248 22904 10248 22904 0 _164_
rlabel metal2 10584 23968 10584 23968 0 _165_
rlabel metal2 6664 32032 6664 32032 0 _166_
rlabel metal2 10360 29960 10360 29960 0 _167_
rlabel metal2 10136 29680 10136 29680 0 _168_
rlabel metal2 10808 23744 10808 23744 0 _169_
rlabel metal2 10360 23856 10360 23856 0 _170_
rlabel metal2 7560 27048 7560 27048 0 _171_
rlabel metal2 5768 24360 5768 24360 0 _172_
rlabel metal2 15176 16464 15176 16464 0 _173_
rlabel metal2 7336 22848 7336 22848 0 _174_
rlabel metal2 7672 33936 7672 33936 0 _175_
rlabel metal2 10248 31640 10248 31640 0 _176_
rlabel metal3 8064 32760 8064 32760 0 _177_
rlabel metal2 6440 33208 6440 33208 0 _178_
rlabel metal2 7616 30408 7616 30408 0 _179_
rlabel metal3 6608 25592 6608 25592 0 _180_
rlabel metal3 10528 24584 10528 24584 0 _181_
rlabel metal3 11760 24696 11760 24696 0 _182_
rlabel metal3 9184 24920 9184 24920 0 _183_
rlabel metal2 12264 31528 12264 31528 0 _184_
rlabel metal3 14168 30744 14168 30744 0 _185_
rlabel metal3 9912 30296 9912 30296 0 _186_
rlabel metal2 7336 26544 7336 26544 0 _187_
rlabel metal2 15512 17360 15512 17360 0 _188_
rlabel metal2 7784 32480 7784 32480 0 _189_
rlabel metal2 9912 32200 9912 32200 0 _190_
rlabel metal2 7224 33376 7224 33376 0 _191_
rlabel metal2 7952 29624 7952 29624 0 _192_
rlabel metal3 11872 27720 11872 27720 0 _193_
rlabel metal2 13048 27384 13048 27384 0 _194_
rlabel metal3 13272 35784 13272 35784 0 _195_
rlabel metal2 15736 26992 15736 26992 0 _196_
rlabel metal2 16296 26208 16296 26208 0 _197_
rlabel metal2 15176 27552 15176 27552 0 _198_
rlabel metal2 10696 28616 10696 28616 0 _199_
rlabel metal3 20720 38696 20720 38696 0 _200_
rlabel metal2 12264 19264 12264 19264 0 _201_
rlabel metal2 12712 19264 12712 19264 0 _202_
rlabel metal3 11536 25928 11536 25928 0 _203_
rlabel metal2 14168 29680 14168 29680 0 _204_
rlabel metal2 14112 19320 14112 19320 0 _205_
rlabel metal2 17528 29792 17528 29792 0 _206_
rlabel metal3 12712 28616 12712 28616 0 _207_
rlabel metal2 23576 18480 23576 18480 0 _208_
rlabel metal2 15960 15204 15960 15204 0 _209_
rlabel metal2 16744 15288 16744 15288 0 _210_
rlabel metal2 28504 18032 28504 18032 0 _211_
rlabel metal2 31528 19936 31528 19936 0 _212_
rlabel metal2 15288 21672 15288 21672 0 _213_
rlabel metal2 32088 20160 32088 20160 0 _214_
rlabel metal2 33096 17528 33096 17528 0 _215_
rlabel metal2 28728 23912 28728 23912 0 _216_
rlabel metal2 29960 21448 29960 21448 0 _217_
rlabel metal2 34048 24472 34048 24472 0 _218_
rlabel metal2 34216 22400 34216 22400 0 _219_
rlabel metal2 33768 22680 33768 22680 0 _220_
rlabel metal3 21224 24584 21224 24584 0 _221_
rlabel metal2 29288 27944 29288 27944 0 _222_
rlabel metal3 32144 20216 32144 20216 0 _223_
rlabel metal2 36232 19376 36232 19376 0 _224_
rlabel metal2 35504 19432 35504 19432 0 _225_
rlabel metal2 7224 11200 7224 11200 0 _226_
rlabel metal2 8568 16128 8568 16128 0 _227_
rlabel metal3 12376 14728 12376 14728 0 _228_
rlabel metal2 8456 18088 8456 18088 0 _229_
rlabel metal3 9968 36456 9968 36456 0 _230_
rlabel metal2 5992 35168 5992 35168 0 _231_
rlabel metal2 6664 29232 6664 29232 0 _232_
rlabel metal2 4368 29400 4368 29400 0 _233_
rlabel metal2 2744 29568 2744 29568 0 _234_
rlabel metal2 3080 30296 3080 30296 0 _235_
rlabel metal2 4984 34104 4984 34104 0 _236_
rlabel metal2 10192 34776 10192 34776 0 _237_
rlabel metal2 3304 29344 3304 29344 0 _238_
rlabel metal2 4480 28840 4480 28840 0 _239_
rlabel metal3 6832 13048 6832 13048 0 _240_
rlabel metal3 6272 36456 6272 36456 0 _241_
rlabel metal2 7336 36680 7336 36680 0 _242_
rlabel metal2 5320 36176 5320 36176 0 _243_
rlabel metal2 2296 33264 2296 33264 0 _244_
rlabel metal2 2632 29792 2632 29792 0 _245_
rlabel metal2 21896 16800 21896 16800 0 _246_
rlabel metal3 18536 19880 18536 19880 0 _247_
rlabel metal2 11480 7616 11480 7616 0 _248_
rlabel metal2 9800 36848 9800 36848 0 _249_
rlabel metal2 8904 37352 8904 37352 0 _250_
rlabel metal2 2744 34160 2744 34160 0 _251_
rlabel metal2 3080 33432 3080 33432 0 _252_
rlabel metal2 12040 8848 12040 8848 0 _253_
rlabel metal2 10584 37072 10584 37072 0 _254_
rlabel metal3 8344 38808 8344 38808 0 _255_
rlabel metal3 10920 8120 10920 8120 0 _256_
rlabel metal2 7784 36848 7784 36848 0 _257_
rlabel metal2 7504 35896 7504 35896 0 _258_
rlabel metal2 10696 8008 10696 8008 0 _259_
rlabel metal2 8120 10808 8120 10808 0 _260_
rlabel metal2 15400 17248 15400 17248 0 _261_
rlabel metal2 11704 11648 11704 11648 0 _262_
rlabel metal2 7224 12040 7224 12040 0 _263_
rlabel metal3 6776 10584 6776 10584 0 _264_
rlabel metal2 11312 11368 11312 11368 0 _265_
rlabel metal2 6552 10080 6552 10080 0 _266_
rlabel metal2 6216 10192 6216 10192 0 _267_
rlabel metal3 10920 12376 10920 12376 0 _268_
rlabel metal2 10136 12376 10136 12376 0 _269_
rlabel metal2 9296 12152 9296 12152 0 _270_
rlabel metal2 6104 11648 6104 11648 0 _271_
rlabel metal2 5544 11088 5544 11088 0 _272_
rlabel metal2 12936 9576 12936 9576 0 _273_
rlabel metal2 12712 10024 12712 10024 0 _274_
rlabel metal2 12488 10472 12488 10472 0 _275_
rlabel metal2 10360 7392 10360 7392 0 _276_
rlabel metal3 11200 8232 11200 8232 0 _277_
rlabel metal2 10696 6888 10696 6888 0 _278_
rlabel metal2 10584 7616 10584 7616 0 _279_
rlabel metal2 11032 6552 11032 6552 0 _280_
rlabel metal2 27720 29400 27720 29400 0 _281_
rlabel metal2 12376 7504 12376 7504 0 _282_
rlabel metal2 12712 7336 12712 7336 0 _283_
rlabel metal2 10136 8568 10136 8568 0 _284_
rlabel metal3 10024 7672 10024 7672 0 _285_
rlabel metal2 13832 7336 13832 7336 0 _286_
rlabel metal2 13272 6664 13272 6664 0 _287_
rlabel metal2 14168 7056 14168 7056 0 _288_
rlabel metal3 8792 15288 8792 15288 0 _289_
rlabel metal3 11816 8344 11816 8344 0 _290_
rlabel metal2 16464 9016 16464 9016 0 _291_
rlabel metal2 16520 8120 16520 8120 0 _292_
rlabel metal2 17584 10584 17584 10584 0 _293_
rlabel metal3 17808 10808 17808 10808 0 _294_
rlabel metal2 16184 7336 16184 7336 0 _295_
rlabel metal3 17360 12152 17360 12152 0 _296_
rlabel metal2 17752 12600 17752 12600 0 _297_
rlabel metal2 17416 8624 17416 8624 0 _298_
rlabel metal2 19320 7728 19320 7728 0 _299_
rlabel metal2 18424 7560 18424 7560 0 _300_
rlabel metal2 18648 7784 18648 7784 0 _301_
rlabel metal3 21000 8232 21000 8232 0 _302_
rlabel metal3 21056 10696 21056 10696 0 _303_
rlabel metal2 21336 8792 21336 8792 0 _304_
rlabel metal2 21896 8176 21896 8176 0 _305_
rlabel metal2 22568 9856 22568 9856 0 _306_
rlabel metal2 22680 8512 22680 8512 0 _307_
rlabel metal2 23240 8624 23240 8624 0 _308_
rlabel metal2 23016 9576 23016 9576 0 _309_
rlabel metal3 22512 10584 22512 10584 0 _310_
rlabel metal2 22064 7672 22064 7672 0 _311_
rlabel metal2 17976 35000 17976 35000 0 _312_
rlabel metal2 15512 36848 15512 36848 0 _313_
rlabel metal2 14728 37296 14728 37296 0 _314_
rlabel metal3 19040 36456 19040 36456 0 _315_
rlabel metal2 16408 38080 16408 38080 0 _316_
rlabel metal2 14056 38248 14056 38248 0 _317_
rlabel metal2 24584 34720 24584 34720 0 _318_
rlabel metal3 18872 38808 18872 38808 0 _319_
rlabel metal2 18312 38136 18312 38136 0 _320_
rlabel metal3 17864 37912 17864 37912 0 _321_
rlabel metal2 15568 37464 15568 37464 0 _322_
rlabel metal2 16072 38416 16072 38416 0 _323_
rlabel metal2 18312 36848 18312 36848 0 _324_
rlabel metal3 18088 37240 18088 37240 0 _325_
rlabel metal2 22344 34496 22344 34496 0 _326_
rlabel metal2 22680 35112 22680 35112 0 _327_
rlabel metal2 23576 35280 23576 35280 0 _328_
rlabel metal2 23352 35952 23352 35952 0 _329_
rlabel metal3 24080 36456 24080 36456 0 _330_
rlabel metal2 24192 34328 24192 34328 0 _331_
rlabel metal2 24136 35168 24136 35168 0 _332_
rlabel metal3 23576 35672 23576 35672 0 _333_
rlabel metal2 23744 35448 23744 35448 0 _334_
rlabel metal2 22064 35448 22064 35448 0 _335_
rlabel metal2 23016 36344 23016 36344 0 _336_
rlabel metal3 23352 28616 23352 28616 0 _337_
rlabel metal2 21336 25424 21336 25424 0 _338_
rlabel metal3 22064 25256 22064 25256 0 _339_
rlabel metal3 23352 29400 23352 29400 0 _340_
rlabel metal2 20776 30408 20776 30408 0 _341_
rlabel metal2 20888 26544 20888 26544 0 _342_
rlabel metal2 22232 27888 22232 27888 0 _343_
rlabel metal2 20888 30576 20888 30576 0 _344_
rlabel metal2 22680 30576 22680 30576 0 _345_
rlabel metal2 21672 26180 21672 26180 0 _346_
rlabel metal2 21672 27440 21672 27440 0 _347_
rlabel metal3 20552 30408 20552 30408 0 _348_
rlabel metal2 20664 30856 20664 30856 0 _349_
rlabel metal2 29176 28448 29176 28448 0 _350_
rlabel metal2 27608 27384 27608 27384 0 _351_
rlabel metal3 29288 28504 29288 28504 0 _352_
rlabel metal2 28112 28392 28112 28392 0 _353_
rlabel metal2 27328 29960 27328 29960 0 _354_
rlabel metal3 28392 30184 28392 30184 0 _355_
rlabel metal2 28448 31080 28448 31080 0 _356_
rlabel metal2 30184 27944 30184 27944 0 _357_
rlabel metal2 30856 28784 30856 28784 0 _358_
rlabel metal2 29512 28952 29512 28952 0 _359_
rlabel metal2 29624 30184 29624 30184 0 _360_
rlabel metal3 18984 15512 18984 15512 0 _361_
rlabel metal2 16576 19096 16576 19096 0 _362_
rlabel metal3 16856 18424 16856 18424 0 _363_
rlabel metal2 16072 19600 16072 19600 0 _364_
rlabel metal2 25928 15568 25928 15568 0 _365_
rlabel metal3 22120 14504 22120 14504 0 _366_
rlabel metal2 21560 14784 21560 14784 0 _367_
rlabel metal3 20440 14504 20440 14504 0 _368_
rlabel metal2 27160 14280 27160 14280 0 _369_
rlabel metal2 19208 18424 19208 18424 0 _370_
rlabel metal2 21560 19992 21560 19992 0 _371_
rlabel metal2 23352 14560 23352 14560 0 _372_
rlabel metal2 28280 14224 28280 14224 0 _373_
rlabel metal2 23800 14392 23800 14392 0 _374_
rlabel metal2 27496 13160 27496 13160 0 _375_
rlabel metal2 26712 13328 26712 13328 0 _376_
rlabel metal3 27160 14392 27160 14392 0 _377_
rlabel metal2 27832 14392 27832 14392 0 _378_
rlabel metal2 29960 16128 29960 16128 0 _379_
rlabel metal2 28952 15568 28952 15568 0 _380_
rlabel metal3 17416 17864 17416 17864 0 _381_
rlabel metal2 24192 20776 24192 20776 0 _382_
rlabel metal3 22400 20664 22400 20664 0 _383_
rlabel metal2 24192 20104 24192 20104 0 _384_
rlabel metal2 23072 19768 23072 19768 0 _385_
rlabel metal3 22960 19096 22960 19096 0 _386_
rlabel metal2 21616 18648 21616 18648 0 _387_
rlabel metal3 23856 20776 23856 20776 0 _388_
rlabel metal2 26824 21560 26824 21560 0 _389_
rlabel metal3 23464 19432 23464 19432 0 _390_
rlabel metal3 30016 23128 30016 23128 0 _391_
rlabel metal2 28392 21784 28392 21784 0 _392_
rlabel metal2 27720 22400 27720 22400 0 _393_
rlabel metal2 27496 21168 27496 21168 0 _394_
rlabel metal2 29008 22904 29008 22904 0 _395_
rlabel metal2 29512 22736 29512 22736 0 _396_
rlabel metal2 1848 3192 1848 3192 0 addr[0]
rlabel metal2 1736 4704 1736 4704 0 addr[1]
rlabel metal2 1736 5768 1736 5768 0 addr[2]
rlabel metal2 1736 7224 1736 7224 0 addr[3]
rlabel metal2 31416 2086 31416 2086 0 bus_cyc
rlabel metal2 33600 3528 33600 3528 0 bus_we
rlabel metal2 27104 27720 27104 27720 0 clknet_0_wb_clk_i
rlabel metal2 18760 9464 18760 9464 0 clknet_3_0__leaf_wb_clk_i
rlabel metal2 6888 6664 6888 6664 0 clknet_3_1__leaf_wb_clk_i
rlabel metal3 28224 13720 28224 13720 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 25368 18088 25368 18088 0 clknet_3_3__leaf_wb_clk_i
rlabel metal2 4760 25480 4760 25480 0 clknet_3_4__leaf_wb_clk_i
rlabel metal3 5824 38808 5824 38808 0 clknet_3_5__leaf_wb_clk_i
rlabel metal2 31024 30184 31024 30184 0 clknet_3_6__leaf_wb_clk_i
rlabel metal3 28000 31864 28000 31864 0 clknet_3_7__leaf_wb_clk_i
rlabel metal3 1246 8344 1246 8344 0 data_in[0]
rlabel metal3 1246 9688 1246 9688 0 data_in[1]
rlabel metal2 1736 11592 1736 11592 0 data_in[2]
rlabel metal3 1750 12376 1750 12376 0 data_in[3]
rlabel metal2 1848 13328 1848 13328 0 data_in[4]
rlabel metal2 1736 14504 1736 14504 0 data_in[5]
rlabel metal2 2408 17416 2408 17416 0 data_in[6]
rlabel metal2 1736 18088 1736 18088 0 data_in[7]
rlabel metal3 1358 19096 1358 19096 0 data_out[0]
rlabel metal3 1358 20440 1358 20440 0 data_out[1]
rlabel metal3 1358 21784 1358 21784 0 data_out[2]
rlabel metal2 1960 22848 1960 22848 0 data_out[3]
rlabel metal3 1358 24472 1358 24472 0 data_out[4]
rlabel metal3 1414 25816 1414 25816 0 data_out[5]
rlabel metal3 1358 27160 1358 27160 0 data_out[6]
rlabel metal3 1358 28504 1358 28504 0 data_out[7]
rlabel metal3 5544 39704 5544 39704 0 io_in[0]
rlabel metal2 15064 42770 15064 42770 0 io_in[10]
rlabel metal2 16184 42714 16184 42714 0 io_in[11]
rlabel metal2 17304 42770 17304 42770 0 io_in[12]
rlabel metal2 18424 42770 18424 42770 0 io_in[13]
rlabel metal2 19544 42770 19544 42770 0 io_in[14]
rlabel metal2 20832 41160 20832 41160 0 io_in[15]
rlabel metal2 4928 41160 4928 41160 0 io_in[1]
rlabel metal2 5656 41664 5656 41664 0 io_in[2]
rlabel metal2 7560 40936 7560 40936 0 io_in[3]
rlabel metal2 8344 42378 8344 42378 0 io_in[4]
rlabel metal2 9464 42770 9464 42770 0 io_in[5]
rlabel metal3 11032 40376 11032 40376 0 io_in[6]
rlabel metal2 11256 41720 11256 41720 0 io_in[7]
rlabel metal2 12992 41160 12992 41160 0 io_in[8]
rlabel metal2 14392 41552 14392 41552 0 io_in[9]
rlabel metal2 2744 2198 2744 2198 0 io_oeb[0]
rlabel metal2 20664 2058 20664 2058 0 io_oeb[10]
rlabel metal2 22456 2030 22456 2030 0 io_oeb[11]
rlabel metal2 24248 854 24248 854 0 io_oeb[12]
rlabel metal2 26040 2058 26040 2058 0 io_oeb[13]
rlabel metal2 27832 2198 27832 2198 0 io_oeb[14]
rlabel metal2 29624 2422 29624 2422 0 io_oeb[15]
rlabel metal2 4536 854 4536 854 0 io_oeb[1]
rlabel metal2 6328 2422 6328 2422 0 io_oeb[2]
rlabel metal2 8120 2030 8120 2030 0 io_oeb[3]
rlabel metal2 9912 2198 9912 2198 0 io_oeb[4]
rlabel metal2 11704 2478 11704 2478 0 io_oeb[5]
rlabel metal2 13496 2422 13496 2422 0 io_oeb[6]
rlabel metal2 15288 2030 15288 2030 0 io_oeb[7]
rlabel metal3 17752 5656 17752 5656 0 io_oeb[8]
rlabel metal2 18872 2198 18872 2198 0 io_oeb[9]
rlabel metal2 21784 42826 21784 42826 0 io_out[0]
rlabel metal2 32984 43106 32984 43106 0 io_out[10]
rlabel metal2 34104 42658 34104 42658 0 io_out[11]
rlabel metal2 35224 42994 35224 42994 0 io_out[12]
rlabel metal2 36344 43050 36344 43050 0 io_out[13]
rlabel metal2 37464 42826 37464 42826 0 io_out[14]
rlabel metal2 38584 42042 38584 42042 0 io_out[15]
rlabel metal2 22904 42042 22904 42042 0 io_out[1]
rlabel metal2 24024 42826 24024 42826 0 io_out[2]
rlabel metal2 25144 42434 25144 42434 0 io_out[3]
rlabel metal2 26264 42826 26264 42826 0 io_out[4]
rlabel metal2 27384 42434 27384 42434 0 io_out[5]
rlabel metal3 28952 39816 28952 39816 0 io_out[6]
rlabel metal2 29624 42826 29624 42826 0 io_out[7]
rlabel metal2 30744 42378 30744 42378 0 io_out[8]
rlabel metal2 31864 42042 31864 42042 0 io_out[9]
rlabel metal2 35000 2198 35000 2198 0 irq0
rlabel metal2 36792 2422 36792 2422 0 irq6
rlabel metal2 38584 2198 38584 2198 0 irq7
rlabel metal3 1358 32536 1358 32536 0 la_data_out[0]
rlabel metal3 1358 33880 1358 33880 0 la_data_out[1]
rlabel metal3 1414 35224 1414 35224 0 la_data_out[2]
rlabel metal3 1358 36568 1358 36568 0 la_data_out[3]
rlabel metal3 1358 37912 1358 37912 0 la_data_out[4]
rlabel metal3 854 39256 854 39256 0 la_data_out[5]
rlabel metal3 1358 40600 1358 40600 0 la_data_out[6]
rlabel metal3 3094 41944 3094 41944 0 la_data_out[7]
rlabel metal2 35000 22680 35000 22680 0 last_irg6_trigger
rlabel metal2 33768 18424 33768 18424 0 last_irq0_trigger
rlabel metal2 36120 19544 36120 19544 0 last_irq7_trigger
rlabel metal3 1792 29624 1792 29624 0 net1
rlabel metal2 7056 12712 7056 12712 0 net10
rlabel metal2 2408 30184 2408 30184 0 net11
rlabel metal2 27272 28392 27272 28392 0 net12
rlabel metal2 2296 14224 2296 14224 0 net13
rlabel metal2 2744 20216 2744 20216 0 net14
rlabel metal2 2072 18368 2072 18368 0 net15
rlabel metal3 5096 38696 5096 38696 0 net16
rlabel metal2 26712 39368 26712 39368 0 net17
rlabel metal2 24360 38920 24360 38920 0 net18
rlabel metal2 17304 40936 17304 40936 0 net19
rlabel metal2 2184 6328 2184 6328 0 net2
rlabel metal2 18760 40936 18760 40936 0 net20
rlabel metal2 19544 40936 19544 40936 0 net21
rlabel metal2 20776 40656 20776 40656 0 net22
rlabel metal2 7336 32368 7336 32368 0 net23
rlabel metal3 5488 40376 5488 40376 0 net24
rlabel metal2 8120 33656 8120 33656 0 net25
rlabel metal2 9576 25844 9576 25844 0 net26
rlabel metal2 9072 40936 9072 40936 0 net27
rlabel metal3 13888 18424 13888 18424 0 net28
rlabel metal2 12768 40936 12768 40936 0 net29
rlabel metal2 2072 5208 2072 5208 0 net3
rlabel metal2 13608 40936 13608 40936 0 net30
rlabel metal2 12432 35896 12432 35896 0 net31
rlabel metal2 29288 32984 29288 32984 0 net32
rlabel metal3 37016 33880 37016 33880 0 net33
rlabel metal2 29736 39816 29736 39816 0 net34
rlabel metal2 42840 4256 42840 4256 0 net35
rlabel metal2 42840 5824 42840 5824 0 net36
rlabel metal3 29400 33432 29400 33432 0 net37
rlabel metal2 4088 31472 4088 31472 0 net38
rlabel metal2 6104 21392 6104 21392 0 net39
rlabel metal2 2072 6048 2072 6048 0 net4
rlabel metal2 1736 20944 1736 20944 0 net40
rlabel metal3 5992 23016 5992 23016 0 net41
rlabel metal2 1736 23800 1736 23800 0 net42
rlabel metal3 2548 25592 2548 25592 0 net43
rlabel metal3 5488 27048 5488 27048 0 net44
rlabel metal2 10024 27496 10024 27496 0 net45
rlabel metal2 6328 28672 6328 28672 0 net46
rlabel metal2 4872 5964 4872 5964 0 net47
rlabel metal2 21224 22232 21224 22232 0 net48
rlabel metal2 21448 4592 21448 4592 0 net49
rlabel metal2 2072 8036 2072 8036 0 net5
rlabel metal2 27160 3584 27160 3584 0 net50
rlabel metal3 29624 4312 29624 4312 0 net51
rlabel metal2 28504 6552 28504 6552 0 net52
rlabel metal2 29960 6944 29960 6944 0 net53
rlabel metal3 7252 4312 7252 4312 0 net54
rlabel metal2 6440 6356 6440 6356 0 net55
rlabel metal3 11424 3528 11424 3528 0 net56
rlabel metal2 12152 4256 12152 4256 0 net57
rlabel metal2 13048 6888 13048 6888 0 net58
rlabel metal2 14168 5096 14168 5096 0 net59
rlabel metal2 32760 8344 32760 8344 0 net6
rlabel metal2 15624 8792 15624 8792 0 net60
rlabel metal2 18368 17864 18368 17864 0 net61
rlabel metal2 19264 12824 19264 12824 0 net62
rlabel metal2 20440 39536 20440 39536 0 net63
rlabel metal2 32256 39032 32256 39032 0 net64
rlabel metal2 33432 39704 33432 39704 0 net65
rlabel metal2 31528 40376 31528 40376 0 net66
rlabel metal2 35336 39536 35336 39536 0 net67
rlabel metal2 36344 40320 36344 40320 0 net68
rlabel metal3 38640 39592 38640 39592 0 net69
rlabel metal2 33432 8456 33432 8456 0 net7
rlabel metal2 21672 39536 21672 39536 0 net70
rlabel metal2 22792 40320 22792 40320 0 net71
rlabel metal3 25032 40488 25032 40488 0 net72
rlabel metal2 27496 40320 27496 40320 0 net73
rlabel metal2 27944 39704 27944 39704 0 net74
rlabel metal2 30856 39312 30856 39312 0 net75
rlabel metal2 28280 39480 28280 39480 0 net76
rlabel metal2 29512 38976 29512 38976 0 net77
rlabel metal2 31528 39312 31528 39312 0 net78
rlabel metal2 36008 3584 36008 3584 0 net79
rlabel metal2 2072 9296 2072 9296 0 net8
rlabel metal2 37016 4424 37016 4424 0 net80
rlabel metal2 39816 3584 39816 3584 0 net81
rlabel metal2 8120 33096 8120 33096 0 net82
rlabel metal2 2632 31248 2632 31248 0 net83
rlabel metal2 8120 37296 8120 37296 0 net84
rlabel metal2 4648 36120 4648 36120 0 net85
rlabel metal2 8344 39368 8344 39368 0 net86
rlabel metal2 2072 34496 2072 34496 0 net87
rlabel metal2 11648 41160 11648 41160 0 net88
rlabel metal2 11928 40544 11928 40544 0 net89
rlabel metal2 4312 11536 4312 11536 0 net9
rlabel metal2 38696 38472 38696 38472 0 net90
rlabel metal2 39480 38304 39480 38304 0 net91
rlabel metal2 4312 41104 4312 41104 0 net92
rlabel metal2 4312 37296 4312 37296 0 net93
rlabel metal2 4312 34216 4312 34216 0 net94
rlabel metal2 4312 33264 4312 33264 0 net95
rlabel metal3 6160 38920 6160 38920 0 net96
rlabel metal2 4368 40376 4368 40376 0 net97
rlabel metal2 4088 37128 4088 37128 0 net98
rlabel metal3 7812 40376 7812 40376 0 net99
rlabel metal2 43176 22792 43176 22792 0 pwm0
rlabel metal2 43176 31528 43176 31528 0 pwm1
rlabel metal3 43722 40376 43722 40376 0 pwm2
rlabel metal2 42168 2478 42168 2478 0 rst
rlabel metal2 39704 41258 39704 41258 0 tmr0_clk
rlabel metal2 43176 4816 43176 4816 0 tmr0_o
rlabel metal2 40824 44170 40824 44170 0 tmr1_clk
rlabel metal2 43176 13608 43176 13608 0 tmr1_o
rlabel metal2 40376 10654 40376 10654 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 45000 45000
<< end >>
