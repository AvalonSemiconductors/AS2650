magic
tech gf180mcuD
magscale 1 5
timestamp 1700526329
<< obsm1 >>
rect 672 1538 99288 68238
<< metal2 >>
rect 1344 69600 1400 70000
rect 3248 69600 3304 70000
rect 5152 69600 5208 70000
rect 7056 69600 7112 70000
rect 8960 69600 9016 70000
rect 10864 69600 10920 70000
rect 12768 69600 12824 70000
rect 14672 69600 14728 70000
rect 16576 69600 16632 70000
rect 18480 69600 18536 70000
rect 20384 69600 20440 70000
rect 22288 69600 22344 70000
rect 24192 69600 24248 70000
rect 26096 69600 26152 70000
rect 28000 69600 28056 70000
rect 29904 69600 29960 70000
rect 31808 69600 31864 70000
rect 33712 69600 33768 70000
rect 35616 69600 35672 70000
rect 37520 69600 37576 70000
rect 39424 69600 39480 70000
rect 41328 69600 41384 70000
rect 43232 69600 43288 70000
rect 45136 69600 45192 70000
rect 47040 69600 47096 70000
rect 48944 69600 49000 70000
rect 50848 69600 50904 70000
rect 52752 69600 52808 70000
rect 54656 69600 54712 70000
rect 56560 69600 56616 70000
rect 58464 69600 58520 70000
rect 60368 69600 60424 70000
rect 62272 69600 62328 70000
rect 64176 69600 64232 70000
rect 66080 69600 66136 70000
rect 67984 69600 68040 70000
rect 69888 69600 69944 70000
rect 71792 69600 71848 70000
rect 73696 69600 73752 70000
rect 75600 69600 75656 70000
rect 77504 69600 77560 70000
rect 79408 69600 79464 70000
rect 81312 69600 81368 70000
rect 83216 69600 83272 70000
rect 85120 69600 85176 70000
rect 87024 69600 87080 70000
rect 88928 69600 88984 70000
rect 90832 69600 90888 70000
rect 92736 69600 92792 70000
rect 94640 69600 94696 70000
rect 96544 69600 96600 70000
rect 98448 69600 98504 70000
rect 4704 0 4760 400
rect 5600 0 5656 400
rect 6496 0 6552 400
rect 7392 0 7448 400
rect 8288 0 8344 400
rect 9184 0 9240 400
rect 10080 0 10136 400
rect 10976 0 11032 400
rect 11872 0 11928 400
rect 12768 0 12824 400
rect 13664 0 13720 400
rect 14560 0 14616 400
rect 15456 0 15512 400
rect 16352 0 16408 400
rect 17248 0 17304 400
rect 18144 0 18200 400
rect 19040 0 19096 400
rect 19936 0 19992 400
rect 20832 0 20888 400
rect 21728 0 21784 400
rect 22624 0 22680 400
rect 23520 0 23576 400
rect 24416 0 24472 400
rect 25312 0 25368 400
rect 26208 0 26264 400
rect 27104 0 27160 400
rect 28000 0 28056 400
rect 28896 0 28952 400
rect 29792 0 29848 400
rect 30688 0 30744 400
rect 31584 0 31640 400
rect 32480 0 32536 400
rect 33376 0 33432 400
rect 34272 0 34328 400
rect 35168 0 35224 400
rect 36064 0 36120 400
rect 36960 0 37016 400
rect 37856 0 37912 400
rect 38752 0 38808 400
rect 39648 0 39704 400
rect 40544 0 40600 400
rect 41440 0 41496 400
rect 42336 0 42392 400
rect 43232 0 43288 400
rect 44128 0 44184 400
rect 45024 0 45080 400
rect 45920 0 45976 400
rect 46816 0 46872 400
rect 47712 0 47768 400
rect 48608 0 48664 400
rect 49504 0 49560 400
rect 50400 0 50456 400
rect 51296 0 51352 400
rect 52192 0 52248 400
rect 53088 0 53144 400
rect 53984 0 54040 400
rect 54880 0 54936 400
rect 55776 0 55832 400
rect 56672 0 56728 400
rect 57568 0 57624 400
rect 58464 0 58520 400
rect 59360 0 59416 400
rect 60256 0 60312 400
rect 61152 0 61208 400
rect 62048 0 62104 400
rect 62944 0 63000 400
rect 63840 0 63896 400
rect 64736 0 64792 400
rect 65632 0 65688 400
rect 66528 0 66584 400
rect 67424 0 67480 400
rect 68320 0 68376 400
rect 69216 0 69272 400
rect 70112 0 70168 400
rect 71008 0 71064 400
rect 71904 0 71960 400
rect 72800 0 72856 400
rect 73696 0 73752 400
rect 74592 0 74648 400
rect 75488 0 75544 400
rect 76384 0 76440 400
rect 77280 0 77336 400
rect 78176 0 78232 400
rect 79072 0 79128 400
rect 79968 0 80024 400
rect 80864 0 80920 400
rect 81760 0 81816 400
rect 82656 0 82712 400
rect 83552 0 83608 400
rect 84448 0 84504 400
rect 85344 0 85400 400
rect 86240 0 86296 400
rect 87136 0 87192 400
rect 88032 0 88088 400
rect 88928 0 88984 400
rect 89824 0 89880 400
rect 90720 0 90776 400
rect 91616 0 91672 400
rect 92512 0 92568 400
rect 93408 0 93464 400
rect 94304 0 94360 400
rect 95200 0 95256 400
<< obsm2 >>
rect 686 69570 1314 69650
rect 1430 69570 3218 69650
rect 3334 69570 5122 69650
rect 5238 69570 7026 69650
rect 7142 69570 8930 69650
rect 9046 69570 10834 69650
rect 10950 69570 12738 69650
rect 12854 69570 14642 69650
rect 14758 69570 16546 69650
rect 16662 69570 18450 69650
rect 18566 69570 20354 69650
rect 20470 69570 22258 69650
rect 22374 69570 24162 69650
rect 24278 69570 26066 69650
rect 26182 69570 27970 69650
rect 28086 69570 29874 69650
rect 29990 69570 31778 69650
rect 31894 69570 33682 69650
rect 33798 69570 35586 69650
rect 35702 69570 37490 69650
rect 37606 69570 39394 69650
rect 39510 69570 41298 69650
rect 41414 69570 43202 69650
rect 43318 69570 45106 69650
rect 45222 69570 47010 69650
rect 47126 69570 48914 69650
rect 49030 69570 50818 69650
rect 50934 69570 52722 69650
rect 52838 69570 54626 69650
rect 54742 69570 56530 69650
rect 56646 69570 58434 69650
rect 58550 69570 60338 69650
rect 60454 69570 62242 69650
rect 62358 69570 64146 69650
rect 64262 69570 66050 69650
rect 66166 69570 67954 69650
rect 68070 69570 69858 69650
rect 69974 69570 71762 69650
rect 71878 69570 73666 69650
rect 73782 69570 75570 69650
rect 75686 69570 77474 69650
rect 77590 69570 79378 69650
rect 79494 69570 81282 69650
rect 81398 69570 83186 69650
rect 83302 69570 85090 69650
rect 85206 69570 86994 69650
rect 87110 69570 88898 69650
rect 89014 69570 90802 69650
rect 90918 69570 92706 69650
rect 92822 69570 94610 69650
rect 94726 69570 96514 69650
rect 96630 69570 98418 69650
rect 98534 69570 99386 69650
rect 686 430 99386 69570
rect 686 350 4674 430
rect 4790 350 5570 430
rect 5686 350 6466 430
rect 6582 350 7362 430
rect 7478 350 8258 430
rect 8374 350 9154 430
rect 9270 350 10050 430
rect 10166 350 10946 430
rect 11062 350 11842 430
rect 11958 350 12738 430
rect 12854 350 13634 430
rect 13750 350 14530 430
rect 14646 350 15426 430
rect 15542 350 16322 430
rect 16438 350 17218 430
rect 17334 350 18114 430
rect 18230 350 19010 430
rect 19126 350 19906 430
rect 20022 350 20802 430
rect 20918 350 21698 430
rect 21814 350 22594 430
rect 22710 350 23490 430
rect 23606 350 24386 430
rect 24502 350 25282 430
rect 25398 350 26178 430
rect 26294 350 27074 430
rect 27190 350 27970 430
rect 28086 350 28866 430
rect 28982 350 29762 430
rect 29878 350 30658 430
rect 30774 350 31554 430
rect 31670 350 32450 430
rect 32566 350 33346 430
rect 33462 350 34242 430
rect 34358 350 35138 430
rect 35254 350 36034 430
rect 36150 350 36930 430
rect 37046 350 37826 430
rect 37942 350 38722 430
rect 38838 350 39618 430
rect 39734 350 40514 430
rect 40630 350 41410 430
rect 41526 350 42306 430
rect 42422 350 43202 430
rect 43318 350 44098 430
rect 44214 350 44994 430
rect 45110 350 45890 430
rect 46006 350 46786 430
rect 46902 350 47682 430
rect 47798 350 48578 430
rect 48694 350 49474 430
rect 49590 350 50370 430
rect 50486 350 51266 430
rect 51382 350 52162 430
rect 52278 350 53058 430
rect 53174 350 53954 430
rect 54070 350 54850 430
rect 54966 350 55746 430
rect 55862 350 56642 430
rect 56758 350 57538 430
rect 57654 350 58434 430
rect 58550 350 59330 430
rect 59446 350 60226 430
rect 60342 350 61122 430
rect 61238 350 62018 430
rect 62134 350 62914 430
rect 63030 350 63810 430
rect 63926 350 64706 430
rect 64822 350 65602 430
rect 65718 350 66498 430
rect 66614 350 67394 430
rect 67510 350 68290 430
rect 68406 350 69186 430
rect 69302 350 70082 430
rect 70198 350 70978 430
rect 71094 350 71874 430
rect 71990 350 72770 430
rect 72886 350 73666 430
rect 73782 350 74562 430
rect 74678 350 75458 430
rect 75574 350 76354 430
rect 76470 350 77250 430
rect 77366 350 78146 430
rect 78262 350 79042 430
rect 79158 350 79938 430
rect 80054 350 80834 430
rect 80950 350 81730 430
rect 81846 350 82626 430
rect 82742 350 83522 430
rect 83638 350 84418 430
rect 84534 350 85314 430
rect 85430 350 86210 430
rect 86326 350 87106 430
rect 87222 350 88002 430
rect 88118 350 88898 430
rect 89014 350 89794 430
rect 89910 350 90690 430
rect 90806 350 91586 430
rect 91702 350 92482 430
rect 92598 350 93378 430
rect 93494 350 94274 430
rect 94390 350 95170 430
rect 95286 350 99386 430
<< metal3 >>
rect 99600 68992 100000 69048
rect 99600 68208 100000 68264
rect 99600 67424 100000 67480
rect 99600 66640 100000 66696
rect 99600 65856 100000 65912
rect 99600 65072 100000 65128
rect 0 64848 400 64904
rect 99600 64288 100000 64344
rect 0 64176 400 64232
rect 0 63504 400 63560
rect 99600 63504 100000 63560
rect 0 62832 400 62888
rect 99600 62720 100000 62776
rect 0 62160 400 62216
rect 99600 61936 100000 61992
rect 0 61488 400 61544
rect 99600 61152 100000 61208
rect 0 60816 400 60872
rect 99600 60368 100000 60424
rect 0 60144 400 60200
rect 99600 59584 100000 59640
rect 0 59472 400 59528
rect 0 58800 400 58856
rect 99600 58800 100000 58856
rect 0 58128 400 58184
rect 99600 58016 100000 58072
rect 0 57456 400 57512
rect 99600 57232 100000 57288
rect 0 56784 400 56840
rect 99600 56448 100000 56504
rect 0 56112 400 56168
rect 99600 55664 100000 55720
rect 0 55440 400 55496
rect 99600 54880 100000 54936
rect 0 54768 400 54824
rect 0 54096 400 54152
rect 99600 54096 100000 54152
rect 0 53424 400 53480
rect 99600 53312 100000 53368
rect 0 52752 400 52808
rect 99600 52528 100000 52584
rect 0 52080 400 52136
rect 99600 51744 100000 51800
rect 0 51408 400 51464
rect 99600 50960 100000 51016
rect 0 50736 400 50792
rect 99600 50176 100000 50232
rect 0 50064 400 50120
rect 0 49392 400 49448
rect 99600 49392 100000 49448
rect 0 48720 400 48776
rect 99600 48608 100000 48664
rect 0 48048 400 48104
rect 99600 47824 100000 47880
rect 0 47376 400 47432
rect 99600 47040 100000 47096
rect 0 46704 400 46760
rect 99600 46256 100000 46312
rect 0 46032 400 46088
rect 99600 45472 100000 45528
rect 0 45360 400 45416
rect 0 44688 400 44744
rect 99600 44688 100000 44744
rect 0 44016 400 44072
rect 99600 43904 100000 43960
rect 0 43344 400 43400
rect 99600 43120 100000 43176
rect 0 42672 400 42728
rect 99600 42336 100000 42392
rect 0 42000 400 42056
rect 99600 41552 100000 41608
rect 0 41328 400 41384
rect 99600 40768 100000 40824
rect 0 40656 400 40712
rect 0 39984 400 40040
rect 99600 39984 100000 40040
rect 0 39312 400 39368
rect 99600 39200 100000 39256
rect 0 38640 400 38696
rect 99600 38416 100000 38472
rect 0 37968 400 38024
rect 99600 37632 100000 37688
rect 0 37296 400 37352
rect 99600 36848 100000 36904
rect 0 36624 400 36680
rect 99600 36064 100000 36120
rect 0 35952 400 36008
rect 0 35280 400 35336
rect 99600 35280 100000 35336
rect 0 34608 400 34664
rect 99600 34496 100000 34552
rect 0 33936 400 33992
rect 99600 33712 100000 33768
rect 0 33264 400 33320
rect 99600 32928 100000 32984
rect 0 32592 400 32648
rect 99600 32144 100000 32200
rect 0 31920 400 31976
rect 99600 31360 100000 31416
rect 0 31248 400 31304
rect 0 30576 400 30632
rect 99600 30576 100000 30632
rect 0 29904 400 29960
rect 99600 29792 100000 29848
rect 0 29232 400 29288
rect 99600 29008 100000 29064
rect 0 28560 400 28616
rect 99600 28224 100000 28280
rect 0 27888 400 27944
rect 99600 27440 100000 27496
rect 0 27216 400 27272
rect 99600 26656 100000 26712
rect 0 26544 400 26600
rect 0 25872 400 25928
rect 99600 25872 100000 25928
rect 0 25200 400 25256
rect 99600 25088 100000 25144
rect 0 24528 400 24584
rect 99600 24304 100000 24360
rect 0 23856 400 23912
rect 99600 23520 100000 23576
rect 0 23184 400 23240
rect 99600 22736 100000 22792
rect 0 22512 400 22568
rect 99600 21952 100000 22008
rect 0 21840 400 21896
rect 0 21168 400 21224
rect 99600 21168 100000 21224
rect 0 20496 400 20552
rect 99600 20384 100000 20440
rect 0 19824 400 19880
rect 99600 19600 100000 19656
rect 0 19152 400 19208
rect 99600 18816 100000 18872
rect 0 18480 400 18536
rect 99600 18032 100000 18088
rect 0 17808 400 17864
rect 99600 17248 100000 17304
rect 0 17136 400 17192
rect 0 16464 400 16520
rect 99600 16464 100000 16520
rect 0 15792 400 15848
rect 99600 15680 100000 15736
rect 0 15120 400 15176
rect 99600 14896 100000 14952
rect 0 14448 400 14504
rect 99600 14112 100000 14168
rect 0 13776 400 13832
rect 99600 13328 100000 13384
rect 0 13104 400 13160
rect 99600 12544 100000 12600
rect 0 12432 400 12488
rect 0 11760 400 11816
rect 99600 11760 100000 11816
rect 0 11088 400 11144
rect 99600 10976 100000 11032
rect 0 10416 400 10472
rect 99600 10192 100000 10248
rect 0 9744 400 9800
rect 99600 9408 100000 9464
rect 0 9072 400 9128
rect 99600 8624 100000 8680
rect 0 8400 400 8456
rect 99600 7840 100000 7896
rect 0 7728 400 7784
rect 0 7056 400 7112
rect 99600 7056 100000 7112
rect 0 6384 400 6440
rect 99600 6272 100000 6328
rect 0 5712 400 5768
rect 99600 5488 100000 5544
rect 0 5040 400 5096
rect 99600 4704 100000 4760
rect 99600 3920 100000 3976
rect 99600 3136 100000 3192
rect 99600 2352 100000 2408
rect 99600 1568 100000 1624
rect 99600 784 100000 840
<< obsm3 >>
rect 400 68962 99570 69034
rect 400 68294 99600 68962
rect 400 68178 99570 68294
rect 400 67510 99600 68178
rect 400 67394 99570 67510
rect 400 66726 99600 67394
rect 400 66610 99570 66726
rect 400 65942 99600 66610
rect 400 65826 99570 65942
rect 400 65158 99600 65826
rect 400 65042 99570 65158
rect 400 64934 99600 65042
rect 430 64818 99600 64934
rect 400 64374 99600 64818
rect 400 64262 99570 64374
rect 430 64258 99570 64262
rect 430 64146 99600 64258
rect 400 63590 99600 64146
rect 430 63474 99570 63590
rect 400 62918 99600 63474
rect 430 62806 99600 62918
rect 430 62802 99570 62806
rect 400 62690 99570 62802
rect 400 62246 99600 62690
rect 430 62130 99600 62246
rect 400 62022 99600 62130
rect 400 61906 99570 62022
rect 400 61574 99600 61906
rect 430 61458 99600 61574
rect 400 61238 99600 61458
rect 400 61122 99570 61238
rect 400 60902 99600 61122
rect 430 60786 99600 60902
rect 400 60454 99600 60786
rect 400 60338 99570 60454
rect 400 60230 99600 60338
rect 430 60114 99600 60230
rect 400 59670 99600 60114
rect 400 59558 99570 59670
rect 430 59554 99570 59558
rect 430 59442 99600 59554
rect 400 58886 99600 59442
rect 430 58770 99570 58886
rect 400 58214 99600 58770
rect 430 58102 99600 58214
rect 430 58098 99570 58102
rect 400 57986 99570 58098
rect 400 57542 99600 57986
rect 430 57426 99600 57542
rect 400 57318 99600 57426
rect 400 57202 99570 57318
rect 400 56870 99600 57202
rect 430 56754 99600 56870
rect 400 56534 99600 56754
rect 400 56418 99570 56534
rect 400 56198 99600 56418
rect 430 56082 99600 56198
rect 400 55750 99600 56082
rect 400 55634 99570 55750
rect 400 55526 99600 55634
rect 430 55410 99600 55526
rect 400 54966 99600 55410
rect 400 54854 99570 54966
rect 430 54850 99570 54854
rect 430 54738 99600 54850
rect 400 54182 99600 54738
rect 430 54066 99570 54182
rect 400 53510 99600 54066
rect 430 53398 99600 53510
rect 430 53394 99570 53398
rect 400 53282 99570 53394
rect 400 52838 99600 53282
rect 430 52722 99600 52838
rect 400 52614 99600 52722
rect 400 52498 99570 52614
rect 400 52166 99600 52498
rect 430 52050 99600 52166
rect 400 51830 99600 52050
rect 400 51714 99570 51830
rect 400 51494 99600 51714
rect 430 51378 99600 51494
rect 400 51046 99600 51378
rect 400 50930 99570 51046
rect 400 50822 99600 50930
rect 430 50706 99600 50822
rect 400 50262 99600 50706
rect 400 50150 99570 50262
rect 430 50146 99570 50150
rect 430 50034 99600 50146
rect 400 49478 99600 50034
rect 430 49362 99570 49478
rect 400 48806 99600 49362
rect 430 48694 99600 48806
rect 430 48690 99570 48694
rect 400 48578 99570 48690
rect 400 48134 99600 48578
rect 430 48018 99600 48134
rect 400 47910 99600 48018
rect 400 47794 99570 47910
rect 400 47462 99600 47794
rect 430 47346 99600 47462
rect 400 47126 99600 47346
rect 400 47010 99570 47126
rect 400 46790 99600 47010
rect 430 46674 99600 46790
rect 400 46342 99600 46674
rect 400 46226 99570 46342
rect 400 46118 99600 46226
rect 430 46002 99600 46118
rect 400 45558 99600 46002
rect 400 45446 99570 45558
rect 430 45442 99570 45446
rect 430 45330 99600 45442
rect 400 44774 99600 45330
rect 430 44658 99570 44774
rect 400 44102 99600 44658
rect 430 43990 99600 44102
rect 430 43986 99570 43990
rect 400 43874 99570 43986
rect 400 43430 99600 43874
rect 430 43314 99600 43430
rect 400 43206 99600 43314
rect 400 43090 99570 43206
rect 400 42758 99600 43090
rect 430 42642 99600 42758
rect 400 42422 99600 42642
rect 400 42306 99570 42422
rect 400 42086 99600 42306
rect 430 41970 99600 42086
rect 400 41638 99600 41970
rect 400 41522 99570 41638
rect 400 41414 99600 41522
rect 430 41298 99600 41414
rect 400 40854 99600 41298
rect 400 40742 99570 40854
rect 430 40738 99570 40742
rect 430 40626 99600 40738
rect 400 40070 99600 40626
rect 430 39954 99570 40070
rect 400 39398 99600 39954
rect 430 39286 99600 39398
rect 430 39282 99570 39286
rect 400 39170 99570 39282
rect 400 38726 99600 39170
rect 430 38610 99600 38726
rect 400 38502 99600 38610
rect 400 38386 99570 38502
rect 400 38054 99600 38386
rect 430 37938 99600 38054
rect 400 37718 99600 37938
rect 400 37602 99570 37718
rect 400 37382 99600 37602
rect 430 37266 99600 37382
rect 400 36934 99600 37266
rect 400 36818 99570 36934
rect 400 36710 99600 36818
rect 430 36594 99600 36710
rect 400 36150 99600 36594
rect 400 36038 99570 36150
rect 430 36034 99570 36038
rect 430 35922 99600 36034
rect 400 35366 99600 35922
rect 430 35250 99570 35366
rect 400 34694 99600 35250
rect 430 34582 99600 34694
rect 430 34578 99570 34582
rect 400 34466 99570 34578
rect 400 34022 99600 34466
rect 430 33906 99600 34022
rect 400 33798 99600 33906
rect 400 33682 99570 33798
rect 400 33350 99600 33682
rect 430 33234 99600 33350
rect 400 33014 99600 33234
rect 400 32898 99570 33014
rect 400 32678 99600 32898
rect 430 32562 99600 32678
rect 400 32230 99600 32562
rect 400 32114 99570 32230
rect 400 32006 99600 32114
rect 430 31890 99600 32006
rect 400 31446 99600 31890
rect 400 31334 99570 31446
rect 430 31330 99570 31334
rect 430 31218 99600 31330
rect 400 30662 99600 31218
rect 430 30546 99570 30662
rect 400 29990 99600 30546
rect 430 29878 99600 29990
rect 430 29874 99570 29878
rect 400 29762 99570 29874
rect 400 29318 99600 29762
rect 430 29202 99600 29318
rect 400 29094 99600 29202
rect 400 28978 99570 29094
rect 400 28646 99600 28978
rect 430 28530 99600 28646
rect 400 28310 99600 28530
rect 400 28194 99570 28310
rect 400 27974 99600 28194
rect 430 27858 99600 27974
rect 400 27526 99600 27858
rect 400 27410 99570 27526
rect 400 27302 99600 27410
rect 430 27186 99600 27302
rect 400 26742 99600 27186
rect 400 26630 99570 26742
rect 430 26626 99570 26630
rect 430 26514 99600 26626
rect 400 25958 99600 26514
rect 430 25842 99570 25958
rect 400 25286 99600 25842
rect 430 25174 99600 25286
rect 430 25170 99570 25174
rect 400 25058 99570 25170
rect 400 24614 99600 25058
rect 430 24498 99600 24614
rect 400 24390 99600 24498
rect 400 24274 99570 24390
rect 400 23942 99600 24274
rect 430 23826 99600 23942
rect 400 23606 99600 23826
rect 400 23490 99570 23606
rect 400 23270 99600 23490
rect 430 23154 99600 23270
rect 400 22822 99600 23154
rect 400 22706 99570 22822
rect 400 22598 99600 22706
rect 430 22482 99600 22598
rect 400 22038 99600 22482
rect 400 21926 99570 22038
rect 430 21922 99570 21926
rect 430 21810 99600 21922
rect 400 21254 99600 21810
rect 430 21138 99570 21254
rect 400 20582 99600 21138
rect 430 20470 99600 20582
rect 430 20466 99570 20470
rect 400 20354 99570 20466
rect 400 19910 99600 20354
rect 430 19794 99600 19910
rect 400 19686 99600 19794
rect 400 19570 99570 19686
rect 400 19238 99600 19570
rect 430 19122 99600 19238
rect 400 18902 99600 19122
rect 400 18786 99570 18902
rect 400 18566 99600 18786
rect 430 18450 99600 18566
rect 400 18118 99600 18450
rect 400 18002 99570 18118
rect 400 17894 99600 18002
rect 430 17778 99600 17894
rect 400 17334 99600 17778
rect 400 17222 99570 17334
rect 430 17218 99570 17222
rect 430 17106 99600 17218
rect 400 16550 99600 17106
rect 430 16434 99570 16550
rect 400 15878 99600 16434
rect 430 15766 99600 15878
rect 430 15762 99570 15766
rect 400 15650 99570 15762
rect 400 15206 99600 15650
rect 430 15090 99600 15206
rect 400 14982 99600 15090
rect 400 14866 99570 14982
rect 400 14534 99600 14866
rect 430 14418 99600 14534
rect 400 14198 99600 14418
rect 400 14082 99570 14198
rect 400 13862 99600 14082
rect 430 13746 99600 13862
rect 400 13414 99600 13746
rect 400 13298 99570 13414
rect 400 13190 99600 13298
rect 430 13074 99600 13190
rect 400 12630 99600 13074
rect 400 12518 99570 12630
rect 430 12514 99570 12518
rect 430 12402 99600 12514
rect 400 11846 99600 12402
rect 430 11730 99570 11846
rect 400 11174 99600 11730
rect 430 11062 99600 11174
rect 430 11058 99570 11062
rect 400 10946 99570 11058
rect 400 10502 99600 10946
rect 430 10386 99600 10502
rect 400 10278 99600 10386
rect 400 10162 99570 10278
rect 400 9830 99600 10162
rect 430 9714 99600 9830
rect 400 9494 99600 9714
rect 400 9378 99570 9494
rect 400 9158 99600 9378
rect 430 9042 99600 9158
rect 400 8710 99600 9042
rect 400 8594 99570 8710
rect 400 8486 99600 8594
rect 430 8370 99600 8486
rect 400 7926 99600 8370
rect 400 7814 99570 7926
rect 430 7810 99570 7814
rect 430 7698 99600 7810
rect 400 7142 99600 7698
rect 430 7026 99570 7142
rect 400 6470 99600 7026
rect 430 6358 99600 6470
rect 430 6354 99570 6358
rect 400 6242 99570 6354
rect 400 5798 99600 6242
rect 430 5682 99600 5798
rect 400 5574 99600 5682
rect 400 5458 99570 5574
rect 400 5126 99600 5458
rect 430 5010 99600 5126
rect 400 4790 99600 5010
rect 400 4674 99570 4790
rect 400 4006 99600 4674
rect 400 3890 99570 4006
rect 400 3222 99600 3890
rect 400 3106 99570 3222
rect 400 2438 99600 3106
rect 400 2322 99570 2438
rect 400 1654 99600 2322
rect 400 1538 99570 1654
rect 400 870 99600 1538
rect 400 798 99570 870
<< metal4 >>
rect 2224 1538 2384 68238
rect 9904 1538 10064 68238
rect 17584 1538 17744 68238
rect 25264 1538 25424 68238
rect 32944 1538 33104 68238
rect 40624 1538 40784 68238
rect 48304 1538 48464 68238
rect 55984 1538 56144 68238
rect 63664 1538 63824 68238
rect 71344 1538 71504 68238
rect 79024 1538 79184 68238
rect 86704 1538 86864 68238
rect 94384 1538 94544 68238
<< obsm4 >>
rect 15638 2641 17554 65175
rect 17774 2641 25234 65175
rect 25454 2641 32914 65175
rect 33134 2641 40594 65175
rect 40814 2641 48274 65175
rect 48494 2641 55954 65175
rect 56174 2641 63634 65175
rect 63854 2641 71314 65175
rect 71534 2641 78994 65175
rect 79214 2641 86674 65175
rect 86894 2641 94354 65175
rect 94574 2641 98938 65175
<< labels >>
rlabel metal3 s 0 44016 400 44072 6 RAM_end_addr[0]
port 1 nsew signal output
rlabel metal3 s 0 50736 400 50792 6 RAM_end_addr[10]
port 2 nsew signal output
rlabel metal3 s 0 51408 400 51464 6 RAM_end_addr[11]
port 3 nsew signal output
rlabel metal3 s 0 52080 400 52136 6 RAM_end_addr[12]
port 4 nsew signal output
rlabel metal3 s 0 52752 400 52808 6 RAM_end_addr[13]
port 5 nsew signal output
rlabel metal3 s 0 53424 400 53480 6 RAM_end_addr[14]
port 6 nsew signal output
rlabel metal3 s 0 54096 400 54152 6 RAM_end_addr[15]
port 7 nsew signal output
rlabel metal3 s 0 44688 400 44744 6 RAM_end_addr[1]
port 8 nsew signal output
rlabel metal3 s 0 45360 400 45416 6 RAM_end_addr[2]
port 9 nsew signal output
rlabel metal3 s 0 46032 400 46088 6 RAM_end_addr[3]
port 10 nsew signal output
rlabel metal3 s 0 46704 400 46760 6 RAM_end_addr[4]
port 11 nsew signal output
rlabel metal3 s 0 47376 400 47432 6 RAM_end_addr[5]
port 12 nsew signal output
rlabel metal3 s 0 48048 400 48104 6 RAM_end_addr[6]
port 13 nsew signal output
rlabel metal3 s 0 48720 400 48776 6 RAM_end_addr[7]
port 14 nsew signal output
rlabel metal3 s 0 49392 400 49448 6 RAM_end_addr[8]
port 15 nsew signal output
rlabel metal3 s 0 50064 400 50120 6 RAM_end_addr[9]
port 16 nsew signal output
rlabel metal3 s 0 30576 400 30632 6 RAM_start_addr[0]
port 17 nsew signal output
rlabel metal3 s 0 37296 400 37352 6 RAM_start_addr[10]
port 18 nsew signal output
rlabel metal3 s 0 37968 400 38024 6 RAM_start_addr[11]
port 19 nsew signal output
rlabel metal3 s 0 38640 400 38696 6 RAM_start_addr[12]
port 20 nsew signal output
rlabel metal3 s 0 39312 400 39368 6 RAM_start_addr[13]
port 21 nsew signal output
rlabel metal3 s 0 39984 400 40040 6 RAM_start_addr[14]
port 22 nsew signal output
rlabel metal3 s 0 40656 400 40712 6 RAM_start_addr[15]
port 23 nsew signal output
rlabel metal3 s 0 31248 400 31304 6 RAM_start_addr[1]
port 24 nsew signal output
rlabel metal3 s 0 31920 400 31976 6 RAM_start_addr[2]
port 25 nsew signal output
rlabel metal3 s 0 32592 400 32648 6 RAM_start_addr[3]
port 26 nsew signal output
rlabel metal3 s 0 33264 400 33320 6 RAM_start_addr[4]
port 27 nsew signal output
rlabel metal3 s 0 33936 400 33992 6 RAM_start_addr[5]
port 28 nsew signal output
rlabel metal3 s 0 34608 400 34664 6 RAM_start_addr[6]
port 29 nsew signal output
rlabel metal3 s 0 35280 400 35336 6 RAM_start_addr[7]
port 30 nsew signal output
rlabel metal3 s 0 35952 400 36008 6 RAM_start_addr[8]
port 31 nsew signal output
rlabel metal3 s 0 36624 400 36680 6 RAM_start_addr[9]
port 32 nsew signal output
rlabel metal2 s 94640 69600 94696 70000 6 WEb_raw
port 33 nsew signal output
rlabel metal3 s 0 43344 400 43400 6 boot_rom_en
port 34 nsew signal output
rlabel metal2 s 67984 69600 68040 70000 6 bus_addr[0]
port 35 nsew signal output
rlabel metal2 s 69888 69600 69944 70000 6 bus_addr[1]
port 36 nsew signal output
rlabel metal2 s 71792 69600 71848 70000 6 bus_addr[2]
port 37 nsew signal output
rlabel metal2 s 73696 69600 73752 70000 6 bus_addr[3]
port 38 nsew signal output
rlabel metal2 s 75600 69600 75656 70000 6 bus_addr[4]
port 39 nsew signal output
rlabel metal2 s 77504 69600 77560 70000 6 bus_addr[5]
port 40 nsew signal output
rlabel metal2 s 66080 69600 66136 70000 6 bus_cyc
port 41 nsew signal output
rlabel metal2 s 50848 69600 50904 70000 6 bus_data_out[0]
port 42 nsew signal output
rlabel metal2 s 52752 69600 52808 70000 6 bus_data_out[1]
port 43 nsew signal output
rlabel metal2 s 54656 69600 54712 70000 6 bus_data_out[2]
port 44 nsew signal output
rlabel metal2 s 56560 69600 56616 70000 6 bus_data_out[3]
port 45 nsew signal output
rlabel metal2 s 58464 69600 58520 70000 6 bus_data_out[4]
port 46 nsew signal output
rlabel metal2 s 60368 69600 60424 70000 6 bus_data_out[5]
port 47 nsew signal output
rlabel metal2 s 62272 69600 62328 70000 6 bus_data_out[6]
port 48 nsew signal output
rlabel metal2 s 64176 69600 64232 70000 6 bus_data_out[7]
port 49 nsew signal output
rlabel metal3 s 99600 47824 100000 47880 6 bus_in_gpios[0]
port 50 nsew signal input
rlabel metal3 s 99600 48608 100000 48664 6 bus_in_gpios[1]
port 51 nsew signal input
rlabel metal3 s 99600 49392 100000 49448 6 bus_in_gpios[2]
port 52 nsew signal input
rlabel metal3 s 99600 50176 100000 50232 6 bus_in_gpios[3]
port 53 nsew signal input
rlabel metal3 s 99600 50960 100000 51016 6 bus_in_gpios[4]
port 54 nsew signal input
rlabel metal3 s 99600 51744 100000 51800 6 bus_in_gpios[5]
port 55 nsew signal input
rlabel metal3 s 99600 52528 100000 52584 6 bus_in_gpios[6]
port 56 nsew signal input
rlabel metal3 s 99600 53312 100000 53368 6 bus_in_gpios[7]
port 57 nsew signal input
rlabel metal2 s 79408 69600 79464 70000 6 bus_in_serial_ports[0]
port 58 nsew signal input
rlabel metal2 s 81312 69600 81368 70000 6 bus_in_serial_ports[1]
port 59 nsew signal input
rlabel metal2 s 83216 69600 83272 70000 6 bus_in_serial_ports[2]
port 60 nsew signal input
rlabel metal2 s 85120 69600 85176 70000 6 bus_in_serial_ports[3]
port 61 nsew signal input
rlabel metal2 s 87024 69600 87080 70000 6 bus_in_serial_ports[4]
port 62 nsew signal input
rlabel metal2 s 88928 69600 88984 70000 6 bus_in_serial_ports[5]
port 63 nsew signal input
rlabel metal2 s 90832 69600 90888 70000 6 bus_in_serial_ports[6]
port 64 nsew signal input
rlabel metal2 s 92736 69600 92792 70000 6 bus_in_serial_ports[7]
port 65 nsew signal input
rlabel metal3 s 99600 63504 100000 63560 6 bus_in_sid[0]
port 66 nsew signal input
rlabel metal3 s 99600 64288 100000 64344 6 bus_in_sid[1]
port 67 nsew signal input
rlabel metal3 s 99600 65072 100000 65128 6 bus_in_sid[2]
port 68 nsew signal input
rlabel metal3 s 99600 65856 100000 65912 6 bus_in_sid[3]
port 69 nsew signal input
rlabel metal3 s 99600 66640 100000 66696 6 bus_in_sid[4]
port 70 nsew signal input
rlabel metal3 s 99600 67424 100000 67480 6 bus_in_sid[5]
port 71 nsew signal input
rlabel metal3 s 99600 68208 100000 68264 6 bus_in_sid[6]
port 72 nsew signal input
rlabel metal3 s 99600 68992 100000 69048 6 bus_in_sid[7]
port 73 nsew signal input
rlabel metal3 s 99600 56448 100000 56504 6 bus_in_timers[0]
port 74 nsew signal input
rlabel metal3 s 99600 57232 100000 57288 6 bus_in_timers[1]
port 75 nsew signal input
rlabel metal3 s 99600 58016 100000 58072 6 bus_in_timers[2]
port 76 nsew signal input
rlabel metal3 s 99600 58800 100000 58856 6 bus_in_timers[3]
port 77 nsew signal input
rlabel metal3 s 99600 59584 100000 59640 6 bus_in_timers[4]
port 78 nsew signal input
rlabel metal3 s 99600 60368 100000 60424 6 bus_in_timers[5]
port 79 nsew signal input
rlabel metal3 s 99600 61152 100000 61208 6 bus_in_timers[6]
port 80 nsew signal input
rlabel metal3 s 99600 61936 100000 61992 6 bus_in_timers[7]
port 81 nsew signal input
rlabel metal3 s 99600 47040 100000 47096 6 bus_we_gpios
port 82 nsew signal output
rlabel metal3 s 99600 55664 100000 55720 6 bus_we_serial_ports
port 83 nsew signal output
rlabel metal3 s 99600 62720 100000 62776 6 bus_we_sid
port 84 nsew signal output
rlabel metal3 s 99600 54880 100000 54936 6 bus_we_timers
port 85 nsew signal output
rlabel metal3 s 0 41328 400 41384 6 cs_port[0]
port 86 nsew signal output
rlabel metal3 s 0 42000 400 42056 6 cs_port[1]
port 87 nsew signal output
rlabel metal3 s 0 42672 400 42728 6 cs_port[2]
port 88 nsew signal output
rlabel metal2 s 1344 69600 1400 70000 6 io_in[0]
port 89 nsew signal input
rlabel metal2 s 20384 69600 20440 70000 6 io_in[10]
port 90 nsew signal input
rlabel metal2 s 22288 69600 22344 70000 6 io_in[11]
port 91 nsew signal input
rlabel metal2 s 24192 69600 24248 70000 6 io_in[12]
port 92 nsew signal input
rlabel metal2 s 26096 69600 26152 70000 6 io_in[13]
port 93 nsew signal input
rlabel metal2 s 28000 69600 28056 70000 6 io_in[14]
port 94 nsew signal input
rlabel metal2 s 29904 69600 29960 70000 6 io_in[15]
port 95 nsew signal input
rlabel metal2 s 31808 69600 31864 70000 6 io_in[16]
port 96 nsew signal input
rlabel metal2 s 33712 69600 33768 70000 6 io_in[17]
port 97 nsew signal input
rlabel metal2 s 35616 69600 35672 70000 6 io_in[18]
port 98 nsew signal input
rlabel metal2 s 3248 69600 3304 70000 6 io_in[1]
port 99 nsew signal input
rlabel metal2 s 5152 69600 5208 70000 6 io_in[2]
port 100 nsew signal input
rlabel metal2 s 7056 69600 7112 70000 6 io_in[3]
port 101 nsew signal input
rlabel metal2 s 8960 69600 9016 70000 6 io_in[4]
port 102 nsew signal input
rlabel metal2 s 10864 69600 10920 70000 6 io_in[5]
port 103 nsew signal input
rlabel metal2 s 12768 69600 12824 70000 6 io_in[6]
port 104 nsew signal input
rlabel metal2 s 14672 69600 14728 70000 6 io_in[7]
port 105 nsew signal input
rlabel metal2 s 16576 69600 16632 70000 6 io_in[8]
port 106 nsew signal input
rlabel metal2 s 18480 69600 18536 70000 6 io_in[9]
port 107 nsew signal input
rlabel metal3 s 0 17808 400 17864 6 io_oeb[0]
port 108 nsew signal output
rlabel metal3 s 0 24528 400 24584 6 io_oeb[10]
port 109 nsew signal output
rlabel metal3 s 0 25200 400 25256 6 io_oeb[11]
port 110 nsew signal output
rlabel metal3 s 0 25872 400 25928 6 io_oeb[12]
port 111 nsew signal output
rlabel metal3 s 0 26544 400 26600 6 io_oeb[13]
port 112 nsew signal output
rlabel metal3 s 0 27216 400 27272 6 io_oeb[14]
port 113 nsew signal output
rlabel metal3 s 0 27888 400 27944 6 io_oeb[15]
port 114 nsew signal output
rlabel metal3 s 0 28560 400 28616 6 io_oeb[16]
port 115 nsew signal output
rlabel metal3 s 0 29232 400 29288 6 io_oeb[17]
port 116 nsew signal output
rlabel metal3 s 0 29904 400 29960 6 io_oeb[18]
port 117 nsew signal output
rlabel metal3 s 0 18480 400 18536 6 io_oeb[1]
port 118 nsew signal output
rlabel metal3 s 0 19152 400 19208 6 io_oeb[2]
port 119 nsew signal output
rlabel metal3 s 0 19824 400 19880 6 io_oeb[3]
port 120 nsew signal output
rlabel metal3 s 0 20496 400 20552 6 io_oeb[4]
port 121 nsew signal output
rlabel metal3 s 0 21168 400 21224 6 io_oeb[5]
port 122 nsew signal output
rlabel metal3 s 0 21840 400 21896 6 io_oeb[6]
port 123 nsew signal output
rlabel metal3 s 0 22512 400 22568 6 io_oeb[7]
port 124 nsew signal output
rlabel metal3 s 0 23184 400 23240 6 io_oeb[8]
port 125 nsew signal output
rlabel metal3 s 0 23856 400 23912 6 io_oeb[9]
port 126 nsew signal output
rlabel metal3 s 0 5040 400 5096 6 io_out[0]
port 127 nsew signal output
rlabel metal3 s 0 11760 400 11816 6 io_out[10]
port 128 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 io_out[11]
port 129 nsew signal output
rlabel metal3 s 0 13104 400 13160 6 io_out[12]
port 130 nsew signal output
rlabel metal3 s 0 13776 400 13832 6 io_out[13]
port 131 nsew signal output
rlabel metal3 s 0 14448 400 14504 6 io_out[14]
port 132 nsew signal output
rlabel metal3 s 0 15120 400 15176 6 io_out[15]
port 133 nsew signal output
rlabel metal3 s 0 15792 400 15848 6 io_out[16]
port 134 nsew signal output
rlabel metal3 s 0 16464 400 16520 6 io_out[17]
port 135 nsew signal output
rlabel metal3 s 0 17136 400 17192 6 io_out[18]
port 136 nsew signal output
rlabel metal3 s 0 5712 400 5768 6 io_out[1]
port 137 nsew signal output
rlabel metal3 s 0 6384 400 6440 6 io_out[2]
port 138 nsew signal output
rlabel metal3 s 0 7056 400 7112 6 io_out[3]
port 139 nsew signal output
rlabel metal3 s 0 7728 400 7784 6 io_out[4]
port 140 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 io_out[5]
port 141 nsew signal output
rlabel metal3 s 0 9072 400 9128 6 io_out[6]
port 142 nsew signal output
rlabel metal3 s 0 9744 400 9800 6 io_out[7]
port 143 nsew signal output
rlabel metal3 s 0 10416 400 10472 6 io_out[8]
port 144 nsew signal output
rlabel metal3 s 0 11088 400 11144 6 io_out[9]
port 145 nsew signal output
rlabel metal3 s 99600 44688 100000 44744 6 irq[0]
port 146 nsew signal output
rlabel metal3 s 99600 45472 100000 45528 6 irq[1]
port 147 nsew signal output
rlabel metal3 s 99600 46256 100000 46312 6 irq[2]
port 148 nsew signal output
rlabel metal2 s 37520 69600 37576 70000 6 irqs[0]
port 149 nsew signal input
rlabel metal2 s 39424 69600 39480 70000 6 irqs[1]
port 150 nsew signal input
rlabel metal2 s 41328 69600 41384 70000 6 irqs[2]
port 151 nsew signal input
rlabel metal2 s 43232 69600 43288 70000 6 irqs[3]
port 152 nsew signal input
rlabel metal2 s 45136 69600 45192 70000 6 irqs[4]
port 153 nsew signal input
rlabel metal2 s 47040 69600 47096 70000 6 irqs[5]
port 154 nsew signal input
rlabel metal2 s 48944 69600 49000 70000 6 irqs[6]
port 155 nsew signal input
rlabel metal3 s 99600 784 100000 840 6 la_data_out[0]
port 156 nsew signal output
rlabel metal3 s 99600 8624 100000 8680 6 la_data_out[10]
port 157 nsew signal output
rlabel metal3 s 99600 9408 100000 9464 6 la_data_out[11]
port 158 nsew signal output
rlabel metal3 s 99600 10192 100000 10248 6 la_data_out[12]
port 159 nsew signal output
rlabel metal3 s 99600 10976 100000 11032 6 la_data_out[13]
port 160 nsew signal output
rlabel metal3 s 99600 11760 100000 11816 6 la_data_out[14]
port 161 nsew signal output
rlabel metal3 s 99600 12544 100000 12600 6 la_data_out[15]
port 162 nsew signal output
rlabel metal3 s 99600 13328 100000 13384 6 la_data_out[16]
port 163 nsew signal output
rlabel metal3 s 99600 14112 100000 14168 6 la_data_out[17]
port 164 nsew signal output
rlabel metal3 s 99600 14896 100000 14952 6 la_data_out[18]
port 165 nsew signal output
rlabel metal3 s 99600 15680 100000 15736 6 la_data_out[19]
port 166 nsew signal output
rlabel metal3 s 99600 1568 100000 1624 6 la_data_out[1]
port 167 nsew signal output
rlabel metal3 s 99600 16464 100000 16520 6 la_data_out[20]
port 168 nsew signal output
rlabel metal3 s 99600 17248 100000 17304 6 la_data_out[21]
port 169 nsew signal output
rlabel metal3 s 99600 18032 100000 18088 6 la_data_out[22]
port 170 nsew signal output
rlabel metal3 s 99600 18816 100000 18872 6 la_data_out[23]
port 171 nsew signal output
rlabel metal3 s 99600 19600 100000 19656 6 la_data_out[24]
port 172 nsew signal output
rlabel metal3 s 99600 20384 100000 20440 6 la_data_out[25]
port 173 nsew signal output
rlabel metal3 s 99600 21168 100000 21224 6 la_data_out[26]
port 174 nsew signal output
rlabel metal3 s 99600 21952 100000 22008 6 la_data_out[27]
port 175 nsew signal output
rlabel metal3 s 99600 22736 100000 22792 6 la_data_out[28]
port 176 nsew signal output
rlabel metal3 s 99600 23520 100000 23576 6 la_data_out[29]
port 177 nsew signal output
rlabel metal3 s 99600 2352 100000 2408 6 la_data_out[2]
port 178 nsew signal output
rlabel metal3 s 99600 24304 100000 24360 6 la_data_out[30]
port 179 nsew signal output
rlabel metal3 s 99600 25088 100000 25144 6 la_data_out[31]
port 180 nsew signal output
rlabel metal3 s 99600 25872 100000 25928 6 la_data_out[32]
port 181 nsew signal output
rlabel metal3 s 99600 26656 100000 26712 6 la_data_out[33]
port 182 nsew signal output
rlabel metal3 s 99600 27440 100000 27496 6 la_data_out[34]
port 183 nsew signal output
rlabel metal3 s 99600 28224 100000 28280 6 la_data_out[35]
port 184 nsew signal output
rlabel metal3 s 99600 29008 100000 29064 6 la_data_out[36]
port 185 nsew signal output
rlabel metal3 s 99600 29792 100000 29848 6 la_data_out[37]
port 186 nsew signal output
rlabel metal3 s 99600 30576 100000 30632 6 la_data_out[38]
port 187 nsew signal output
rlabel metal3 s 99600 31360 100000 31416 6 la_data_out[39]
port 188 nsew signal output
rlabel metal3 s 99600 3136 100000 3192 6 la_data_out[3]
port 189 nsew signal output
rlabel metal3 s 99600 32144 100000 32200 6 la_data_out[40]
port 190 nsew signal output
rlabel metal3 s 99600 32928 100000 32984 6 la_data_out[41]
port 191 nsew signal output
rlabel metal3 s 99600 33712 100000 33768 6 la_data_out[42]
port 192 nsew signal output
rlabel metal3 s 99600 34496 100000 34552 6 la_data_out[43]
port 193 nsew signal output
rlabel metal3 s 99600 35280 100000 35336 6 la_data_out[44]
port 194 nsew signal output
rlabel metal3 s 99600 36064 100000 36120 6 la_data_out[45]
port 195 nsew signal output
rlabel metal3 s 99600 36848 100000 36904 6 la_data_out[46]
port 196 nsew signal output
rlabel metal3 s 99600 37632 100000 37688 6 la_data_out[47]
port 197 nsew signal output
rlabel metal3 s 99600 38416 100000 38472 6 la_data_out[48]
port 198 nsew signal output
rlabel metal3 s 99600 39200 100000 39256 6 la_data_out[49]
port 199 nsew signal output
rlabel metal3 s 99600 3920 100000 3976 6 la_data_out[4]
port 200 nsew signal output
rlabel metal3 s 99600 39984 100000 40040 6 la_data_out[50]
port 201 nsew signal output
rlabel metal3 s 99600 40768 100000 40824 6 la_data_out[51]
port 202 nsew signal output
rlabel metal3 s 99600 41552 100000 41608 6 la_data_out[52]
port 203 nsew signal output
rlabel metal3 s 99600 42336 100000 42392 6 la_data_out[53]
port 204 nsew signal output
rlabel metal3 s 99600 43120 100000 43176 6 la_data_out[54]
port 205 nsew signal output
rlabel metal3 s 99600 43904 100000 43960 6 la_data_out[55]
port 206 nsew signal output
rlabel metal3 s 99600 4704 100000 4760 6 la_data_out[5]
port 207 nsew signal output
rlabel metal3 s 99600 5488 100000 5544 6 la_data_out[6]
port 208 nsew signal output
rlabel metal3 s 99600 6272 100000 6328 6 la_data_out[7]
port 209 nsew signal output
rlabel metal3 s 99600 7056 100000 7112 6 la_data_out[8]
port 210 nsew signal output
rlabel metal3 s 99600 7840 100000 7896 6 la_data_out[9]
port 211 nsew signal output
rlabel metal2 s 98448 69600 98504 70000 6 le_hi_act
port 212 nsew signal output
rlabel metal2 s 96544 69600 96600 70000 6 le_lo_act
port 213 nsew signal output
rlabel metal3 s 99600 54096 100000 54152 6 reset_out
port 214 nsew signal output
rlabel metal3 s 0 60144 400 60200 6 rom_bus_in[0]
port 215 nsew signal input
rlabel metal3 s 0 60816 400 60872 6 rom_bus_in[1]
port 216 nsew signal input
rlabel metal3 s 0 61488 400 61544 6 rom_bus_in[2]
port 217 nsew signal input
rlabel metal3 s 0 62160 400 62216 6 rom_bus_in[3]
port 218 nsew signal input
rlabel metal3 s 0 62832 400 62888 6 rom_bus_in[4]
port 219 nsew signal input
rlabel metal3 s 0 63504 400 63560 6 rom_bus_in[5]
port 220 nsew signal input
rlabel metal3 s 0 64176 400 64232 6 rom_bus_in[6]
port 221 nsew signal input
rlabel metal3 s 0 64848 400 64904 6 rom_bus_in[7]
port 222 nsew signal input
rlabel metal3 s 0 54768 400 54824 6 rom_bus_out[0]
port 223 nsew signal output
rlabel metal3 s 0 55440 400 55496 6 rom_bus_out[1]
port 224 nsew signal output
rlabel metal3 s 0 56112 400 56168 6 rom_bus_out[2]
port 225 nsew signal output
rlabel metal3 s 0 56784 400 56840 6 rom_bus_out[3]
port 226 nsew signal output
rlabel metal3 s 0 57456 400 57512 6 rom_bus_out[4]
port 227 nsew signal output
rlabel metal3 s 0 58128 400 58184 6 rom_bus_out[5]
port 228 nsew signal output
rlabel metal3 s 0 58800 400 58856 6 rom_bus_out[6]
port 229 nsew signal output
rlabel metal3 s 0 59472 400 59528 6 rom_bus_out[7]
port 230 nsew signal output
rlabel metal4 s 2224 1538 2384 68238 6 vdd
port 231 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 68238 6 vdd
port 231 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 68238 6 vdd
port 231 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 68238 6 vdd
port 231 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 68238 6 vdd
port 231 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 68238 6 vdd
port 231 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 68238 6 vdd
port 231 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 68238 6 vss
port 232 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 68238 6 vss
port 232 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 68238 6 vss
port 232 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 68238 6 vss
port 232 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 68238 6 vss
port 232 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 68238 6 vss
port 232 nsew ground bidirectional
rlabel metal2 s 4704 0 4760 400 6 wb_clk_i
port 233 nsew signal input
rlabel metal2 s 5600 0 5656 400 6 wb_rst_i
port 234 nsew signal input
rlabel metal2 s 6496 0 6552 400 6 wbs_ack_o
port 235 nsew signal output
rlabel metal2 s 10080 0 10136 400 6 wbs_adr_i[0]
port 236 nsew signal input
rlabel metal2 s 36960 0 37016 400 6 wbs_adr_i[10]
port 237 nsew signal input
rlabel metal2 s 39648 0 39704 400 6 wbs_adr_i[11]
port 238 nsew signal input
rlabel metal2 s 42336 0 42392 400 6 wbs_adr_i[12]
port 239 nsew signal input
rlabel metal2 s 45024 0 45080 400 6 wbs_adr_i[13]
port 240 nsew signal input
rlabel metal2 s 47712 0 47768 400 6 wbs_adr_i[14]
port 241 nsew signal input
rlabel metal2 s 50400 0 50456 400 6 wbs_adr_i[15]
port 242 nsew signal input
rlabel metal2 s 53088 0 53144 400 6 wbs_adr_i[16]
port 243 nsew signal input
rlabel metal2 s 55776 0 55832 400 6 wbs_adr_i[17]
port 244 nsew signal input
rlabel metal2 s 58464 0 58520 400 6 wbs_adr_i[18]
port 245 nsew signal input
rlabel metal2 s 61152 0 61208 400 6 wbs_adr_i[19]
port 246 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 wbs_adr_i[1]
port 247 nsew signal input
rlabel metal2 s 63840 0 63896 400 6 wbs_adr_i[20]
port 248 nsew signal input
rlabel metal2 s 66528 0 66584 400 6 wbs_adr_i[21]
port 249 nsew signal input
rlabel metal2 s 69216 0 69272 400 6 wbs_adr_i[22]
port 250 nsew signal input
rlabel metal2 s 71904 0 71960 400 6 wbs_adr_i[23]
port 251 nsew signal input
rlabel metal2 s 74592 0 74648 400 6 wbs_adr_i[24]
port 252 nsew signal input
rlabel metal2 s 77280 0 77336 400 6 wbs_adr_i[25]
port 253 nsew signal input
rlabel metal2 s 79968 0 80024 400 6 wbs_adr_i[26]
port 254 nsew signal input
rlabel metal2 s 82656 0 82712 400 6 wbs_adr_i[27]
port 255 nsew signal input
rlabel metal2 s 85344 0 85400 400 6 wbs_adr_i[28]
port 256 nsew signal input
rlabel metal2 s 88032 0 88088 400 6 wbs_adr_i[29]
port 257 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 wbs_adr_i[2]
port 258 nsew signal input
rlabel metal2 s 90720 0 90776 400 6 wbs_adr_i[30]
port 259 nsew signal input
rlabel metal2 s 93408 0 93464 400 6 wbs_adr_i[31]
port 260 nsew signal input
rlabel metal2 s 18144 0 18200 400 6 wbs_adr_i[3]
port 261 nsew signal input
rlabel metal2 s 20832 0 20888 400 6 wbs_adr_i[4]
port 262 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 wbs_adr_i[5]
port 263 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 wbs_adr_i[6]
port 264 nsew signal input
rlabel metal2 s 28896 0 28952 400 6 wbs_adr_i[7]
port 265 nsew signal input
rlabel metal2 s 31584 0 31640 400 6 wbs_adr_i[8]
port 266 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 wbs_adr_i[9]
port 267 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 wbs_cyc_i
port 268 nsew signal input
rlabel metal2 s 10976 0 11032 400 6 wbs_dat_i[0]
port 269 nsew signal input
rlabel metal2 s 37856 0 37912 400 6 wbs_dat_i[10]
port 270 nsew signal input
rlabel metal2 s 40544 0 40600 400 6 wbs_dat_i[11]
port 271 nsew signal input
rlabel metal2 s 43232 0 43288 400 6 wbs_dat_i[12]
port 272 nsew signal input
rlabel metal2 s 45920 0 45976 400 6 wbs_dat_i[13]
port 273 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 wbs_dat_i[14]
port 274 nsew signal input
rlabel metal2 s 51296 0 51352 400 6 wbs_dat_i[15]
port 275 nsew signal input
rlabel metal2 s 53984 0 54040 400 6 wbs_dat_i[16]
port 276 nsew signal input
rlabel metal2 s 56672 0 56728 400 6 wbs_dat_i[17]
port 277 nsew signal input
rlabel metal2 s 59360 0 59416 400 6 wbs_dat_i[18]
port 278 nsew signal input
rlabel metal2 s 62048 0 62104 400 6 wbs_dat_i[19]
port 279 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 wbs_dat_i[1]
port 280 nsew signal input
rlabel metal2 s 64736 0 64792 400 6 wbs_dat_i[20]
port 281 nsew signal input
rlabel metal2 s 67424 0 67480 400 6 wbs_dat_i[21]
port 282 nsew signal input
rlabel metal2 s 70112 0 70168 400 6 wbs_dat_i[22]
port 283 nsew signal input
rlabel metal2 s 72800 0 72856 400 6 wbs_dat_i[23]
port 284 nsew signal input
rlabel metal2 s 75488 0 75544 400 6 wbs_dat_i[24]
port 285 nsew signal input
rlabel metal2 s 78176 0 78232 400 6 wbs_dat_i[25]
port 286 nsew signal input
rlabel metal2 s 80864 0 80920 400 6 wbs_dat_i[26]
port 287 nsew signal input
rlabel metal2 s 83552 0 83608 400 6 wbs_dat_i[27]
port 288 nsew signal input
rlabel metal2 s 86240 0 86296 400 6 wbs_dat_i[28]
port 289 nsew signal input
rlabel metal2 s 88928 0 88984 400 6 wbs_dat_i[29]
port 290 nsew signal input
rlabel metal2 s 16352 0 16408 400 6 wbs_dat_i[2]
port 291 nsew signal input
rlabel metal2 s 91616 0 91672 400 6 wbs_dat_i[30]
port 292 nsew signal input
rlabel metal2 s 94304 0 94360 400 6 wbs_dat_i[31]
port 293 nsew signal input
rlabel metal2 s 19040 0 19096 400 6 wbs_dat_i[3]
port 294 nsew signal input
rlabel metal2 s 21728 0 21784 400 6 wbs_dat_i[4]
port 295 nsew signal input
rlabel metal2 s 24416 0 24472 400 6 wbs_dat_i[5]
port 296 nsew signal input
rlabel metal2 s 27104 0 27160 400 6 wbs_dat_i[6]
port 297 nsew signal input
rlabel metal2 s 29792 0 29848 400 6 wbs_dat_i[7]
port 298 nsew signal input
rlabel metal2 s 32480 0 32536 400 6 wbs_dat_i[8]
port 299 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 wbs_dat_i[9]
port 300 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 wbs_dat_o[0]
port 301 nsew signal output
rlabel metal2 s 38752 0 38808 400 6 wbs_dat_o[10]
port 302 nsew signal output
rlabel metal2 s 41440 0 41496 400 6 wbs_dat_o[11]
port 303 nsew signal output
rlabel metal2 s 44128 0 44184 400 6 wbs_dat_o[12]
port 304 nsew signal output
rlabel metal2 s 46816 0 46872 400 6 wbs_dat_o[13]
port 305 nsew signal output
rlabel metal2 s 49504 0 49560 400 6 wbs_dat_o[14]
port 306 nsew signal output
rlabel metal2 s 52192 0 52248 400 6 wbs_dat_o[15]
port 307 nsew signal output
rlabel metal2 s 54880 0 54936 400 6 wbs_dat_o[16]
port 308 nsew signal output
rlabel metal2 s 57568 0 57624 400 6 wbs_dat_o[17]
port 309 nsew signal output
rlabel metal2 s 60256 0 60312 400 6 wbs_dat_o[18]
port 310 nsew signal output
rlabel metal2 s 62944 0 63000 400 6 wbs_dat_o[19]
port 311 nsew signal output
rlabel metal2 s 14560 0 14616 400 6 wbs_dat_o[1]
port 312 nsew signal output
rlabel metal2 s 65632 0 65688 400 6 wbs_dat_o[20]
port 313 nsew signal output
rlabel metal2 s 68320 0 68376 400 6 wbs_dat_o[21]
port 314 nsew signal output
rlabel metal2 s 71008 0 71064 400 6 wbs_dat_o[22]
port 315 nsew signal output
rlabel metal2 s 73696 0 73752 400 6 wbs_dat_o[23]
port 316 nsew signal output
rlabel metal2 s 76384 0 76440 400 6 wbs_dat_o[24]
port 317 nsew signal output
rlabel metal2 s 79072 0 79128 400 6 wbs_dat_o[25]
port 318 nsew signal output
rlabel metal2 s 81760 0 81816 400 6 wbs_dat_o[26]
port 319 nsew signal output
rlabel metal2 s 84448 0 84504 400 6 wbs_dat_o[27]
port 320 nsew signal output
rlabel metal2 s 87136 0 87192 400 6 wbs_dat_o[28]
port 321 nsew signal output
rlabel metal2 s 89824 0 89880 400 6 wbs_dat_o[29]
port 322 nsew signal output
rlabel metal2 s 17248 0 17304 400 6 wbs_dat_o[2]
port 323 nsew signal output
rlabel metal2 s 92512 0 92568 400 6 wbs_dat_o[30]
port 324 nsew signal output
rlabel metal2 s 95200 0 95256 400 6 wbs_dat_o[31]
port 325 nsew signal output
rlabel metal2 s 19936 0 19992 400 6 wbs_dat_o[3]
port 326 nsew signal output
rlabel metal2 s 22624 0 22680 400 6 wbs_dat_o[4]
port 327 nsew signal output
rlabel metal2 s 25312 0 25368 400 6 wbs_dat_o[5]
port 328 nsew signal output
rlabel metal2 s 28000 0 28056 400 6 wbs_dat_o[6]
port 329 nsew signal output
rlabel metal2 s 30688 0 30744 400 6 wbs_dat_o[7]
port 330 nsew signal output
rlabel metal2 s 33376 0 33432 400 6 wbs_dat_o[8]
port 331 nsew signal output
rlabel metal2 s 36064 0 36120 400 6 wbs_dat_o[9]
port 332 nsew signal output
rlabel metal2 s 8288 0 8344 400 6 wbs_stb_i
port 333 nsew signal input
rlabel metal2 s 9184 0 9240 400 6 wbs_we_i
port 334 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 14466372
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/AS2650/openlane/wrapped_as2650/runs/23_11_21_01_04/results/signoff/wrapped_as2650.magic.gds
string GDS_START 568484
<< end >>

