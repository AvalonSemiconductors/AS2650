* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

.subckt wrapped_as2650 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vdd vss wb_clk_i
XFILLER_39_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7957__A2 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7963_ _4444_ _3126_ _3134_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5968__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _0405_ _2128_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6425__I _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7894_ _2971_ _2951_ _2284_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7709__A2 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8906__A1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7965__B _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ _1910_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8382__A2 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6776_ _1976_ _0744_ _1974_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8921__A4 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_3_3__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6932__A3 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8515_ _1033_ _2155_ _3659_ _3668_ _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5727_ _1046_ _1048_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4943__A2 _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8134__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8446_ _2903_ _3581_ _3396_ _3273_ _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ _0984_ _0965_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4609_ as2650.cycle\[7\] as2650.cycle\[6\] as2650.cycle\[5\] as2650.cycle\[4\] _4190_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__6696__A2 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7893__A1 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8377_ _2217_ _2934_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _4197_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7328_ _2528_ _2495_ _2345_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6448__A2 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7259_ _2460_ _2407_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5120__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5959__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6335__I _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4631__A1 as2650.alu_op\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4934__A2 _4514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7166__I _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7884__A1 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6439__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8725__I _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_wb_clk_i clknet_opt_4_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8061__A1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8600__A3 _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4960_ _4524_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4622__A1 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _4471_ _4472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8364__A2 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _1028_ _1871_ _1878_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6561_ _1817_ _1820_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8116__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8300_ _0901_ _4363_ _3461_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5512_ as2650.stack\[7\]\[14\] _0392_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9280_ _0229_ clknet_leaf_43_wb_clk_i as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6492_ _1750_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8231_ _3360_ _3394_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7875__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5443_ _0592_ as2650.stack\[1\]\[13\] as2650.stack\[0\]\[13\] _0586_ _0778_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7804__I _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8162_ _0385_ _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5374_ _0698_ _0700_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7113_ _1572_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8093_ _1544_ _2482_ _3259_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7044_ _2238_ _2247_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7679__C _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8052__A1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8995_ _0495_ _4054_ _4059_ _3970_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7946_ _2199_ _3105_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7877_ _3051_ _3052_ _3054_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8355__A2 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6828_ _2035_ _2042_ _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8303__C _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6759_ _1957_ _1988_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9118__D _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6118__A1 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7866__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8429_ _2177_ _2334_ _3349_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7618__A1 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8291__A1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7094__A2 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6841__A2 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4852__A1 as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8594__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6065__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8346__A2 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9328__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5332__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7609__A1 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8282__A1 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7085__A2 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8282__B2 _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5090_ _0420_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5096__A1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7499__C _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6045__B1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7800_ _2986_ _2987_ _2988_ _2982_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_64_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8780_ _4118_ _1168_ _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5992_ _0541_ _1192_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7731_ _4427_ _4425_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6060__A3 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4943_ as2650.holding_reg\[1\] _4319_ _4523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8337__A2 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7662_ _2854_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4874_ _4451_ _4455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6613_ _1115_ _1862_ _1867_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6899__A2 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7593_ _0985_ _1595_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6544_ _1737_ _1806_ _1807_ _1783_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_9332_ _0281_ clknet_leaf_62_wb_clk_i net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5571__A2 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9263_ _0212_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6475_ _1727_ _1741_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8214_ _3343_ _3346_ _3378_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5426_ _0759_ _0760_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9194_ _0143_ clknet_opt_3_0_wb_clk_i net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8145_ _3308_ _3309_ _3310_ _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5357_ _0691_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5054__I _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8273__A1 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7076__A2 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8076_ as2650.stack\[6\]\[1\] _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ _0524_ _0527_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4893__I _4473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7027_ _0404_ _4123_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8025__A1 _4471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8576__A2 _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8978_ _1551_ _4017_ _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7929_ _2220_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8328__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6339__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7000__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5562__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7839__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8500__A2 _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6511__A1 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5865__A3 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8264__A1 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7067__A2 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5078__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4825__A1 _4404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8016__A1 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9150__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8319__A2 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5250__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__B2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5002__A1 _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6750__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _4150_ _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6750__B2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _1544_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5305__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5211_ _4300_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6191_ _1450_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8255__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5142_ _4455_ _4452_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7058__A2 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5069__A1 _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ as2650.holding_reg\[2\] _4320_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8007__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8901_ as2650.stack\[2\]\[1\] _3976_ _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6281__A3 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8558__A2 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8832_ _2021_ _3919_ _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7957__C _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6569__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7230__A2 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5975_ _1249_ _1181_ _1266_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8763_ as2650.stack\[7\]\[8\] _3871_ _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7714_ _2476_ _2899_ _2905_ _2695_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4926_ _4506_ _4507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8694_ _1027_ _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7645_ _2838_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4857_ _4437_ _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8730__A2 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7576_ _1631_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4788_ _4365_ _4368_ _4369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5544__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4888__I _4468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6527_ _1791_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9315_ _0264_ clknet_leaf_47_wb_clk_i as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7264__I _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6458_ _1724_ _1725_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9246_ _0195_ clknet_leaf_54_wb_clk_i as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5409_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9177_ _0126_ clknet_leaf_15_wb_clk_i as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6389_ _1659_ _1664_ _1473_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8128_ as2650.stack\[3\]\[2\] _3243_ _3241_ _3294_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7049__A2 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8059_ _2803_ _2130_ _2141_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6272__A3 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5480__B2 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7221__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6024__A3 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8044__B _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5232__A1 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6980__A1 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7883__B _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5535__A2 _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7288__A2 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7902__I _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8237__A1 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7460__A2 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5471__A1 _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7212__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5223__A1 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8960__A2 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7763__A3 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6253__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5760_ as2650.pc\[3\] _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6971__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4711_ _4291_ _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _1018_ _1009_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7430_ _4242_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8712__A2 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4642_ _4220_ _4222_ _4180_ _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6723__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7361_ _2558_ _2560_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4573_ _4153_ _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9216__D _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6312_ _1595_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9100_ _0049_ clknet_leaf_65_wb_clk_i as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8476__A1 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7292_ _2383_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9031_ _4088_ _4090_ _1428_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6243_ _4148_ _1522_ _1524_ _1527_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_89_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8908__I _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7812__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8228__A1 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6174_ _4123_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8779__A2 _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5125_ _0459_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7987__B1 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ as2650.stack\[2\]\[9\] _4473_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5462__A1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7203__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8815_ _0845_ _3893_ _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8746_ _1896_ _3856_ _3860_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5958_ _0506_ _1224_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4909_ _4489_ _4490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8677_ _3814_ _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5889_ _0332_ _0696_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7628_ _4248_ _2731_ _2730_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8311__C _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7559_ _2664_ _2752_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5507__I _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8467__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9229_ _0178_ clknet_leaf_30_wb_clk_i as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8219__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8039__B _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8981__C _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__A3 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7878__B _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8553__I _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7__f_wb_clk_i clknet_0_wb_clk_i clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7169__I _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8942__A2 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6953__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9069__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5508__A2 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_14_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_14_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5417__I _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8458__A1 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7681__A2 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8891__C _3970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7433__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8630__A1 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5444__A1 as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4991__I _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6930_ _2128_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7197__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6861_ _0860_ _2085_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8933__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8600_ _3678_ _3739_ _3749_ _3750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5812_ _1087_ _1120_ _1125_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6792_ _1993_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5743_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8531_ _1564_ _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8462_ as2650.pc\[13\] as2650.pc\[12\] _2854_ _3553_ _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5674_ _0657_ as2650.r123_2\[0\]\[3\] _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8131__C _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7413_ _2600_ _2185_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4625_ _4186_ _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8393_ _3551_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5327__I _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6172__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8449__A1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7344_ _2543_ _1271_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8449__B2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4556_ _4136_ _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_5_0_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_opt_5_0_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7275_ _2476_ _2469_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7121__A1 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9014_ _1404_ _2300_ _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6226_ _1458_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7672__A2 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6158__I _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ _4193_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\] _0339_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8621__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6088_ _1367_ _1371_ _1364_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8373__I _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5435__B2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _4469_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7188__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9211__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8924__A2 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8729_ _3821_ _3845_ _3850_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6163__A2 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5910__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput20 net20 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7112__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput31 net31 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5674__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8612__A1 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9379__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8216__C _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7627__I _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7351__A1 _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6154__A2 _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7351__B2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5390_ _0626_ _0723_ _0721_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7362__I _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__C _4499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7060_ _0929_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7654__A2 _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8851__A1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ _1285_ _1286_ _1300_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8603__A1 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9234__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7962_ _3132_ _3133_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6913_ _4190_ _0949_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout49_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7893_ _3069_ _2264_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8906__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6917__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6844_ _2068_ _2070_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7590__A1 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6775_ _2002_ _2003_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8514_ _1438_ _3662_ _3666_ _3667_ _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5726_ _1050_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8445_ _3600_ _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5657_ _0986_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4608_ as2650.cycle\[2\] _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8376_ _3089_ _3263_ _3534_ _3034_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5588_ _0917_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7893__A2 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4896__I as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7327_ _2340_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8368__I _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4539_ as2650.cycle\[2\] _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7272__I _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8842__A1 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7258_ as2650.pc\[1\] _0349_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ _0870_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7189_ _2389_ _2391_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7581__A1 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6384__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7884__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4698__A2 _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7182__I _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9257__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8061__A2 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A2 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9010__A1 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4890_ _4469_ _4470_ _4471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7357__I _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6375__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6261__I _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _1331_ _1696_ _1823_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5511_ _4348_ _0814_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6491_ _1735_ _1751_ _1756_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7324__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8230_ _2595_ _2184_ _3393_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5442_ _0491_ _0775_ _0776_ _0502_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7875__A2 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8161_ _3195_ _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5373_ _4467_ _0708_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7112_ _2313_ _2315_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8092_ _1074_ _1616_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8824__A1 _4463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7043_ _1385_ _2238_ _2247_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8137__B _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8052__A2 _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5340__I _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8994_ _0495_ _4055_ _4058_ _4054_ _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7945_ as2650.cycle\[4\] _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5810__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4613__A2 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9001__A1 _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7876_ _3043_ _4267_ _2200_ _3053_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6827_ _2039_ _2040_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7563__A1 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6366__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6171__I _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6758_ _1959_ _1987_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5709_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6118__A2 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6689_ _1919_ _1848_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8428_ _1616_ _2910_ _3584_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7866__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8359_ _2315_ _3511_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8815__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__A1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7177__I _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A2 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__I _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7306__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8806__A1 _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8282__A2 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4843__A2 _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _1271_ _1193_ _1281_ _1192_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7730_ _1387_ _2273_ _1473_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4942_ _4377_ _4381_ _4522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_45_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7661_ as2650.pc\[11\] _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4873_ _4451_ _4453_ _4454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ as2650.stack\[5\]\[7\] _1863_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7592_ _2777_ _2316_ _2783_ _2786_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5020__A2 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9331_ _0280_ clknet_3_1__leaf_wb_clk_i as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6543_ _0442_ _1717_ _1780_ as2650.r0\[1\] _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9008__S _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9262_ _0211_ clknet_leaf_37_wb_clk_i as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6474_ _1728_ _1740_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8213_ _3368_ _3377_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5425_ _4136_ _4263_ _0356_ _0640_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_9193_ _0142_ clknet_leaf_25_wb_clk_i net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8144_ _1465_ _2298_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5356_ _4164_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8075_ _0380_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5287_ _0622_ _0521_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5087__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6284__A1 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7481__B1 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7026_ _2230_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__A2 _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8025__A2 _4483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5070__I _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8977_ _1680_ _2195_ _4040_ _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7784__A1 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4598__A1 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7928_ _3096_ _3099_ _3103_ _3031_ _0927_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_93_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7859_ _1154_ _2298_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7839__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8264__A2 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_39_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__A2 _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8016__A2 _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8505__B _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6025__B _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5002__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4761__A1 _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5583__C _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\] _4301_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6190_ _1368_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ _4456_ _0472_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8255__A2 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7058__A3 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7303__C _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _4442_ _4272_ _4264_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_96_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8900_ _3975_ _1062_ _3977_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8007__A2 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6018__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8831_ _0488_ _3915_ _3917_ as2650.r123\[2\]\[2\] _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8762_ _3869_ _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5974_ _1186_ _1251_ _1265_ _1218_ _1220_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8134__C _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7713_ net51 _0936_ _2904_ _2187_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4925_ _4504_ _4505_ _4506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8693_ _3825_ _3816_ _3826_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7644_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4856_ _4398_ _4436_ _4437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7575_ _2763_ _2770_ _2586_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4787_ as2650.r123\[1\]\[7\] as2650.r123\[0\]\[7\] as2650.r123_2\[1\]\[7\] as2650.r123_2\[0\]\[7\]
+ _4367_ _4112_ _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9314_ _0263_ clknet_leaf_47_wb_clk_i as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6526_ _1766_ _1768_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9245_ _0194_ clknet_leaf_54_wb_clk_i as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5065__I as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6457_ _1265_ _1705_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5408_ as2650.r0\[6\] _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9176_ _0125_ clknet_leaf_15_wb_clk_i as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6388_ _1663_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8127_ _3292_ _4472_ _3204_ _3293_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5339_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7049__A3 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6257__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8058_ _2380_ _2604_ _3225_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__A2 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7009_ _2136_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6272__A4 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6009__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6009__B2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6__f_wb_clk_i clknet_0_wb_clk_i clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7757__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7509__A1 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7883__C _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4743__A1 _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6496__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8237__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6248__A1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7996__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5578__C _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _4155_ _4196_ _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7793__C _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5690_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _4221_ _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6723__A2 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7360_ _2512_ _2516_ _2559_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4572_ as2650.alu_op\[0\] _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6311_ net2 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7291_ _2491_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6487__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9030_ _3006_ _4089_ _4082_ _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6242_ _1429_ _1525_ _0431_ _1526_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6173_ _4225_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5613__I _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6239__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8779__A3 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5124_ _4212_ _0460_ _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7987__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7987__B2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5055_ _0384_ as2650.stack\[1\]\[9\] as2650.stack\[0\]\[9\] _0393_ _0394_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5462__A2 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8145__B _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7739__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8814_ as2650.r123\[1\]\[6\] _3901_ _3898_ _1822_ _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5214__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6411__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8745_ as2650.stack\[7\]\[2\] _3857_ _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ as2650.r123_2\[0\]\[2\] _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4908_ _4488_ _4489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8676_ _3813_ _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8164__A1 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5888_ _4170_ _1157_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7627_ _2820_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4839_ _4182_ _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7911__A1 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _2666_ _2752_ _2753_ _2699_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _1772_ _1773_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8467__A2 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7489_ _2647_ _2493_ _2686_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6478__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9228_ _0177_ clknet_leaf_29_wb_clk_i as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5150__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9159_ _0108_ clknet_leaf_45_wb_clk_i as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7978__A1 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9290__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7978__B2 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7878__C _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8055__B _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6354__I _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__A1 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7894__B _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8942__A3 _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4964__A1 _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8155__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8502__C _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7185__I _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6705__A2 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8458__A2 _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7913__I _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_54_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6469__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7969__A1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8630__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5444__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6264__I _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6860_ _0782_ _2082_ _2061_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8394__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5811_ as2650.stack\[0\]\[3\] _1121_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8933__A3 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _1995_ _2019_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8530_ _3682_ _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5742_ as2650.pc\[1\] _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8146__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8461_ _3123_ _3616_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5673_ _0958_ _1001_ _1002_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9227__D _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7412_ _2607_ _2610_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9163__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _4180_ _4204_ _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8392_ _1693_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6172__A3 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7343_ _0554_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ as2650.ins_reg\[4\] _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7274_ _2475_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7121__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9013_ _3638_ _4075_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6225_ _1166_ _0884_ _1491_ _1507_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_106_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _4232_ _4167_ _4340_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_97_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8082__B1 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8654__I _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5107_ _0444_ _4176_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8621__A2 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6087_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5435__A2 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6632__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _0376_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6174__I _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8385__A1 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7188__A2 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8385__B2 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ _2190_ _2195_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4946__A1 _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8728_ as2650.stack\[3\]\[10\] _3848_ _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8137__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8659_ as2650.stack\[6\]\[2\] _3800_ _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6699__A1 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5371__A1 as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7648__B1 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput21 net21 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput32 net32 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7112__A2 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput43 net43 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6349__I _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5123__A1 _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5674__A2 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4721__I1 as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6218__A4 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8612__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8376__A1 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__A1 _4503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8679__A2 _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7351__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6154__A3 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__A1 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8739__I _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8300__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6259__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8851__A2 _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6010_ _1219_ _1297_ _1299_ _1180_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8603__A2 _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7961_ _2562_ _3131_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6912_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7892_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6843_ _2046_ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6917__A2 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7818__I _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8119__A1 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _1978_ _1982_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7590__A2 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8513_ _0924_ _1449_ _2235_ _1444_ _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5338__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8444_ as2650.pc\[13\] _3599_ _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5656_ _0964_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4607_ as2650.cycle\[3\] _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8375_ _2815_ _3533_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4787__S0 _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5587_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7326_ _2474_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4538_ as2650.cycle\[0\] _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6169__I _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7257_ as2650.pc\[2\] net8 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6302__B1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8842__A2 _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6208_ _0873_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7188_ _0352_ _0320_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_58_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9059__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6139_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__I _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8317__C _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8358__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7728__I _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4919__A1 _4495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4919__B2 _4474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5248__I _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5647__A2 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A2 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8349__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9010__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7021__A1 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5510_ _0542_ _0821_ _0843_ _0321_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_125_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6490_ _1753_ _1754_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7324__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8521__A1 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5441_ as2650.stack\[6\]\[13\] _0588_ _4484_ as2650.stack\[7\]\[13\] _0776_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5335__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7373__I _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8160_ _3127_ _3312_ _3315_ _2313_ _3190_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5372_ _0702_ _0703_ _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7111_ _2314_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7088__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8091_ _1074_ _3256_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5099__B1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6835__A1 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7042_ _2240_ _2246_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9240__D _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8588__A1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8993_ _4056_ _4057_ _3503_ _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7944_ _3104_ _4188_ _3112_ _3117_ _3118_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5110__I1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7875_ _2531_ _2339_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9001__A2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7548__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7012__A1 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _2009_ _2034_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6757_ _1961_ _1986_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5574__A1 _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ _1031_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6688_ _1827_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6118__A3 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8512__A1 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8427_ _2886_ _1543_ _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5639_ _0946_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7866__A3 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5877__A2 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8358_ _3263_ _3517_ _3064_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7309_ _2350_ _2504_ _2509_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8289_ _2184_ _2703_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8815__A2 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8328__B _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8047__C _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7251__A1 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7003__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8200__B1 _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__A2 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8751__A1 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5565__A1 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6762__B1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7306__A2 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8503__A1 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__A1 _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9224__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__A2 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7126__C _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7921__I _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7490__A1 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7242__A1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _1193_ _1278_ _1280_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8990__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4941_ as2650.r123\[0\]\[1\] _4521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7660_ _2646_ _2851_ _2853_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4872_ _4452_ _4453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8742__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6611_ _1108_ _1862_ _1866_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5556__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7591_ _2332_ _2784_ _2785_ _2695_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9330_ _0279_ clknet_leaf_62_wb_clk_i as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6542_ as2650.r0\[3\] _1014_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4721__S _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9261_ _0210_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6473_ _1729_ _1730_ _1739_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5616__I _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8212_ _3369_ _3376_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5424_ _0670_ _0669_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9192_ _0141_ clknet_leaf_25_wb_clk_i net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8143_ _1075_ _3264_ _2492_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5355_ _4367_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8074_ _1590_ as2650.stack\[3\]\[1\] as2650.stack\[2\]\[1\] _0377_ _3241_ _3242_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5286_ _0514_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7481__A1 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7025_ _1424_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7481__B2 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5__f_wb_clk_i clknet_0_wb_clk_i clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8976_ _3638_ _4042_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7784__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8981__A1 _4466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7927_ _3086_ _3102_ _0963_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7858_ _3035_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8733__A1 _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6809_ _0611_ _2036_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5547__A1 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9247__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7789_ _1488_ _2969_ _2978_ _1573_ _2225_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5526__I _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7472__A1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5261__I _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6027__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8972__A1 _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8505__C _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4605__I _4126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8724__A1 _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7916__I _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8521__B _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4761__A2 _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5436__I _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _0314_ _0469_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7058__A4 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7463__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6267__I _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8830_ _3921_ _3922_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8963__A1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8761_ _3869_ _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5973_ _0437_ _1228_ _1264_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7712_ _2903_ _2338_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4924_ _4132_ _4177_ _4505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8692_ as2650.stack\[5\]\[12\] _3819_ _3826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7643_ _1475_ _1663_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4855_ _4433_ _4435_ _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8191__A2 _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7574_ _2322_ _2767_ _2769_ _2421_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4786_ _4366_ _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8150__C _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9313_ _0262_ clknet_leaf_47_wb_clk_i as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6525_ _1774_ _1789_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_109_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9244_ _0193_ clknet_leaf_14_wb_clk_i as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ as2650.r123_2\[1\]\[2\] _1699_ _1722_ _1723_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _0638_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9175_ _0124_ clknet_leaf_45_wb_clk_i as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6387_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8126_ _3245_ as2650.stack\[1\]\[2\] as2650.stack\[0\]\[2\] _3205_ _3293_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5338_ net10 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8057_ _2184_ _2425_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5269_ as2650.holding_reg\[4\] _0422_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7008_ _1513_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6009__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7206__A1 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8392__I _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6905__I _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7757__A2 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8954__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8959_ _2999_ _1363_ _1399_ _1405_ _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_43_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6193__A1 _4465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8995__C _3970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7693__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6496__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8567__I _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6248__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6087__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7996__A2 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4763__C _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4640_ _4125_ _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6184__A1 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4571_ _4133_ _4145_ _4151_ _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6310_ _0691_ _4182_ _4332_ _1381_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7290_ as2650.pc\[3\] _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6241_ _0692_ _0833_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _1454_ _1456_ _1382_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7436__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6239__A2 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ _4384_ _0358_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8779__A4 _4446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5054_ _0386_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9092__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8936__A1 _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7739__A2 _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8813_ _3908_ _3909_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5956_ _1222_ _1181_ _1248_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8744_ _1894_ _3856_ _3859_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4907_ _4487_ _4488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8675_ _0917_ _3812_ _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5887_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7626_ as2650.addr_buff\[0\] as2650.addr_buff\[1\] as2650.addr_buff\[2\] _2820_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4838_ _4352_ _4418_ _4419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7911__A2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7557_ _1110_ _0830_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5922__A1 _4459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5076__I _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _4349_ _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6508_ _0438_ _1006_ _1023_ _4353_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7488_ _2676_ _2685_ _2374_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6478__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9227_ _0176_ clknet_3_6__leaf_wb_clk_i as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6439_ _0331_ _0962_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7291__I _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5804__I _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9158_ _0107_ clknet_leaf_45_wb_clk_i as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5150__A2 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8109_ _0349_ _4380_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9089_ _0038_ clknet_leaf_60_wb_clk_i as2650.r123_2\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5989__A1 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A1 _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8927__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6402__A2 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4964__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8155__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6166__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5913__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7666__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6469__A2 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7418__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_23_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_23_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7969__A2 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8918__A1 _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8394__A2 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _1079_ _1120_ _1124_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8760__I _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6790_ _1998_ _2018_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_62_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ _0331_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8146__A2 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8460_ _1025_ _3528_ _3615_ _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5672_ as2650.stack\[2\]\[10\] _0991_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7411_ _2540_ _0675_ _2609_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4623_ _4183_ _4187_ _4203_ _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8391_ _3095_ _3532_ _3547_ _3549_ _3299_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7342_ _2350_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4554_ _4134_ _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7657__A1 _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7657__B2 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7273_ _0951_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9243__D _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9012_ as2650.overflow _4070_ _4074_ _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6224_ _1503_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7409__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6155_ _1438_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5106_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8082__B2 _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _0931_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ _4468_ as2650.psu\[1\] _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8909__A1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8385__A2 _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6988_ _2194_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8603__C _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8727_ _3818_ _3845_ _3849_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4946__A2 _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5939_ _4445_ _4448_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_139_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8137__A2 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6190__I _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4703__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6148__A1 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7345__B1 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8658_ _1894_ _3799_ _3802_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6123__C _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7609_ _2735_ _2733_ _2803_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7896__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8589_ _0673_ _2797_ _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5371__A2 _4485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7648__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7648__B2 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput11 net11 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput22 net22 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput33 net33 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput44 net44 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6871__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7820__A1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6623__A2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4634__A1 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8376__A2 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__A2 _4510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8128__A2 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7336__B1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7924__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7145__B _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8300__A2 _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4873__A1 _4451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8064__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6275__I _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6614__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7960_ _2562_ _3131_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_82_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6911_ _4425_ _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7891_ _3035_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ _1993_ _2020_ _2047_ _2024_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__6378__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6917__A3 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6773_ _1975_ _1977_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9238__D _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5724_ _0585_ _0954_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8512_ _1472_ _2261_ _3665_ _1462_ _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7878__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5655_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8443_ _2886_ _2854_ _3553_ _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_opt_4_0_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9280__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _4185_ _4186_ _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8374_ _0985_ _3516_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5586_ _4486_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5353__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__S1 _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7325_ _0936_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4537_ _4113_ _4117_ _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7256_ _2350_ _2457_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__A1 _4477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__B2 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6207_ as2650.psl\[1\] _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7187_ _4386_ _4458_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4864__A1 _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8055__A1 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6138_ _4116_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__A1 _4451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ as2650.psl\[6\] _4367_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8614__B _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__B1 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5529__I _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5592__A2 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__B _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7744__I _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5344__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8818__B1 _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7097__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8046__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9153__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8349__A2 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7021__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5032__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5583__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8521__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5440_ _0585_ as2650.stack\[5\]\[13\] as2650.stack\[4\]\[13\] _0393_ _0775_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5371_ as2650.stack\[7\]\[12\] _4485_ _4490_ _0706_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5174__I as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7110_ _0938_ _1455_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8285__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7088__A2 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8090_ _1074_ _3256_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_113_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5099__B2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7041_ _2202_ _2241_ _2245_ _1574_ _1459_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__8485__I _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6835__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5902__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8037__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8037__B2 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6219__B _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8588__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_4__f_wb_clk_i clknet_0_wb_clk_i clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6599__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8992_ _4503_ _3009_ _4467_ _0972_ _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_94_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout54_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7943_ _1427_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5110__I2 as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7874_ _2324_ _2941_ _2368_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7012__A2 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _2033_ _2043_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6220__B1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6756_ _1964_ _1985_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5574__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5707_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6687_ _1824_ _1916_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8512__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8426_ _2144_ _3582_ _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5638_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8357_ _0986_ _3516_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5569_ _0901_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7308_ _2358_ _2507_ _2508_ _2135_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8276__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8288_ _3449_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6908__I _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6826__A2 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7239_ _2440_ _0319_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9176__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4837__A1 _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8028__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8028__B2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5968__B _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8200__A1 _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7003__A2 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8200__B2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6762__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8503__A2 _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6514__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__A2 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5722__I _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4828__A1 _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8238__C _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8019__A1 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6039__B _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7242__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ _4107_ _4287_ _4520_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8990__A2 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ as2650.idx_ctrl\[0\] _4452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5169__I _4508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6610_ as2650.stack\[5\]\[6\] _1863_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7590_ _2780_ _2526_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5556__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6541_ _1700_ _1803_ _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4801__I _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6505__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6472_ _1733_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9260_ _0209_ clknet_leaf_37_wb_clk_i as2650.stack\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5423_ _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8211_ _3371_ _3372_ _3374_ _3375_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_9191_ _0140_ clknet_leaf_25_wb_clk_i net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8258__A1 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8142_ _2491_ _1073_ _3264_ _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5354_ _4348_ _0634_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7333__B _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8073_ _4487_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5285_ _0616_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4819__A1 _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7024_ _4141_ _2228_ _2229_ _1644_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7481__A2 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8430__A1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8975_ _4025_ _1048_ _4041_ _4042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7784__A3 _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8981__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7926_ _3101_ _2382_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5795__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7857_ _2141_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _1979_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6744__A1 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7788_ _2348_ _2975_ _2977_ _2223_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _1941_ _1945_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__I _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8497__A1 _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8497__B2 _4169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8409_ _3091_ _3565_ _3566_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8249__A1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7243__B _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5483__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8853__I _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__A2 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5235__A1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8972__A2 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8724__A2 _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5717__I _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8488__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5710__A2 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7463__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5070_ _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8660__A1 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8412__A1 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8963__A2 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8760_ _3868_ _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5972_ _1253_ _1261_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7711_ as2650.addr_buff\[4\] _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4923_ _4135_ _4217_ _4294_ _4504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8691_ _1020_ _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7642_ _2153_ _2835_ _2386_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4854_ _4434_ as2650.addr_buff\[5\] _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8431__C _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7328__B _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7573_ _2744_ _2768_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4785_ _4173_ _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9312_ _0261_ clknet_leaf_17_wb_clk_i net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4531__I _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8479__A1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ _1777_ _1788_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9243_ _0192_ clknet_leaf_0_wb_clk_i as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8938__I _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7151__A1 _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6455_ _1702_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5406_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9174_ _0123_ clknet_leaf_44_wb_clk_i as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6386_ _0922_ _1661_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8125_ as2650.stack\[2\]\[2\] _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5337_ _0667_ _0668_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_115_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8056_ _2420_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8651__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5268_ _0432_ _0427_ _0523_ _0533_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7007_ _2205_ _2213_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8673__I _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _0295_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8403__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8403__B2 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9214__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8958_ _3078_ _4023_ _4024_ _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7909_ _2137_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8889_ net20 _3962_ _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8622__B _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6921__I _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7390__A1 _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6368__I _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8642__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7199__I _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8945__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6708__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5447__I _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6184__A2 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ _4148_ _4150_ _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6240_ _0832_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5695__A1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6171_ _1455_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5182__I _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5122_ _4378_ _4382_ _4397_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7436__A2 _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8633__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9237__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8493__I _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5053_ _4483_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8936__A2 _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8812_ _0774_ _3893_ _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8743_ as2650.stack\[7\]\[1\] _3857_ _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5955_ _1186_ _1226_ _1247_ _1219_ _1220_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _4486_ _4483_ _4487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8674_ _4495_ _1050_ _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5886_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7625_ _2388_ _2798_ _2802_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4837_ _4354_ _4355_ _4417_ _4418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7372__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7911__A3 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7556_ _2700_ _2698_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4768_ _4280_ _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6507_ _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7124__A1 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7487_ _2647_ _2575_ _2684_ _2586_ _2588_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7572__I _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4699_ _4207_ _4269_ _4279_ _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_9226_ _0175_ clknet_leaf_32_wb_clk_i as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8872__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6438_ _0329_ _0984_ _1701_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6883__B1 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9157_ _0106_ clknet_leaf_45_wb_clk_i as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6369_ as2650.stack\[6\]\[9\] _1650_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8108_ _0453_ _0340_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9088_ _0037_ clknet_leaf_59_wb_clk_i as2650.r123_2\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8039_ as2650.stack\[7\]\[0\] _3202_ _0501_ _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6137__B _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4661__A2 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6938__A1 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7363__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6166__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5913__A2 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8863__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6098__I _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8615__A1 _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5429__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7969__A3 _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5730__I as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_63_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8918__A2 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9040__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6929__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4790__B _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _1053_ _1062_ _1064_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5671_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7410_ _2608_ _2581_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4622_ _4195_ _4202_ _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8390_ _0505_ _3369_ _3287_ _3548_ _3251_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_129_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5904__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7341_ _2540_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4553_ as2650.alu_op\[0\] _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5905__I _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7657__A2 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6314__C1 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8854__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7272_ _2473_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5212__S0 _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9011_ _2215_ _4071_ _4073_ _4070_ _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6223_ _4330_ _0291_ _0421_ _0532_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7409__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8606__A1 _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _4311_ _4410_ _1374_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__B _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5105_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8082__A2 _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6085_ _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_85_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6093__A1 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _4509_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7593__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6987_ _0969_ _2193_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8790__B1 _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8726_ as2650.stack\[3\]\[9\] _3848_ _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5938_ _1229_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4946__A3 _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8657_ as2650.stack\[6\]\[1\] _3800_ _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7345__A1 _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6148__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5869_ _4220_ _4125_ _1158_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7608_ as2650.addr_buff\[1\] _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7896__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8588_ _2779_ _0634_ _3640_ _3737_ _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7539_ _2160_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7235__C _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7648__A2 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8845__A1 _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput12 net12 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput23 net23 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9209_ _0158_ clknet_leaf_6_wb_clk_i as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput45 net45 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4882__A2 _4347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6084__A1 _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_0__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7820__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9022__A1 _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7033__B1 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8376__A3 _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7336__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7336__B2 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__I _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4570__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6847__B1 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4873__A2 _4453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8064__A2 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_3__f_wb_clk_i clknet_0_wb_clk_i clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6075__A1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5822__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6910_ _2121_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__9013__A1 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7890_ _3066_ _2284_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6841_ _2052_ _2067_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_62_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7575__A1 _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6378__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4804__I _4373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6772_ _1999_ _2000_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5050__A2 _4475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8511_ _4251_ _3664_ _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5723_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8442_ _0781_ _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5654_ as2650.pc\[9\] _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7878__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4605_ _4126_ _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8373_ _3531_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5635__I _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5585_ _4477_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7324_ _1545_ _2522_ _2524_ _2421_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4536_ _4115_ _4116_ _4117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _2447_ _2456_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__A2 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ _0736_ _1489_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_132_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7186_ _4446_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4864__A2 _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8055__A2 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _1418_ _1421_ _1422_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__A2 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ as2650.psl\[7\] _4150_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6861__I0 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8681__I _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9004__A1 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5019_ as2650.ins_reg\[4\] _4262_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7297__I _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7566__B2 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8709_ as2650.stack\[4\]\[10\] _3836_ _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7318__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8630__B _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8818__B2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8856__I _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8046__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6057__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_4_0_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_opt_4_0_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7557__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5883__C _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8521__A3 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6532__A2 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8809__A1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _0491_ _0704_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8285__A2 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6296__A1 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7040_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8991_ _1669_ _4017_ _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7796__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ _2797_ _3113_ _3116_ _3104_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__I3 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8434__C _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout47_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7873_ _4444_ _4408_ _2361_ _2187_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6824_ _2028_ _2029_ _2044_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6220__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5023__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6220__B2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6755_ _1968_ _1984_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ _0332_ _0946_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ _1826_ _1850_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8425_ _2903_ _3581_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5637_ _0944_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7720__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8356_ _0966_ _1110_ _3456_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5568_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7307_ _1555_ _2358_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8676__I _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8276__A2 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8287_ _1112_ _3448_ _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5499_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6287__A1 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7238_ net7 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8028__A2 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4709__I _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7169_ _1446_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6039__A1 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7787__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8200__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5275__I _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6514__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6278__A1 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9120__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4828__A2 _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8019__A2 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7778__A1 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9270__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__I _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__A1 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ as2650.idx_ctrl\[1\] _4451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6540_ _0744_ _0960_ _1038_ _4316_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4764__A1 _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6471_ _1715_ _1735_ _1736_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7702__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__A2 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8210_ _1590_ as2650.stack\[3\]\[4\] as2650.stack\[2\]\[4\] _0377_ _3241_ _3375_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_5422_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9190_ _0139_ clknet_leaf_25_wb_clk_i net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8141_ _3218_ _3306_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8258__A2 _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5353_ _0542_ _0643_ _0688_ _0321_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8072_ _3204_ _3239_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5284_ _0294_ _4312_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4819__A2 _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7023_ net22 _2228_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7769__A1 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8430__A2 _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8974_ _1683_ _2195_ _4040_ _4041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5244__A2 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7925_ _3100_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7856_ _2327_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8194__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6807_ _2009_ _2034_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7787_ _1633_ _2976_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7941__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6744__A2 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _4385_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4755__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _1965_ _1966_ _1967_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _1900_ _1901_ _1903_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8497__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8408_ _1395_ _3555_ _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8400__S _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9143__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7524__B _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6919__I _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8249__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8339_ _2991_ _3486_ _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5483__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8074__C _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5235__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__B1 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8488__A2 _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_17_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7160__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5733__I _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8249__C _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6671__A1 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8412__A2 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5226__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5971_ _0485_ _1253_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7710_ _2617_ _2892_ _2901_ _2370_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4922_ _4354_ _4503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8690_ _3823_ _3815_ _3824_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7641_ _2830_ _2834_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7609__B _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4853_ as2650.addr_buff\[6\] _4434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7395__I _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7923__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5908__I _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4737__A1 _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7572_ _2426_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9166__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4784_ _4303_ _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9311_ _0260_ clknet_leaf_17_wb_clk_i net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _1778_ _1787_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9242_ _0191_ clknet_leaf_3_wb_clk_i as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6454_ _1707_ _1721_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7151__A2 _4459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _4436_ _0662_ _0737_ _0470_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5162__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9173_ _0122_ clknet_leaf_44_wb_clk_i as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5162__B2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6385_ _4216_ _1660_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8124_ as2650.stack\[7\]\[2\] _3243_ _0501_ _3290_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5336_ _0667_ _0568_ _0669_ _0670_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__8100__A1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8055_ _2596_ _3221_ _3222_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5267_ _4286_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7006_ _4202_ _1463_ _2208_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ _0532_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8957_ _4490_ _3444_ _4019_ _3047_ _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_71_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7908_ _3078_ _3083_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8888_ _1102_ _3958_ _3967_ _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7839_ _0783_ _2999_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7914__A1 _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7678__B1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7254__B _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6649__I _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8069__C _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5456__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5221__C _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8158__A1 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6708__A2 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5728__I _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7905__A1 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A1 _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5392__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7943__I _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8330__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6892__A1 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5695__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6170_ _0931_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5121_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5052_ as2650.stack\[7\]\[9\] _4484_ _4489_ _0390_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_111_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8811_ as2650.r123\[1\]\[5\] _3901_ _3898_ _1792_ _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5131__C _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8742_ _1888_ _3856_ _3858_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5954_ _0313_ _1228_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_81_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8149__A1 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4905_ as2650.psu\[2\] _4486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8673_ _0976_ _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5885_ _4170_ _1157_ _1178_ _4284_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_61_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5638__I _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7624_ _2816_ _2817_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8014__I _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4836_ _4356_ _4371_ _4415_ _4416_ _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7372__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7555_ as2650.pc\[8\] _1595_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7911__A4 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5383__A1 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ _4289_ _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6506_ _1728_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7486_ _2678_ _2679_ _2683_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8321__A1 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7124__A2 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4698_ _4272_ _4278_ _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_140_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9225_ _0174_ clknet_3_6__leaf_wb_clk_i as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5135__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6437_ _1704_ _1706_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6883__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9156_ _0105_ clknet_leaf_45_wb_clk_i as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6883__B2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6368_ _1645_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8107_ _3273_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5319_ _4147_ _4149_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9087_ _0036_ clknet_leaf_58_wb_clk_i as2650.r123_2\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8624__A2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6299_ net27 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8617__C _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7521__C _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8038_ _3203_ _4472_ _3204_ _3206_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4717__I _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9331__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8927__A3 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4949__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7363__A2 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8560__A1 _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8859__I _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5913__A3 _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2__f_wb_clk_i clknet_0_wb_clk_i clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6626__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7431__C _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5232__B _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__I _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8379__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9040__A2 _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6929__A2 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5458__I _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_32_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_32_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _0996_ _0965_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5365__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4621_ _4184_ _4201_ _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5365__B2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5904__A3 _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7340_ _2539_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4552_ _4132_ _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8303__A1 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8303__B2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6289__I _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6314__B1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7271_ _2331_ _0935_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9204__CLK clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6314__C2 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8854__A2 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9010_ _2317_ _3012_ _4072_ _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__S1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _1166_ _1506_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6153_ _1183_ _1434_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5104_ as2650.r0\[3\] _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6084_ _4292_ _4199_ _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_131_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6093__A2 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _4348_ _0313_ _0322_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__4723__S0 _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _2191_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8790__B2 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8725_ _3843_ _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5937_ _1197_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4800__B1 _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8656_ _1888_ _3799_ _3801_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _1160_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7345__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8542__B2 _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7607_ _2629_ _2801_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4819_ _4399_ _4395_ _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8587_ _2362_ _0643_ _2439_ _3736_ _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5799_ _1089_ _1115_ _1116_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7538_ _2161_ _2733_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7469_ _1105_ _1597_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8845__A2 _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput13 net47 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput24 net24 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9208_ _0157_ clknet_leaf_3_wb_clk_i as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput35 net35 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6927__I _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9139_ _0088_ clknet_leaf_51_wb_clk_i as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6608__A1 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5052__B _4489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7281__A1 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6084__A2 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8363__B _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7033__A1 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6662__I _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8781__A1 _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7336__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8533__A1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5347__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9227__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7493__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6847__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8538__B _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5741__I _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6075__A2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5822__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7024__A1 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6840_ _2053_ _2066_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_63_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8772__A1 as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6771_ _1968_ _1984_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5188__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8510_ _2333_ _4263_ _4424_ _3663_ _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _0919_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8441_ _1018_ _3300_ _3596_ _3597_ _3122_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5653_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5889__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _4184_ _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8372_ _0998_ _3508_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5584_ _0858_ _0603_ _0864_ _0916_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7323_ _2523_ _2323_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4535_ net5 _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7254_ _1552_ _2394_ _2455_ _2135_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6205_ _0313_ _0437_ _0814_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7185_ _2353_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5651__I _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6136_ _1389_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7263__A1 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6067_ _4362_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5018_ _4306_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_73_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5577__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5098__I _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6969_ _1585_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8708_ _3818_ _3833_ _3837_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7318__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8515__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8639_ _3784_ _3785_ _3641_ _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4730__I _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8279__B1 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8358__B _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5501__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__I _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7006__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__I as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7557__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8754__A1 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8506__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4640__I _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A2 _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8809__A2 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6296__A2 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7245__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8990_ _1478_ _3503_ _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7941_ _3114_ _3115_ _3107_ _2917_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4815__I _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7872_ _2215_ _3049_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8745__A1 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5559__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6823_ _2023_ _2050_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6220__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6754_ _1971_ _1983_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5705_ _4270_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6685_ _1826_ _1850_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6251__B _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5646__I _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8022__I _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5636_ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8424_ as2650.addr_buff\[3\] _2333_ _2820_ _3493_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7720__A2 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8355_ _3066_ _3512_ _3514_ _3183_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5567_ net3 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7861__I _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7306_ _0556_ _0575_ _2506_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8286_ as2650.pc\[6\] _2593_ _3381_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7484__A1 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7237_ _1487_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5381__I _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7168_ _2318_ _2349_ _2371_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6119_ _1402_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7099_ _2292_ _2299_ _2302_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8984__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9072__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4725__I _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7101__I _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8200__A3 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5970__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7771__I _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7475__A1 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6387__I _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7720__B _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7227__B2 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7778__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4635__I _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8107__I _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6450__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8727__A1 _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8551__B _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7167__B _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5961__A1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _1734_ _1717_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8140_ _1083_ _3305_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5352_ _0323_ _0683_ _0687_ _4350_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7466__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6297__I _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8071_ _0493_ as2650.stack\[1\]\[1\] as2650.stack\[0\]\[1\] _3238_ _3239_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5283_ _0536_ _0617_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_134_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7022_ _2220_ _2223_ _2225_ _2227_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_101_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7218__A1 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8415__B1 _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4973__C _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7769__A2 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6246__B _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8973_ _4028_ _4033_ _4037_ _4039_ _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_55_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4545__I _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7924_ _2235_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8718__A1 _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7855_ _2230_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7856__I _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8194__A2 _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _0745_ _1023_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7786_ net49 _2967_ _1436_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4998_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6737_ _0744_ _1004_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4755__A2 _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6668_ as2650.stack\[3\]\[4\] _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8407_ _2531_ _3558_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5619_ _4122_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6599_ _1071_ _1856_ _1859_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__C _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8338_ _3274_ _3481_ _3498_ _3089_ _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7457__A1 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8269_ _1559_ _2528_ _3273_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6935__I _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8355__C _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8957__A1 _4490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8957__B2 _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5060__B _4517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7766__I _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6670__I _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__B2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4746__A2 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__I _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7715__B _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7696__A1 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8597__I _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5171__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_57_wb_clk_i clknet_opt_5_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6120__A1 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8546__B _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6671__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5970_ _4265_ _1170_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8963__A4 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4921_ _4464_ _4467_ _4501_ _4502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7640_ _2832_ _2833_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4852_ as2650.addr_buff\[6\] _4432_ _4433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7923__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7571_ _2765_ _2766_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4783_ _4362_ _4363_ _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4737__A2 _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5196__I _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5934__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9310_ _0259_ clknet_leaf_17_wb_clk_i net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6522_ _1782_ _1786_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7687__A1 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6453_ _1714_ _1720_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9241_ _0190_ clknet_leaf_67_wb_clk_i as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5404_ _0571_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9172_ _0121_ clknet_leaf_45_wb_clk_i as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5162__A2 as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6384_ _4511_ _1366_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_47_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7439__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8123_ _3288_ _4472_ _3204_ _3289_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5335_ _0670_ _0636_ _0552_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8100__A2 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8054_ _0352_ _2338_ _2216_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ as2650.r123\[0\]\[4\] _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7005_ _1446_ _1675_ _2210_ _2211_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5197_ _0432_ _0427_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8939__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8175__C _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8956_ _4018_ _4022_ _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7907_ _3079_ _2190_ _3082_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8887_ _1539_ _3959_ _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7838_ _0607_ _2997_ _3020_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9110__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7914__A2 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7769_ _1447_ _2287_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7678__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7678__B2 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9260__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7254__C _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4900__A2 _4474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_1__f_wb_clk_i clknet_0_wb_clk_i clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6665__I _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7850__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8085__C _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8880__I _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8158__A2 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4913__I as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7905__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5916__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5916__B2 _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7669__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7669__B2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8330__A2 _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8120__I _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6341__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5120_ _0341_ _0345_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8094__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8276__B _4498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5051_ _0382_ _0388_ _0389_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8810_ _3906_ _3907_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8936__A4 _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9133__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8741_ as2650.stack\[7\]\[0\] _3857_ _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__A2 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5953_ _0320_ _1232_ _1245_ _1227_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5080__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8149__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4823__I _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4904_ _4484_ _4485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5884_ _4171_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8672_ _1908_ _3805_ _3810_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7623_ net37 net36 _2746_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__9283__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4835_ _4230_ _4416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7554_ _2352_ _2743_ _2749_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6580__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5383__A2 _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _4298_ _4308_ _4346_ _4347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4979__B _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6505_ _1769_ _0647_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7485_ _2671_ _2324_ _2329_ _2682_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4697_ _4277_ _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8321__A2 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9224_ _0173_ clknet_leaf_32_wb_clk_i as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6436_ _1217_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9155_ _0104_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6367_ _0977_ _1647_ _1649_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8106_ _1443_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8085__A1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5318_ _0651_ _4165_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9086_ _0035_ clknet_leaf_58_wb_clk_i as2650.r123_2\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6298_ _0378_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7832__A1 _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8037_ _0493_ as2650.stack\[5\]\[0\] as2650.stack\[4\]\[0\] _3205_ _3206_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5249_ _0387_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_2_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8927__A4 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8939_ _0624_ _4006_ _1499_ _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4949__A2 _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7899__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6571__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5913__A4 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5126__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8875__I _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4908__I _4488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6626__A2 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9156__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7051__A2 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4643__I _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8000__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7954__I _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8551__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4620_ _4196_ _4200_ _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8839__B1 _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4551_ _4131_ _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7270_ _2341_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6314__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6314__B2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ _1492_ _1493_ _1499_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8067__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _4185_ _1436_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5103_ _0316_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7814__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ _0922_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5034_ _0323_ _0328_ _0372_ _4449_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_85_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4723__S1 _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8453__C _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6985_ _1362_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8790__A2 _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4553__I as2650.alu_op\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8724_ _3811_ _3845_ _3847_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _4441_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4800__A1 _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4800__B2 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8655_ as2650.stack\[6\]\[0\] _3800_ _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ _4441_ _4412_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8542__A2 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7606_ _2160_ as2650.addr_buff\[1\] _2730_ _2732_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4818_ _4211_ _4398_ _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8586_ _2983_ _0686_ _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5798_ as2650.stack\[1\]\[7\] _1094_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7085__B _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7537_ _2730_ _2732_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4749_ _4325_ _4329_ _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7468_ _2593_ _0755_ _2665_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xoutput14 net14 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9207_ _0156_ clknet_leaf_4_wb_clk_i as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput25 net25 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6419_ _4141_ _1673_ _1690_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput36 net36 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7399_ net33 _2597_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4867__A1 _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9179__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8628__C _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8058__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9138_ _0087_ clknet_leaf_52_wb_clk_i as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6608__A2 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__I _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7805__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9069_ _0018_ clknet_leaf_46_wb_clk_i as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7104__I _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4619__A1 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7281__A2 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6084__A3 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8230__A1 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7033__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8533__A2 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A1 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8297__A1 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7014__I _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7949__I _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7024__A2 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8221__A1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8772__A2 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6770_ _1971_ _1983_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5721_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8440_ _3078_ _3578_ _3166_ _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5652_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6535__A1 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ _4128_ _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8371_ _3123_ _3530_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5583_ _4290_ _0884_ _0915_ _4288_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7322_ net53 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4534_ _4114_ _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9321__CLK clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7253_ _2450_ _2453_ _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__A1 _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5897__I0 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6204_ _4347_ _0541_ _0633_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7184_ _4447_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5510__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _0651_ _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8460__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _1349_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _4450_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8212__A1 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8763__A2 _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6968_ _2178_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7971__B1 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8707_ as2650.stack\[4\]\[9\] _3836_ _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5919_ _4371_ _1199_ _1211_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6899_ as2650.stack\[4\]\[5\] _2115_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8638_ _3139_ _0891_ _2370_ _3785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7723__B1 _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8569_ _2273_ _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8279__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8279__B2 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5501__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6159__B _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5063__B _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8451__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5265__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6673__I _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8203__A1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7006__A2 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8203__B2 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7309__A3 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8506__A2 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6517__A1 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7190__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7009__I _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6296__A3 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8690__A1 _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7245__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5256__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5256__B2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8993__A2 _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7940_ _2217_ _1660_ _2968_ _3085_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7871_ _2993_ _3034_ _2225_ _3048_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6822_ _1915_ _2049_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5559__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _1978_ _1982_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5704_ as2650.pc\[14\] _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6508__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6684_ _1702_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6508__B2 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8423_ _1018_ _3579_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5635_ _0966_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8354_ _3066_ _3513_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4987__B _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5566_ _0666_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7305_ _2450_ _2451_ _2505_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5497_ _0830_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8285_ _1105_ _3341_ _3447_ _3254_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7484__A2 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6287__A3 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7236_ _1380_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5495__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7167_ _2352_ _2363_ _2369_ _2370_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8433__A1 _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6118_ _4133_ _4145_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8433__B2 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7098_ _4224_ _2301_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8984__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6049_ net3 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8922__B _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6747__A1 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5970__A2 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7172__A1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7172__B2 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5572__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8672__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5486__B2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6683__B1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8424__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7227__A2 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7720__C _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6986__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8727__A2 _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__A1 _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5747__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4651__I _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7167__C _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5961__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7163__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5420_ net1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6910__A1 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5351_ _4431_ _0686_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7466__A2 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8070_ _0379_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5282_ _0531_ _0616_ _0604_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_142_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5477__A1 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7021_ _2202_ _2226_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7218__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8415__A1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8415__B2 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5229__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8972_ _2949_ _3152_ _4038_ _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout52_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7923_ _0409_ _3086_ _3098_ _2280_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_82_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8718__A2 _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7854_ _3031_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6805_ _2012_ _2016_ _2032_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7785_ _2793_ _2970_ _2974_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4997_ _0333_ _4422_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4561__I as2650.alu_op\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8033__I _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _0611_ _0648_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6667_ _1890_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8406_ _2839_ _3563_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5618_ _4252_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6598_ as2650.stack\[5\]\[1\] _1857_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7093__B _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8337_ _3274_ _3497_ _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5549_ _4313_ _0876_ _0878_ _0620_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8103__B1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7457__A2 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_0__f_wb_clk_i clknet_0_wb_clk_i clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8268_ _0833_ _0747_ _3430_ _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_79_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7219_ _1465_ _2421_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8199_ _3350_ _3356_ _3363_ _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8406__A1 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8957__A2 _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4736__I _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8009__I1 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8709__A2 _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6951__I as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7917__B1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6196__A2 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9186__D _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7393__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5567__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7696__A2 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8893__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8645__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6120__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8546__C _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4646__I _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8948__A2 _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_26_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_26_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8562__B _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4920_ _4481_ _4491_ _4493_ _4500_ _4501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ as2650.addr_buff\[5\] _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7384__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6187__A2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7570_ _2751_ _2754_ _2764_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_127_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4782_ as2650.r123\[2\]\[7\] as2650.r123_2\[2\]\[7\] _4112_ _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5934__A2 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _1783_ _1784_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_53_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9240_ _0189_ clknet_leaf_67_wb_clk_i as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7687__A2 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8884__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6452_ _1715_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9062__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _0669_ _0660_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9171_ _0120_ clknet_leaf_55_wb_clk_i as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6383_ _1658_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8122_ _0493_ as2650.stack\[5\]\[2\] as2650.stack\[4\]\[2\] _3205_ _3289_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7439__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5334_ _0355_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8636__A1 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8053_ _0351_ _4380_ _3220_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5265_ _0511_ _4287_ _0601_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5940__I _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7004_ _1324_ _1363_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5196_ _0419_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4556__I _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8955_ _4466_ _4499_ _4021_ _2226_ _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5622__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7906_ _2190_ _2198_ _3081_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8886_ _3957_ _3965_ _3966_ _3953_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_93_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7837_ _2998_ _3019_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7375__A1 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7768_ _1466_ _2957_ _1183_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6719_ _1926_ _1949_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7699_ as2650.pc\[12\] _0831_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7678__A2 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7107__I _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8627__A1 _4508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6946__I _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7850__A2 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7777__I _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9085__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8866__A1 _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6341__A2 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7017__I _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8618__A1 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6856__I _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8094__A2 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5760__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5050_ as2650.stack\[6\]\[9\] _4475_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5852__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9043__A1 _4515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8740_ _3855_ _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5952_ _1242_ _1244_ _1232_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5080__A2 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4903_ _4483_ _4484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8671_ as2650.stack\[6\]\[7\] _3806_ _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5883_ _4204_ _1158_ _1162_ _1176_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_107_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7622_ net52 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4834_ _4374_ _4384_ _4402_ _4414_ _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5000__I _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7553_ _2365_ _2747_ _2748_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _4313_ _4331_ _4345_ _4346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8306__B1 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6504_ _0342_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7355__C _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8857__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7484_ _2321_ _2681_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4696_ _4276_ _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9223_ _0172_ clknet_leaf_23_wb_clk_i as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6868__B1 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _1697_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9154_ _0103_ clknet_leaf_54_wb_clk_i as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8609__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6366_ as2650.stack\[6\]\[8\] _1648_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8105_ _3263_ _3265_ _3271_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5317_ _4361_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8085__A2 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9085_ _0034_ clknet_leaf_59_wb_clk_i as2650.r123_2\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6297_ _0933_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6096__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8036_ _0379_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7832__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _0494_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9034__A1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5179_ _0445_ _0447_ _0449_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_68_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8938_ _1503_ _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8869_ _3551_ _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8930__B _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__A1 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6571__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__A3 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7520__A1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6676__I _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9025__A1 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7587__A1 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6344__C _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8000__A2 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8839__A1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4550_ _4130_ _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7511__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6314__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ _1492_ _1493_ _1499_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6865__A3 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6151_ _1435_ _4200_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9100__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5102_ _4356_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7814__A2 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6082_ _4390_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9016__A1 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5033_ _0323_ _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7578__A1 _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7578__B2 _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9250__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6984_ _1206_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8723_ as2650.stack\[3\]\[8\] _3846_ _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5935_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_80_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4800__A2 _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8654_ _3798_ _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5866_ _1159_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6002__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7605_ _2162_ _2741_ _2165_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _4397_ _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8585_ _3014_ _3683_ _3735_ _3552_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5797_ _1114_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8041__I _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7536_ _4428_ _2731_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4748_ _4308_ _4327_ _4328_ _4329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_108_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7467_ _1096_ _1584_ _2619_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7502__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ _4259_ _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9206_ _0155_ clknet_leaf_3_wb_clk_i as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6418_ _1689_ _1684_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput15 net15 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput26 net26 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7398_ net32 _2567_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xoutput37 net37 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4867__A2 _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8058__A2 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9137_ _0086_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6349_ _0970_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9068_ _0017_ clknet_leaf_56_wb_clk_i as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7805__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5816__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4619__A2 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8019_ _2412_ _3186_ _3187_ _3036_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9007__A1 _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8230__A2 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7120__I _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6241__A1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8781__A3 _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7741__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8297__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9123__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4858__A2 _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5243__C _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9273__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4654__I as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8221__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5686__S _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7980__A1 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5720_ _0393_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5651_ _0981_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6535__A2 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7732__A1 _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4546__A1 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _4155_ _4182_ _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8370_ _2777_ _3303_ _3529_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5582_ _4290_ _0914_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7321_ _2514_ _2521_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7914__B _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4533_ as2650.halted _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7496__B1 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7252_ _2450_ _2453_ _2357_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__A2 _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6203_ _1487_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5897__I1 _4501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7183_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6134_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7799__A1 _4452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5649__I1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8460__A2 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A2 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6471__B2 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5016_ as2650.ins_reg\[4\] _4407_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8212__A2 _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6223__A1 _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _2176_ _2177_ _2174_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7971__A1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8706_ _3831_ _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5918_ _1160_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6898_ _1900_ _2114_ _2116_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8515__A3 _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8637_ _3701_ _0894_ _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5849_ as2650.stack\[1\]\[10\] _1146_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7723__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7723__B2 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__A1 _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8568_ _4409_ _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7519_ _0933_ _0891_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_135_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8279__A2 as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8499_ _3645_ _3651_ _3652_ _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9296__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4739__I _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7115__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6159__C _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6954__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8203__A2 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7006__A3 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6214__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8506__A3 _4514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7714__A1 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5254__B _4490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8690__A2 _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7025__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8284__C _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7870_ _2839_ _3042_ _3046_ _3047_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6205__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6821_ _2025_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_91_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7953__A1 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ _1980_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9169__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5703_ _0978_ _1028_ _1029_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6683_ _1217_ _1911_ _1913_ as2650.r123_2\[2\]\[0\] _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7705__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6508__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7705__B2 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8422_ _2855_ _2814_ _3533_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5634_ as2650.pc\[8\] _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8353_ _2803_ _3496_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5565_ _4370_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5943__I _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8459__C _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7304_ _0454_ _0475_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8284_ _3095_ _3416_ _3436_ _3446_ _3299_ _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5496_ net2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7235_ _2379_ _2433_ _2435_ _2437_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_137_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6692__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7166_ _1487_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6117_ _0691_ _0692_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_140_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8433__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7097_ _2259_ _2300_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6444__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _0863_ _1186_ _1180_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8197__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7999_ _2939_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5955__B1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8369__C _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4930__A1 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__A4 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5486__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6683__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6683__B2 as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8424__A2 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6986__A2 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4997__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8188__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9311__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7935__A1 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5961__A3 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7163__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8360__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6910__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8279__C _4488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5350_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4921__A1 _4464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ _0531_ _0604_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6674__A1 as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5477__A2 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7020_ _1638_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7871__B1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6594__I _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8415__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__A1 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8966__A3 _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8971_ _1351_ _1374_ _2193_ _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4988__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7922_ _1349_ _3097_ _0334_ _1471_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__5003__I as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8179__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7853_ _2220_ _2230_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7926__A1 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4842__I _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6804_ _2004_ _2031_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7784_ net49 _2967_ _2971_ _2973_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4996_ _4131_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6735_ _1936_ _1937_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6666_ _1890_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8405_ _3347_ _3555_ _3562_ _1639_ _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5165__A1 _4494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ _4238_ _4189_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5165__B2 _4476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6597_ _1062_ _1856_ _1858_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6901__A2 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8336_ _3495_ _3496_ _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4912__A1 _4474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5548_ _4341_ _0879_ _0872_ _0431_ _0880_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8103__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_3_0_wb_clk_i clknet_3_3__leaf_wb_clk_i clknet_opt_3_0_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8103__B2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8267_ _3428_ _3387_ _3429_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5479_ _0306_ _0801_ _0812_ _0311_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7218_ _2420_ _1663_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8198_ _3357_ _3345_ _3359_ _3360_ _3362_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5622__B _4421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7149_ _2126_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7614__B1 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9334__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7090__A1 _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4979__A1 _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7917__B2 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8590__A1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout50 net26 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8645__A2 _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9004__B _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7081__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_wb_clk_i clknet_opt_1_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7908__A1 _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__I as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _4430_ _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7384__A2 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8581__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4781_ _4361_ _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7973__I as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6520_ _0442_ _1752_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8333__A1 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _1716_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6589__I _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9207__CLK clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5493__I _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ _0668_ _0660_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9170_ _0119_ clknet_leaf_55_wb_clk_i as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6382_ _4405_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8121_ as2650.stack\[6\]\[2\] _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5333_ _0558_ _0516_ _0609_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_138_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8636__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8052_ net6 _4302_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5264_ _0512_ _0583_ _0600_ _0401_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7003_ _2209_ _2192_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5195_ _0531_ _0523_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7072__A1 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8954_ _0972_ _4019_ _4020_ _4466_ _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5622__A2 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7905_ _2967_ _1398_ _3080_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8885_ net19 _3962_ _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5668__I _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4572__I as2650.alu_op\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7836_ _1090_ _3009_ _3018_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_63_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7375__A2 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8572__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4979_ _4450_ _4454_ _0317_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7767_ _2956_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6718_ _1932_ _1948_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7698_ _2833_ _2887_ _2889_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8324__A1 _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6649_ _1061_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7832__B _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8319_ _0967_ _3479_ _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9299_ _0248_ clknet_leaf_1_wb_clk_i as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8627__A2 _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5310__A1 _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7123__I _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6962__I _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7063__A1 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8260__B1 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6810__A1 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8563__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8315__A1 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6326__B1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6202__I _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8079__B1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8618__A2 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8557__C _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5301__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5852__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9043__A2 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7968__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7054__A1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__A2 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _0328_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4902_ _4482_ _4483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8670_ _1906_ _3805_ _3809_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5882_ _1165_ _1171_ _1174_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__8554__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7621_ _2814_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5368__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4833_ _4413_ _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5368__B2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7552_ _2405_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4764_ _4334_ _4337_ _4344_ _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8306__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8306__B2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _1749_ _1758_ _1767_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7483_ _2667_ _2680_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4591__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4695_ _4275_ _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7208__I _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6868__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6112__I _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9222_ _0171_ clknet_leaf_23_wb_clk_i as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6434_ as2650.r123_2\[1\]\[0\] _1699_ _1701_ _1703_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9153_ _0102_ clknet_leaf_54_wb_clk_i as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6365_ _1646_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8609__A2 _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8104_ _3266_ _3258_ _3267_ _3270_ _3068_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8467__C _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5316_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _4111_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9084_ _0033_ clknet_leaf_66_wb_clk_i as2650.r123_2\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6296_ _1454_ _1579_ _1521_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5172__B _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8035_ _3194_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6096__A2 _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _0381_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5178_ as2650.holding_reg\[3\] _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__9034__A2 _4515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__A1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8242__B1 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7596__A2 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8793__A1 _4463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7099__B _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8937_ _3989_ _4004_ _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8868_ net43 _3945_ _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7348__A2 _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8545__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5359__A1 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7819_ _1680_ _1639_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8799_ as2650.r123\[1\]\[2\] _3889_ _3898_ _1722_ _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8848__A2 _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7118__I _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5531__A1 _4517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__I _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7284__A1 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9025__A2 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7036__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8784__A1 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6795__B1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9052__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5101__I _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6011__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8839__A2 _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7028__I _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6150_ _4143_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6088__B _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7275__A1 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6078__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8472__B1 _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_135_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _0331_ _0337_ _0366_ _0370_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9016__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7027__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_10_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_10_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8775__A1 _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7822__I0 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6983_ _1436_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8722_ _3844_ _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5011__I _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ _4265_ _1170_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8527__A1 _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8527__B2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8653_ _3798_ _3799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5865_ _4186_ _4229_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4850__I _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7604_ _2388_ _2798_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4816_ _4305_ _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5796_ _0862_ _1081_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8584_ _2239_ _3730_ _3731_ _3734_ _3735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7535_ _1336_ _0894_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4747_ _4322_ _4320_ _4328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4564__A2 _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7466_ _2558_ _2560_ _2607_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4678_ _4258_ _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6417_ _1560_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9205_ _0154_ clknet_leaf_6_wb_clk_i as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5513__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7397_ _4256_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput16 net16 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput27 net27 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput38 net38 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9136_ _0085_ clknet_leaf_61_wb_clk_i as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6348_ _1631_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7266__A1 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6069__A2 _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9067_ _0016_ clknet_leaf_56_wb_clk_i as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6279_ _1324_ _1419_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5816__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8018_ _2311_ _1659_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9007__A2 _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7401__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7569__A2 _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8766__A1 as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4961__S _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6241__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8518__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4760__I _4340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__B1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5504__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7257__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8757__A1 as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5991__A1 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4670__I _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5650_ _0980_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7732__A2 _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _4181_ _4182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5581_ _0542_ _0891_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4546__A2 _4126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7320_ _2515_ _2520_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_129_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4532_ _4112_ _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7914__C _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7496__A1 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7251_ _2451_ _2452_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7496__B2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ _1486_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4849__A3 _4429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7182_ _1451_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9098__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _0333_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7799__A2 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8996__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _0333_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__I as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5015_ _4395_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6471__A2 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8748__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7420__A1 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6966_ as2650.addr_buff\[4\] _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7971__A2 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8705_ _3811_ _3833_ _3835_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ _1200_ _1201_ _1202_ _1210_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5676__I _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5982__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6897_ as2650.stack\[4\]\[4\] _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8636_ _3079_ _0884_ _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _0990_ _1143_ _1147_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7723__A2 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6526__A3 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8920__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4537__A2 _4117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7891__I _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8567_ _3689_ _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5779_ _0784_ _1081_ _1098_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7518_ _2656_ _2659_ _2714_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8498_ _1519_ _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7487__A1 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7487__B2 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7449_ _1103_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8001__B _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6300__I _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7239__A1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9119_ _0068_ clknet_leaf_5_wb_clk_i as2650.alu_op\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8987__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6998__B1 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7411__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8390__C _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8506__A4 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7714__A2 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8911__A1 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8897__I _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7478__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8978__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7650__A1 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6205__A2 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6820_ _2046_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6751_ _0443_ _1769_ _1979_ _1039_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5964__A1 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ as2650.stack\[2\]\[13\] _0957_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6682_ _1912_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8902__A1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8421_ _3577_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5633_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5716__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8352_ _3511_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5564_ _0895_ _0752_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7469__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7303_ _2498_ _2502_ _2503_ _2127_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8283_ _3212_ _3445_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5495_ _0792_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7234_ _2436_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7165_ _2337_ _2365_ _2368_ _2325_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6692__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _0946_ _1401_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7096_ _4133_ _4145_ _1353_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6444__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6047_ as2650.r123_2\[0\]\[7\] _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7886__I _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8197__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ _3166_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9113__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7944__A2 _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6949_ _2162_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8619_ _3682_ _3767_ _2230_ _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9263__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6380__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4930__A2 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6132__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6965__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7880__A1 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8424__A3 _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7632__A1 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4997__A2 _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8188__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6199__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5946__B2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7699__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8360__A2 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6371__A1 as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4921__A2 _4467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ _0606_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6123__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6674__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7871__A1 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4685__A1 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7623__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6426__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8970_ _1433_ _4034_ _4035_ _4036_ _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_67_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9136__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7921_ _1420_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4988__A2 _4522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8179__A2 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7852_ _3030_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7926__A2 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6803_ _2011_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7783_ _2413_ _2972_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4995_ _4217_ _4228_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _1962_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6665_ _1092_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8404_ _3536_ _3557_ _3561_ _2935_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5616_ _0925_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6596_ as2650.stack\[5\]\[0\] _1857_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8335_ _2160_ _2475_ _3493_ _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_69_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5547_ _4295_ _0873_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8103__A2 _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8266_ _2606_ _0652_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5478_ _0309_ _0800_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7390__B _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7217_ _0932_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7862__A1 _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8197_ _2150_ _3361_ _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7148_ _2351_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7614__A1 _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7614__B2 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7079_ _4194_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7090__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7917__A2 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__B1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8590__A2 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout51 net40 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7565__B _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6353__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6105__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7853__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9159__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6120__A4 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9004__C _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__A1 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5104__I as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7081__A2 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5092__A1 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7369__B1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5919__A1 _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6967__I0 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8581__A2 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4780_ _4300_ _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6450_ _4299_ _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6344__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5401_ _0726_ _0734_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6381_ _1621_ _1456_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8120_ _3077_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5332_ _4450_ _0639_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8051_ _3218_ _3217_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5263_ _0375_ _0597_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7844__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7002_ _1475_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5442__C _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5194_ _0522_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5014__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7072__A2 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8953_ _0439_ _0972_ _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4853__I as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7904_ _0927_ _2283_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8884_ _0784_ _3958_ _3964_ _3965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4830__A1 _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7835_ _2176_ _2226_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8572__A2 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7766_ _2272_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4978_ _4451_ _4453_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6717_ _1935_ _1947_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7697_ _2866_ _2831_ _2888_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8324__A2 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6648_ _1887_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6579_ as2650.r0\[6\] _0980_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8318_ _1111_ _3448_ _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9301__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9298_ _0247_ clknet_leaf_1_wb_clk_i as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7835__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8249_ _3168_ _3382_ _3412_ _3299_ _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4649__A1 _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5310__A2 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8944__B _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8260__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7063__A2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8260__B2 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5859__I as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6810__A2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4821__A1 _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8012__A1 _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5594__I _4404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6326__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__B2 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8079__A1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9015__B _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7826__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__A2 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5769__I _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6801__A2 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5950_ _4248_ _1173_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_46_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8003__A1 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ as2650.psu\[0\] as2650.psu\[1\] _4482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5881_ _4268_ _4446_ _1173_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8554__A2 _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7620_ as2650.pc\[10\] _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4832_ _4403_ _4412_ _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7917__C _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6565__A1 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7551_ _2744_ _2746_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_92_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4763_ _4338_ _4330_ _4343_ _4297_ _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8306__A2 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _1750_ _1757_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7482_ _2608_ _2581_ _2618_ _2666_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4694_ _4274_ _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9324__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9221_ _0170_ clknet_leaf_42_wb_clk_i as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6433_ _1702_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6868__A2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4879__A1 _4449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5009__I _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9152_ _0101_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6364_ _1646_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8103_ _1552_ _2778_ _2961_ _3257_ _3269_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5315_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_66_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9083_ _0032_ clknet_leaf_57_wb_clk_i as2650.r123_2\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6295_ _1458_ _4333_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7293__A2 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8034_ as2650.stack\[6\]\[0\] _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6096__A3 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5246_ _0410_ _0541_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5177_ _0422_ _0450_ _0513_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9034__A3 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8242__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5679__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5056__A1 as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8793__A2 _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8936_ _3991_ _3996_ _3999_ _4003_ _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8867_ _0506_ _3941_ _3950_ _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7818_ _1395_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5359__A2 _4506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8798_ _3890_ _3898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7749_ _2939_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8939__B _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5531__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7808__A1 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7808__B2 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7134__I _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7284__A2 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8481__A1 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8233__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7036__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5589__I _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8784__A2 _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6795__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5522__A2 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6088__C _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ _0414_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7275__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8472__A1 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _4367_ _4150_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _4215_ _0368_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7027__A2 _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5499__I _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8775__A2 _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7822__I1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6982_ net24 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6786__A1 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8721_ _3844_ _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _0398_ _1223_ _1225_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_50_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8527__A2 _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8652_ _1889_ _1854_ _1118_ _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_59_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5864_ _4177_ _1156_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7603_ _2161_ _2165_ _2741_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4815_ _4395_ _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8583_ _3639_ _0541_ _3641_ _3733_ _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5795_ _1112_ _0974_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7534_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4746_ _4274_ _4306_ _4326_ _4327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7465_ _2648_ _2655_ _2662_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5962__I _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4677_ as2650.idx_ctrl\[1\] as2650.idx_ctrl\[0\] _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9204_ _0153_ clknet_leaf_4_wb_clk_i as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6416_ _4311_ _1687_ _1688_ _1668_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ _2594_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput17 net17 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput28 net28 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9135_ _0084_ clknet_leaf_61_wb_clk_i as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput39 net39 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6347_ _1476_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7266__A2 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9066_ _0015_ clknet_leaf_56_wb_clk_i as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _1513_ _1542_ _1547_ _1562_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7889__I _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5277__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8017_ _1203_ _3185_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5229_ _0543_ _4355_ _0565_ _4352_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9007__A3 _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8215__A1 _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8766__A2 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6777__A1 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8919_ _2176_ _1686_ _3988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8518__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_112_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6529__A1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7129__I _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__B2 _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5872__I _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7257__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8206__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6768__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5440__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5440__B2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7193__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8390__B1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4600_ _4137_ _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5580_ _0314_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6940__A1 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6878__I _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4531_ _4111_ _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7496__A2 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7250_ _0456_ _0476_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8693__A1 _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6201_ _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7181_ _2383_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _1411_ _1413_ _1414_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8996__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6063_ _4226_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5014_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7420__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _0677_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5957__I as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8704_ as2650.stack\[4\]\[8\] _3834_ _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ _1203_ _1205_ _1208_ _4399_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _2107_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8635_ _0862_ _3680_ _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5847_ as2650.stack\[1\]\[9\] _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8920__A2 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8566_ _1254_ _3683_ _3717_ _3552_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5778_ _1097_ _1059_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6931__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8489__B _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7517_ _0831_ _0821_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4729_ _4309_ _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8497_ _3647_ _0962_ _3650_ _4169_ _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7448_ _2434_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7487__A2 _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8684__A1 _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7379_ _1558_ _2577_ _2568_ _2578_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_122_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8436__A1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9118_ _0067_ clknet_leaf_5_wb_clk_i as2650.alu_op\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8436__B2 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8987__A2 _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9049_ _3016_ _4103_ _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6998__A1 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6998__B2 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5670__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7411__A2 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4771__I _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4704__C _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7175__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6922__A1 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7478__A2 _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5535__C _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8427__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4700__A3 _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6989__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5661__A1 as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6205__A3 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5777__I _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5413__A1 _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7197__C _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6750_ _1769_ _1979_ _1039_ _0444_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5701_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _1693_ _1694_ _1910_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8420_ _1017_ _3576_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8902__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5632_ _0963_ _0947_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6913__A1 _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8351_ _3508_ _3510_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9065__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5563_ _4212_ _0817_ _0752_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7302_ _1556_ _2498_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6401__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7469__A2 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8282_ _2241_ _3416_ _3443_ _3444_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5494_ _0759_ _0760_ _0662_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7941__B _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7233_ _1693_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5017__I _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7164_ _2367_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6115_ _4171_ _1400_ _1348_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8969__A2 _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7095_ _4206_ _2298_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _1317_ _1286_ _1333_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7997_ _3165_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5687__I _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8063__I _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _2158_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4758__A3 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6879_ _2088_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8618_ _3747_ _3684_ _3756_ _3766_ _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6904__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8549_ _2983_ _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7407__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6380__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6311__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6132__A2 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8409__A1 _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7880__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5371__B _4490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7142__I _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7632__A2 _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5643__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A3 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7298__B _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6199__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9088__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8701__I _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7699__A2 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6371__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8648__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4921__A3 _4501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7761__B _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6123__A2 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8576__C _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7871__A2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4685__A2 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__I _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7623__A2 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8820__A1 _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7920_ _3084_ _3094_ _3095_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7851_ _2231_ _3029_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6802_ _2028_ _2029_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7782_ _0948_ _2968_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4994_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6733_ _1932_ _1948_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7139__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7655__C _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8887__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6664_ _1898_ _1891_ _1899_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8403_ _2315_ _3554_ _3558_ _3419_ _3560_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5615_ _0945_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6595_ _1855_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6131__I _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8334_ _2735_ _3494_ _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5546_ _0871_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7671__B _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8265_ _2606_ _0652_ _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7311__A1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ _4310_ _0798_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7216_ _0970_ _2418_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8196_ _0677_ _2206_ _2130_ as2650.addr_buff\[4\] _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7862__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5873__A1 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7147_ _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7614__A2 _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7078_ _0405_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8811__B2 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_5__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ as2650.r123_2\[0\]\[6\] _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7090__A3 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9230__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6050__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__B2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout52 net38 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8878__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6353__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5085__C _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7581__B _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6976__I _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7302__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6105__A2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7853__A2 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5864__A1 _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5092__A2 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7369__B2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_90 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__6967__I1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6344__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ _0436_ _0729_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6380_ _1043_ _1648_ _1656_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8587__B _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6886__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5331_ _4136_ _4262_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8097__A2 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8050_ _2193_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5262_ _0598_ _0507_ _4516_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7844__A2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4658__A2 as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7001_ _2207_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_130_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9046__A1 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _4334_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5607__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9253__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8952_ _4494_ _3331_ _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6280__A1 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout50_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7903_ _2339_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8883_ _3747_ _3959_ _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4830__A2 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7834_ _0515_ _2997_ _3017_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6032__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6032__B2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7765_ _1631_ _2949_ _2954_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4977_ _4522_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6716_ _1938_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7696_ as2650.pc\[11\] _0831_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6647_ as2650.r123\[3\]\[7\] _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7532__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6578_ _1753_ _1839_ _1840_ _1809_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_69_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8317_ _1112_ _3341_ _3477_ _3478_ _3122_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5529_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9297_ _0246_ clknet_leaf_1_wb_clk_i as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8248_ _3403_ _3411_ _3251_ _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7835__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8179_ _1083_ _3305_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5205__I _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7599__A1 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5074__A2 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6036__I _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5096__B _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8079__A2 _4471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5316__S _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9015__C _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7826__A2 _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9276__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5115__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9031__B _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4954__I _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7330__I _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6262__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4812__A2 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ as2650.stack\[6\]\[8\] _4474_ _4480_ _4481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8003__A2 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ _4247_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__A1 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _4406_ _4409_ _4411_ _4412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__I _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6565__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8161__I _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7550_ _2745_ _2691_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4576__A1 _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4762_ _4339_ _4341_ _4342_ _4329_ _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6501_ _1746_ _1760_ _1765_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7481_ _2671_ _2472_ _2577_ _1559_ _2346_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__7514__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6317__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4693_ _4273_ _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9220_ _0169_ clknet_leaf_23_wb_clk_i as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6432_ _1694_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4879__A2 _4459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9151_ _0100_ clknet_leaf_58_wb_clk_i as2650.r123\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6363_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8102_ _1155_ _3268_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5314_ as2650.r0\[5\] _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9082_ _0031_ clknet_leaf_58_wb_clk_i as2650.r123_2\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6294_ _4151_ _1370_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8033_ _0380_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9019__A1 _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5245_ _0542_ _0577_ _0581_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7293__A3 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6096__A4 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8490__A2 _4347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ as2650.holding_reg\[3\] _4161_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9034__A4 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8242__A2 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5056__A2 _4473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8935_ _1564_ _2235_ _2254_ _4002_ _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_43_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8866_ _3690_ _3942_ _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6005__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7817_ _1065_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8797_ _3896_ _3897_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7753__A1 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7748_ _2244_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7679_ _2578_ _2859_ _2871_ _2695_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7505__A1 _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6308__A2 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9299__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7808__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__A2 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4774__I _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8233__A2 _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7150__I _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6244__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7441__B1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7992__A1 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7325__I _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8472__A2 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6483__A1 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8584__C _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5030_ _0336_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8224__A2 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7060__I _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6981_ _2186_ _2163_ _2188_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6786__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7983__A1 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5932_ _1065_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8720_ _3843_ _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8651_ _1644_ _3782_ _3797_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_62_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ _1155_ _1156_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7602_ _1477_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4814_ _4179_ _4394_ _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8582_ _3701_ _0575_ _2557_ _3732_ _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5794_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7533_ _2650_ _2652_ _2728_ _2709_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _4317_ _4274_ _4160_ _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7464_ _1559_ _2387_ _2354_ _2661_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4676_ _4177_ _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8160__A1 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8160__B2 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9203_ _0152_ clknet_leaf_14_wb_clk_i as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6415_ _1411_ _1672_ _1678_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7395_ _2593_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput18 net18 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9134_ _0083_ clknet_leaf_61_wb_clk_i as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput29 net29 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6346_ _1573_ _1547_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9065_ _0014_ clknet_leaf_48_wb_clk_i as2650.stack\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6277_ _1548_ _1557_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8016_ _2340_ _4302_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5228_ _0440_ _0348_ _0564_ _4416_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4594__I _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8215__A2 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5159_ _0495_ as2650.stack\[5\]\[10\] as2650.stack\[4\]\[10\] _0496_ _0497_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7974__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8918_ _3047_ _1687_ _3987_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8849_ _2105_ _3904_ _3934_ _3912_ _3935_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7726__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8015__B _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8151__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8151__B2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4769__I _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6984__I _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9314__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6768__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4779__A1 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8390__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6940__A2 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ _4110_ _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8142__A1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7055__I _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8693__A2 _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6200_ _1458_ _1387_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7180_ _1564_ _2382_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__A2 _4485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _4158_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8996__A3 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6223__A4 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6964_ _2175_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5431__A2 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8703_ _3832_ _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1163_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7708__A1 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6895_ _2107_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6134__I _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8634_ _3680_ _3780_ _3781_ _3752_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5846_ _1141_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8381__A1 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5777_ _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8565_ _3682_ _3704_ _3716_ _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_124_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6931__A2 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7516_ _2185_ _2394_ _2712_ _2134_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4942__A1 _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4728_ _4135_ _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8496_ _4335_ _3648_ _3649_ _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4589__I _4169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7447_ _2307_ _2642_ _2645_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4659_ as2650.cycle\[6\] _4239_ _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8684__A2 _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7378_ _2475_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9117_ _0066_ clknet_leaf_11_wb_clk_i as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6329_ _1454_ _1612_ _1521_ _1579_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_89_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8436__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6447__A1 _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9048_ _3015_ _4096_ as2650.psu\[3\] _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6998__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8524__I _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6044__I _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7175__A2 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8372__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6979__I _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6922__A2 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8124__A1 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8427__A2 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6438__A1 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9023__C _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5661__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7938__A1 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_29_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_29_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8060__B1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7478__C _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5413__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ _1024_ _0987_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ _1910_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5177__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ _4421_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5793__I _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8350_ _0986_ _3509_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4924__A1 _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5562_ _0667_ _0815_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_129_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8115__A1 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7301_ _0556_ _1271_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8281_ _2210_ _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5493_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7232_ _2403_ _2434_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7941__C _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7163_ _2366_ _2131_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6114_ _4132_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8969__A3 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7094_ _4183_ _2296_ _2297_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _1185_ _1319_ _1332_ _1218_ _1179_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_86_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6129__I _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4872__I _4452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7996_ _3159_ _3164_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _2161_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8354__A1 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _2072_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8617_ _3114_ _2293_ _3765_ _2772_ _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ as2650.r123_2\[3\]\[3\] _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__A1 as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8548_ _3003_ _3683_ _3700_ _3552_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_124_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8012__C _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8657__A2 _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8479_ _3287_ _3619_ _3622_ _3632_ _3633_ _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_120_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7617__B1 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5891__A2 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7093__A1 _4512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8042__B1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8345__A1 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5159__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5159__B2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8896__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5118__I _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5331__A1 _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5882__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_opt_5_0_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8820__A2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7489__B _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7850_ _1634_ _2259_ _2288_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8584__A1 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _0859_ _1007_ _2014_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7781_ _2327_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _4406_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6732_ _1935_ _1947_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7139__A2 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6663_ as2650.stack\[3\]\[3\] _1892_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8402_ _3559_ _3322_ _2217_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ _4132_ _4151_ _4158_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__9182__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9382_ net48 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6594_ _1855_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6362__A3 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8333_ _2528_ _3493_ _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5545_ _0873_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5570__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__I _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7671__C _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8264_ _3038_ _3416_ _3426_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5476_ _0620_ _0808_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_132_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7311__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5472__B _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7215_ _2417_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5322__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8195_ _0932_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7862__A3 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7146_ _2131_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5873__A2 _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7075__A1 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8272__B1 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8275__S _4468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7077_ _1384_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6822__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6028_ _1301_ _1286_ _1316_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5698__I as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7090__A4 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7979_ net4 _3004_ _1457_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8327__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout53 net31 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6889__A1 as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6105__A3 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4777__I as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7153__I _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5864__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7066__A1 _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8263__B1 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9055__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8566__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6577__B1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_80 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_91 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7756__C _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6232__I _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7772__B _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ _4422_ _4203_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _0543_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7000_ _2206_ _1485_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4658__A3 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9046__A2 _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5192_ _0524_ _0527_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7998__I _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_44_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7057__A1 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5607__A2 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8951_ _1683_ _4017_ _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7012__B _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7902_ _3077_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8882_ _3957_ _3961_ _3963_ _3953_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_64_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8557__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4830__A3 _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7947__B _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7833_ _2998_ _3016_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7764_ _2952_ _2953_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8309__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4976_ _4305_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8309__B2 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6715_ _1941_ _1945_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7695_ _2829_ _2865_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7238__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6142__I _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6646_ _1886_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7532__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8778__B _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _0544_ _1752_ _1780_ as2650.r0\[2\] _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5981__I _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8316_ _3255_ _3449_ _3166_ _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ _0860_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9296_ _0245_ clknet_leaf_2_wb_clk_i as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7296__A1 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6099__A2 _4404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8247_ _3218_ _3382_ _3410_ _3210_ _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5459_ _0745_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_59_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4649__A3 _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_opt_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8178_ _3342_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9078__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7048__A1 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8245__B1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7129_ _2129_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7599__A2 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8796__A1 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8548__A1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__B1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7148__I _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5534__A1 _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7287__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9028__A2 _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6227__I _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6262__A2 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8539__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_opt_2_0_wb_clk_i clknet_3_3__leaf_wb_clk_i clknet_opt_2_0_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7211__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4970__I _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8442__I _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4830_ _4372_ _4172_ _4410_ _4411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5222__B1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7762__A2 _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4761_ _4309_ _4292_ _4342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6500_ _1748_ _1759_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7480_ _2677_ _2673_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ as2650.idx_ctrl\[1\] as2650.idx_ctrl\[0\] _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7514__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8598__B _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6431_ _1700_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9150_ _0099_ clknet_leaf_59_wb_clk_i as2650.r123\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6362_ _1045_ _1047_ _1117_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_66_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7278__A1 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8101_ _2168_ _2197_ _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5313_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__9220__CLK clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6293_ _1394_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9081_ _0030_ clknet_leaf_45_wb_clk_i as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8032_ _0918_ as2650.stack\[3\]\[0\] as2650.stack\[2\]\[0\] _3200_ _4488_ _3201_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5244_ _4350_ _0580_ _4289_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9019__A2 _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _4283_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8778__A1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8934_ _4312_ _2207_ _4000_ _2194_ _4001_ _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_65_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8865_ _3939_ _3948_ _3949_ _3752_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5976__I as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8352__I _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7816_ _4322_ _2997_ _3002_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8796_ _0374_ _3894_ _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8950__A1 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7747_ _1574_ _2936_ _2203_ _2239_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5764__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4959_ _0289_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7678_ _2857_ _2526_ _2527_ _2173_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5516__A1 _4499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ as2650.stack\[0\]\[13\] _1869_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__C1 _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7269__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5216__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9279_ _0228_ clknet_leaf_43_wb_clk_i as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8955__C _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5819__A2 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8769__A1 _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7441__A1 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__I as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6244__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7992__A2 _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6547__A3 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8941__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__B1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8865__C _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9042__B as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5570__B _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A2 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7341__I _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7432__A1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6980_ _2187_ _2174_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7983__A2 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5931_ _1190_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8650_ _0898_ _2797_ _3783_ _3786_ _3796_ _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ _4113_ _4172_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_94_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8932__A1 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7735__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7601_ _1691_ _2792_ _2794_ _2795_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5746__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4813_ _4389_ _4393_ _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8581_ _2648_ _0580_ _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5793_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7532_ _1599_ _0893_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7944__C _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4744_ _4308_ _4321_ _4324_ _4325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7499__A1 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7463_ _2389_ _2660_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4675_ _4255_ _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__I _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9202_ _0151_ clknet_leaf_14_wb_clk_i as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6414_ _1686_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7394_ as2650.pc\[5\] _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9133_ _0082_ clknet_leaf_61_wb_clk_i as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6345_ _1574_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8999__A1 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6276_ _1558_ _1410_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_9064_ _0013_ clknet_leaf_42_wb_clk_i as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8015_ _3170_ _3175_ _3181_ _3183_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5227_ _0365_ _0563_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _0387_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7423__A1 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5089_ _0290_ _0292_ _0307_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7974__A2 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8917_ _2171_ _1687_ _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__A2 _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8848_ as2650.r123\[2\]\[7\] _3928_ _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8923__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7726__A2 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9266__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8779_ _1450_ _4179_ _4269_ _4446_ _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4960__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6162__A1 _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4785__I _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7161__I _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7414__A1 _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7965__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6768__A3 _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__A2 _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8390__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8720__I _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4951__A2 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8142__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6240__I _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6153__A1 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6130_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7653__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6456__A2 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ _1334_ _1286_ _1335_ _1347_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8167__I as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8850__B1 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9203__D _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9139__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5012_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6963_ _2171_ _2173_ _2174_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5967__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8116__B _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9289__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8702_ _3832_ _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6894_ _1898_ _2108_ _2113_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7708__A2 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8633_ _1102_ _3680_ _3781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5719__A1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5845_ _0977_ _1143_ _1145_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8381__A2 _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8564_ _3690_ _2373_ _2533_ _0463_ _3715_ _3716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5776_ as2650.pc\[5\] _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7515_ _4428_ _2711_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4727_ _4160_ _4306_ _4307_ _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8495_ _4478_ _2956_ _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4942__A2 _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6150__I _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7446_ _2600_ _2643_ _2644_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4658_ _4121_ as2650.cycle\[4\] _4238_ _4120_ _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_107_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7690__B _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7377_ _2413_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4589_ _4169_ _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9116_ _0065_ clknet_leaf_7_wb_clk_i as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6328_ _1603_ _1606_ _1611_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6447__A2 _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8841__B1 _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9047_ _4100_ _4104_ _1428_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6259_ _1543_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5958__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6325__I _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5186__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8124__A2 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6135__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6995__I _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7883__A1 _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6686__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7635__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6438__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7938__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8060__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5949__A1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6610__A2 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6235__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4621__A1 _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_69_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_69_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5630_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5177__A2 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6374__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5561_ _0893_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4924__A2 _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8115__A2 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7300_ _2443_ _2499_ _2500_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6126__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5492_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8280_ _3437_ _3439_ _3441_ _3442_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7231_ _2305_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7874__A1 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6677__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7162_ _2122_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6113_ _0697_ _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7093_ _4512_ _1356_ _1357_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_99_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5314__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7669__C _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8051__A1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7995_ _3160_ _3161_ _3163_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6145__I _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _2160_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _2093_ _2101_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8354__A2 _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8616_ _2179_ _1546_ _3757_ _3764_ _3062_ _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5828_ _1134_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8547_ _1200_ _3684_ _3687_ _3699_ _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5759_ _1034_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6117__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9304__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8478_ _0854_ _3444_ _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6668__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7429_ _2622_ _2626_ _2357_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7617__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7617__B2 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8290__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7093__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8535__I _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8042__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8042__B2 _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5894__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8345__A2 _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6356__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A2 _4483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6939__B _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5331__A2 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__A1 _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9050__B _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6800_ _0782_ _1024_ _1981_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7780_ _2327_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5398__A2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4992_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6731_ _1798_ _1929_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8336__A2 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6662_ _1086_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9327__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8401_ _2172_ _2778_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9381_ net47 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _1046_ _1854_ _1051_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8332_ _3491_ _3461_ _3492_ _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_118_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5544_ _0799_ _0797_ _0808_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7847__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8263_ _3010_ _3423_ _3425_ _3231_ _3183_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5475_ _0725_ _0802_ _0807_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_117_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7214_ _0930_ _4195_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8194_ _0902_ _2582_ _3358_ _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7145_ _2330_ _2347_ _2348_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5873__A3 _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8272__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7075__A2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8272__B2 _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7076_ _1450_ _2242_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6822__A2 _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6027_ _1219_ _1312_ _1315_ _1220_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_86_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8575__A2 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5389__A2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7978_ _1457_ _3145_ _3146_ _3147_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6929_ _1372_ _2140_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout54 net28 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6338__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8023__C _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6889__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5219__I _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6105__A4 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6510__A1 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8974__B _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8263__A1 _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7066__A2 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8263__B2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4793__I _4373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8015__A1 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_70 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6577__B2 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_81 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_61_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_92 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8318__A2 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A1 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5552__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5260_ _0591_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_142_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5191_ _0524_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8254__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7057__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5068__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8950_ _2999_ _1412_ _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8006__A1 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7901_ _2193_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7012__C _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8881_ net45 _3962_ _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8557__A2 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7832_ _3014_ _3004_ _3015_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7763_ _4237_ _2145_ _2144_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8124__B _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4975_ _4349_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6714_ _1943_ _1944_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6423__I _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7694_ as2650.pc\[12\] _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5791__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7963__B _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6645_ as2650.r123\[3\]\[6\] _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6576_ as2650.r0\[4\] _1014_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8315_ _3343_ _3476_ _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4878__I _4458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5527_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9295_ _0244_ clknet_leaf_69_wb_clk_i as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7296__A2 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8246_ _3405_ _3406_ _3408_ _3409_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5458_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8177_ _2587_ _2381_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5389_ _0626_ _0722_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7128_ _2331_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7048__A2 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8245__B2 as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8796__A2 _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7059_ _1033_ _2262_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A1 as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5231__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5782__A2 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6731__A1 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5534__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7287__A2 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6936__C _4421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8236__A1 _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8236__B2 _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9172__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5470__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7211__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7339__I as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5222__A1 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7762__A3 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5222__B2 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _4340_ _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _4271_ _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8172__B1 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8711__A2 _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6430_ as2650.r0\[0\] _0960_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6722__A1 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6361_ _1483_ _1642_ _1643_ _1644_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_143_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8100_ _3224_ _3260_ _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5312_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7278__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8475__A1 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9080_ _0029_ clknet_leaf_46_wb_clk_i as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6292_ _1361_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5289__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8031_ _3199_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5243_ _0481_ _0557_ _0572_ _0483_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__8227__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5174_ as2650.r123\[0\]\[3\] _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8778__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8933_ _2136_ _1403_ _1371_ _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A1 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8864_ net42 _3945_ _3949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7738__B1 _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7815_ _2998_ _3001_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8795_ as2650.r123\[1\]\[1\] _3889_ _3891_ _1711_ _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5213__A1 _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8950__A2 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7746_ _2935_ _2936_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4958_ _0291_ _0292_ _0296_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7677_ _2864_ _2869_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4889_ as2650.psu\[1\] _4470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6628_ _1021_ _1871_ _1877_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6713__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__B1 _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6559_ as2650.r123_2\[1\]\[6\] _1726_ _1822_ _1723_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4724__C2 _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7269__A2 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8466__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9278_ _0227_ clknet_leaf_43_wb_clk_i as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8229_ _1581_ _2611_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8769__A2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7441__A2 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6244__A3 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7992__A3 _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7729__B1 _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5204__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6063__I _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__I _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8457__A1 _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__B2 _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7622__I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8209__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5691__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6238__I _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7432__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5443__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5443__B2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ _1190_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5861_ _1154_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7069__I _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7600_ _1420_ _2329_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8932__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4812_ _4390_ _4392_ _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8580_ _0681_ _1446_ _2533_ _0560_ _3677_ _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5792_ as2650.pc\[7\] _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7531_ _2383_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4743_ _4322_ _4323_ _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8402__B _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7499__A2 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7462_ _2656_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8696__A1 _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4674_ _4252_ _4254_ _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9201_ _0150_ clknet_leaf_22_wb_clk_i net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6413_ _0963_ _1473_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7393_ _2307_ _2591_ _2592_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9132_ _0081_ clknet_leaf_55_wb_clk_i as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8448__A1 as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6344_ _1575_ _0905_ _1518_ _1627_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9063_ _0012_ clknet_leaf_48_wb_clk_i as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6275_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8014_ _3182_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5226_ _0363_ _0553_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7671__A2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5682__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5157_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7423__A2 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8620__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5088_ _0421_ _0424_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5434__A1 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4891__I _4471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8916_ _3981_ _1115_ _3986_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7187__A1 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8847_ _3927_ _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8384__B1 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8923__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8778_ _1229_ _1378_ _1375_ _4116_ _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6934__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7729_ _1486_ _2125_ _2917_ _2919_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8687__A1 _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__A2 _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8439__A1 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6767__B _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6465__A3 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8982__B _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5673__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7414__A2 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5425__A1 _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7178__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9210__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8914__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6925__A1 _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6776__I1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8142__A3 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7350__A1 _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4976__I _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7653__A2 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8850__A1 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _4171_ _1177_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8850__B2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5011_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6962_ _2158_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8116__C _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8701_ _3831_ _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5913_ _1206_ _0931_ _4201_ _1172_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6893_ as2650.stack\[4\]\[3\] _2109_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8366__B1 _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8905__A2 _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8632_ _0829_ _1677_ _3771_ _3779_ _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5844_ as2650.stack\[1\]\[8\] _1144_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6916__A1 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5719__A2 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8563_ _1683_ _3688_ _3712_ _3714_ _2411_ _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5775_ _1089_ _1093_ _1095_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7527__I _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7514_ _1599_ _0893_ _2710_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4726_ as2650.holding_reg\[0\] _4160_ _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8494_ _2273_ _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7445_ _1424_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4657_ as2650.cycle\[3\] _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5047__I _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7376_ _2566_ _2472_ _2346_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4588_ _4152_ _4168_ _4169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9115_ _0064_ clknet_leaf_7_wb_clk_i as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4886__I _4466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6327_ _1607_ _0555_ _0675_ _4403_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9046_ _3019_ _4103_ _4104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6258_ _1336_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6447__A3 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8841__A1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _0545_ _4175_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _4114_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9233__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6080__A1 _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4630__A2 as2650.alu_op\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7580__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8977__B _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6135__A2 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7635__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6438__A3 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7399__A1 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7938__A3 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5420__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8060__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6071__A1 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4621__A2 _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6374__A2 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7571__A1 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _0825_ _0567_ _0886_ _0324_ _0892_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5295__C _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_38_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5491_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6126__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7230_ _2380_ _2384_ _2432_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9106__CLK clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7874__A2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5885__A1 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7161_ _2364_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8178__I _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6112_ _1397_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7626__A2 as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7092_ _2293_ _0829_ _0898_ _2295_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_99_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9256__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _1329_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7810__I _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8051__A2 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7994_ _2280_ _2285_ _2954_ _3162_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6945_ as2650.addr_buff\[0\] _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9000__A1 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6876_ _1703_ _2100_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5827_ as2650.r123_2\[3\]\[2\] _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8615_ _3689_ _3763_ _1546_ _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5758_ _1053_ _1079_ _1080_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5573__B1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8546_ _0361_ _1677_ _3678_ _3698_ _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ _4289_ _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7314__A1 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8477_ _3034_ _3629_ _3631_ _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6117__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5689_ as2650.pc\[12\] _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7428_ _2622_ _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8088__I _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7359_ _2492_ _0555_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7617__A2 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8814__B2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9029_ _4080_ _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8290__A2 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6336__I _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8042__A2 _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A1 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7876__B _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6356__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9129__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9382__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7305__A1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8500__B _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9279__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6020__B _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5095__A2 _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4991_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _0782_ _1007_ _1930_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6661_ _1896_ _1891_ _1897_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7077__I _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8400_ _2855_ _2879_ _2604_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5612_ _0943_ _0926_ _4123_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_9380_ net46 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6592_ _4495_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8331_ _0900_ _4363_ _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5543_ _0873_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8262_ _2647_ _3424_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5474_ _0725_ _0807_ _0802_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7847__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5858__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7213_ _2412_ _1664_ _2415_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_105_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9049__A1 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8193_ _2541_ _1543_ _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5325__I _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7144_ _2313_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5873__A4 _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8272__A2 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7075_ _2126_ _2132_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5086__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6283__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6026_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7783__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5995__I as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7977_ _0861_ _1467_ _3097_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4597__A1 _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6928_ _1442_ _2142_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7535__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6859_ _2083_ _2084_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6338__A2 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9119__D _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8529_ _3677_ _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5849__A1 as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7450__I _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_60 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_71 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8281__I _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_82 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_93 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7526__A1 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6329__A2 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5145__I _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5190_ _0420_ _0424_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4984__I _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8254__A2 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8006__A2 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7900_ _0404_ _3032_ _3076_ _1031_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8880_ _3938_ _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__A1 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7831_ _2171_ _2226_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4974_ _0297_ _0305_ _0312_ _0284_ _4298_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_7762_ _2146_ _2950_ _2951_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_53_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_53_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6713_ as2650.r0\[7\] _0981_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7693_ _2379_ _2884_ _2885_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7517__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6644_ _1885_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6575_ _1833_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8314_ _3466_ _3467_ _3475_ _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5526_ _4359_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4751__A1 _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9294_ _0243_ clknet_leaf_69_wb_clk_i as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8245_ as2650.stack\[6\]\[5\] _3199_ _0380_ as2650.stack\[7\]\[5\] _4497_ _3409_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5457_ _0746_ _0748_ _0750_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7296__A3 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8176_ _3214_ _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5388_ _0628_ _0615_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7127_ _4426_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4894__I _4471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7048__A3 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7270__I _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7058_ _4222_ _2259_ _2260_ _2261_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_86_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6009_ _0709_ _1157_ _1182_ _1298_ _0700_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_39_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7756__A1 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5231__A2 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7508__A1 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7445__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8236__A2 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6247__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7995__A1 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7747__A1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5222__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4690_ _4250_ _4270_ _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8172__B2 _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4733__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6360_ _1427_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ _4301_ _0645_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8475__A2 _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6291_ _1396_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8030_ _0376_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5289__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5242_ _0578_ _0570_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8227__A2 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5173_ _0403_ _4287_ _0510_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__I _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8778__A3 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7986__A1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8932_ _4234_ _1455_ _1370_ _1408_ _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_84_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A2 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8863_ _1065_ _3941_ _3947_ _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7738__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7738__B2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7814_ _2120_ _1638_ _3000_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8794_ _3892_ _3895_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__A2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7745_ net50 _2615_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4957_ _0291_ _0292_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7676_ _2617_ _2868_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8163__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ _4468_ _4469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8163__B2 _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4889__I as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6627_ as2650.stack\[0\]\[12\] _1873_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7265__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6713__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4724__A1 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _1821_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4724__B2 _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ _0323_ _0838_ _0842_ _4349_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8466__A2 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6489_ _4299_ _1016_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9277_ _0226_ clknet_leaf_54_wb_clk_i as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6477__A1 as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8228_ _2595_ _3391_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8096__I _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8159_ _2971_ _3318_ _3324_ _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7977__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5452__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7729__A1 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5204__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7884__B _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A2 _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A1 _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8457__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7903__I _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5423__I _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5691__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6254__I _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5860_ _0332_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _4143_ _4391_ _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8932__A3 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _1089_ _1108_ _1109_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7530_ _2377_ _2725_ _2726_ _2437_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4742_ _4129_ _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8145__A1 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7461_ _2633_ _2657_ _2658_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4673_ _4122_ _4253_ _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8696__A2 _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9200_ _0149_ clknet_3_6__leaf_wb_clk_i net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6412_ _1682_ _1668_ _1685_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7392_ _2566_ _2377_ _1425_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9131_ _0080_ clknet_leaf_55_wb_clk_i as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6343_ _1576_ _1626_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8448__A2 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9062_ _0011_ clknet_leaf_52_wb_clk_i as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6274_ _1525_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5131__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8013_ _0948_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5225_ _0556_ _0457_ _0561_ _4374_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7969__B _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5087_ _0421_ _0424_ _4333_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8915_ as2650.stack\[2\]\[7\] _3982_ _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8846_ _3932_ _3933_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8384__A1 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7187__A2 _4458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8384__B2 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5198__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8777_ _3829_ _3871_ _3879_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _0575_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7728_ _2918_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7659_ net52 _2306_ _2852_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8687__A2 _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9162__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6162__A3 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5952__B _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8439__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9329_ _0278_ clknet_leaf_9_wb_clk_i as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5370__A1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A1 _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__A4 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5673__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8611__A2 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6622__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5425__A2 _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8375__A1 _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7178__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5189__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6925__A2 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4787__I1 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5418__I _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7350__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4795__S0 _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8850__A2 _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__I _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ net7 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4992__I _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6613__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5416__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6961_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8700_ _0917_ _1047_ _1117_ _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5912_ _4216_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8366__A1 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _1896_ _2108_ _2112_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8366__B2 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8631_ _1539_ _3684_ _3777_ _3778_ _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5843_ _1142_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6916__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9185__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8562_ _3713_ _0681_ _1515_ _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5774_ as2650.stack\[1\]\[4\] _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7513_ _2650_ _2652_ _2709_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8669__A2 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4725_ _4305_ _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5328__I _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8493_ _3646_ _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7444_ _2305_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4656_ _4236_ _4119_ _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7375_ _2573_ _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4587_ _4158_ _4167_ _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9114_ _0063_ clknet_leaf_49_wb_clk_i as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6326_ _1608_ _0933_ _1609_ as2650.overflow _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9045_ _3058_ _1413_ _4102_ _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6257_ _1515_ _1537_ _1541_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6447__A4 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8841__A2 _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5208_ _0544_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ _1384_ _4237_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5998__I _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5139_ _4431_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_8_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8357__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4630__A3 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8829_ _1989_ _3919_ _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8109__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A1 _4512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__I _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8549__I _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6540__B1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8993__B _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7096__A1 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8832__A2 _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7399__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8596__A1 _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6071__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8233__B _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8899__A2 _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5490_ _4360_ _4364_ _4369_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_129_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7323__A2 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8520__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7160_ _4240_ _2282_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5885__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _1396_ _4213_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7087__A1 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _0673_ _2294_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _0814_ _1171_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9230__D _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8587__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7993_ _4115_ _2302_ _2926_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6944_ _2158_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8339__A1 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9000__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8143__B _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6875_ _2096_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7011__A1 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8614_ _1517_ _3761_ _3762_ _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5826_ _1133_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7982__B _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8545_ _1680_ _3688_ _3697_ _2411_ _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5757_ as2650.stack\[1\]\[2\] _1063_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5573__B2 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4708_ _4266_ _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8476_ _3274_ _3619_ _3630_ _2960_ _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7314__A2 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5688_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8511__A1 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4897__I _4468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7427_ _2550_ _2624_ _2551_ _2625_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_68_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7273__I _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4639_ _4216_ _4219_ _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7358_ _2539_ _0674_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9200__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6309_ _0455_ _0347_ _0451_ _1554_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7289_ _2379_ _2489_ _2490_ _2437_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9028_ _3005_ _4080_ _1492_ _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8578__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7250__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7448__I _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__I _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7553__A2 _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7305__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8502__A1 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_2__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7183__I _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4600__I _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5095__A3 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ _4379_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6660_ as2650.stack\[3\]\[2\] _1892_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8741__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5611_ _4192_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5555__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ _1346_ _1696_ _1853_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8330_ _0900_ _4363_ _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5542_ _0800_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8261_ _2594_ _2539_ _3308_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__9223__CLK clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__I _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7212_ _2403_ _2341_ _2413_ _0353_ _2414_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5858__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8192_ _2314_ _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9049__A2 _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7143_ _2332_ _2336_ _2343_ _2346_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7821__I _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7074_ _2258_ _2263_ _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7480__A1 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6025_ _0784_ _4510_ _1185_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5341__I _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7977__B _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7232__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7976_ net4 _1404_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5243__B1 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7783__A2 _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8980__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6927_ _0928_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4597__A2 _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6858_ _0859_ _2036_ _2061_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__7535__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6338__A3 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5809_ as2650.stack\[0\]\[2\] _1121_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6789_ _2001_ _2017_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8601__B _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8528_ _3638_ _3681_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7299__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8459_ _3095_ _3613_ _3614_ _3528_ _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5849__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6347__I _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__I _4475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_61 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8971__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_72 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_83 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_94 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9246__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__B _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7214__A1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7830_ _0543_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8962__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7765__A2 _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7761_ _2145_ _1385_ _2140_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ _0306_ _0291_ _0310_ _0311_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_6712_ _1839_ _1942_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7692_ _2857_ _2306_ _2852_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7517__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8714__A1 _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6643_ as2650.r123\[3\]\[5\] _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6725__B1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8190__A2 _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6574_ _1834_ _1836_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8313_ _3218_ _3449_ _3474_ _3369_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_22_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_22_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5525_ as2650.r123\[0\]\[7\] _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9293_ _0242_ clknet_leaf_8_wb_clk_i as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4751__A2 _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8244_ _3195_ _3407_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5456_ _0712_ _0751_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7296__A4 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8175_ _1084_ _3167_ _3340_ _3254_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5700__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5387_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7828__I0 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7126_ _2319_ _2322_ _2326_ _2329_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6256__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5071__I _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7057_ _4257_ _0334_ _1349_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9119__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6008_ _1184_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7205__A1 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8953__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7959_ _3105_ _3130_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9269__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5231__A3 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7508__A2 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8705__A1 _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5519__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6192__A1 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7692__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6247__A2 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7747__A2 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8944__A1 _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8172__A2 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5156__I _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8895__C _3970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5310_ _4375_ as2650.r123_2\[0\]\[5\] _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _1514_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7683__A1 _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5241_ _4456_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _4288_ _0488_ _0509_ _0401_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7435__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8931_ _3997_ _3998_ _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5997__A1 _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8862_ _0441_ _3942_ _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8935__A1 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7738__A2 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7813_ _4353_ _2999_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5749__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8793_ _4463_ _3894_ _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6410__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7744_ _2934_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4956_ _0294_ _4293_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7675_ _2865_ _2867_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ as2650.psu\[0\] _4468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6626_ _1012_ _1870_ _1876_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6557_ _1817_ _1820_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4724__A2 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5921__A1 _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ _4430_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9276_ _0225_ clknet_leaf_54_wb_clk_i as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8466__A3 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6488_ _0442_ _0981_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8227_ _2540_ _3308_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _0736_ _0773_ _0321_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8158_ _2841_ _3306_ _3323_ _3088_ _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7426__A1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7109_ _2312_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8623__B1 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8089_ _1066_ _1056_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7977__A2 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4660__A1 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7729__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8926__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6360__I _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8996__B _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4715__A2 _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7417__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7417__B2 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5979__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8917__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8750__I _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4810_ _4208_ _4153_ _4198_ _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ as2650.stack\[1\]\[6\] _1094_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8932__A4 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6943__A3 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ as2650.holding_reg\[0\] _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7366__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6270__I _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7460_ _0756_ _0770_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6156__A1 _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4672_ _4188_ _4120_ _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6411_ _1683_ _1684_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7391_ _2541_ _2493_ _2590_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9130_ _0079_ clknet_leaf_56_wb_clk_i as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6342_ _1577_ _1623_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4939__B _4519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7656__A1 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9061_ _0010_ clknet_leaf_50_wb_clk_i as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ _0677_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8012_ _4183_ _3178_ _3180_ _1351_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5224_ _4396_ _0560_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7408__A1 _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5155_ _0378_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5550__S _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5086_ _0299_ _0303_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7050__B _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8914_ _3981_ _1108_ _3985_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8845_ _2100_ _3891_ _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8384__A2 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8776_ as2650.stack\[7\]\[14\] _3869_ _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6395__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7592__B1 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _1243_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6934__A3 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7727_ _2320_ _2367_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4939_ _4288_ _4463_ _4519_ _4286_ _4520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6180__I _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7658_ _1424_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7895__A1 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6609_ _1100_ _1862_ _1865_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7589_ _2165_ _2778_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_opt_1_0_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9328_ _0277_ clknet_leaf_6_wb_clk_i as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8844__B1 _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9259_ _0208_ clknet_leaf_37_wb_clk_i as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A2 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6355__I _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6622__A2 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5425__A3 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4633__A1 _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6386__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8503__C _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7186__I _4446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__I2 as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6090__I _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4603__I _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5361__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4795__S1 _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7789__C _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6265__I _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6960_ as2650.addr_buff\[3\] _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _1204_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6891_ as2650.stack\[4\]\[2\] _2109_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8366__A2 _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8630_ _1560_ _1548_ _2438_ _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5842_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6377__A1 as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6916__A3 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8561_ _1396_ _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5773_ _1052_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7512_ _1597_ _0841_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4724_ _4299_ _4175_ _4300_ _4302_ _4303_ _4304_ _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_8492_ _4152_ _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7443_ _2595_ _2493_ _2641_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7877__A1 _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4655_ as2650.cycle\[1\] _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7824__I _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7374_ _2417_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4586_ _4163_ _4166_ _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7629__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9113_ _0062_ clknet_leaf_50_wb_clk_i as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6325_ _0454_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_107_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9044_ _3097_ _4101_ _4076_ _4095_ _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_88_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6256_ _1538_ _0905_ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5207_ as2650.r0\[4\] _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6187_ _1445_ _1471_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8054__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5138_ _0475_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7801__A1 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6175__I _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5069_ _4190_ _0406_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5663__I0 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8828_ _0374_ _3915_ _3917_ as2650.r123\[2\]\[1\] _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8759_ _1045_ _3812_ _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8109__A2 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A2 _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7868__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6540__B2 _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8293__A1 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7096__A2 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6085__I _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4606__A1 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__A3 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8348__A2 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7909__I _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6359__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8233__C _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6034__B _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5031__A1 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5582__A2 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7859__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7644__I _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8520__A2 _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5164__I _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6110_ _4219_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8284__A1 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7087__A2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7090_ _4399_ _0361_ _0463_ _0560_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_112_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _1327_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8587__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7992_ _2143_ _2950_ _2972_ _2266_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__9152__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6943_ _2133_ _2139_ _2149_ _2157_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__8339__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6874_ _2088_ _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7011__A2 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8613_ _1360_ _0638_ _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5825_ as2650.r123_2\[3\]\[1\] _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5339__I _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7982__C _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8544_ _3689_ _3690_ _3696_ _1514_ _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5756_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _4283_ _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8475_ _2841_ _3421_ _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5687_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8511__A2 _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7426_ _2623_ _0685_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4638_ _4209_ _4135_ _4217_ _4218_ _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7357_ _1487_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4569_ _4149_ _4150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6308_ as2650.psu\[7\] _1581_ _1587_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7288_ _2467_ _2434_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5089__A1 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9027_ _4085_ _4086_ _4087_ _3118_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _1523_ _0969_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4836__A1 _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8578__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7250__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5564__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8502__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6513__A1 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8266__A1 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5712__I _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9175__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8018__A1 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5610_ _0934_ _0937_ _0940_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6590_ as2650.r123_2\[1\]\[7\] _1726_ _1852_ _1702_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5555__A2 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ _0798_ _0803_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7374__I _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8260_ _2961_ _3415_ _3418_ _3419_ _3422_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5472_ _0718_ _0719_ _0729_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7211_ _0408_ _2404_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8191_ _3351_ _3354_ _3355_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7142_ _2345_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8257__A1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6807__A2 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7073_ _2224_ _2149_ _2276_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9241__D _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6024_ _4509_ _0781_ _1157_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7480__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7232__A2 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7975_ as2650.psu\[7\] _1691_ _3144_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7549__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5243__B2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6926_ _2140_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6857_ _0822_ _2082_ _1040_ _0859_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xfanout46 net48 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8732__A2 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5808_ _1071_ _1120_ _1123_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6743__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6788_ _2012_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8527_ _3644_ _3657_ _3679_ _3680_ _1054_ _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5739_ as2650.stack\[1\]\[0\] _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8458_ _3212_ _3601_ _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8496__A1 _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7409_ _1091_ net10 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8389_ _3532_ _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8799__A2 _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5482__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6363__I _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_62 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8971__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7774__A3 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_73 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_84 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_95 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_72_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7797__C _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8411__A1 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7214__A2 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6273__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8962__A2 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7760_ _2281_ _2148_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4972_ _4296_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _0743_ _0993_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7691_ _2856_ _2727_ _2883_ _2724_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8714__A2 _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6642_ _1884_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6725__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6573_ as2650.r0\[0\] _1835_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8312_ _3469_ _3470_ _3472_ _3473_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_5524_ _0788_ _0603_ _0857_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8478__A1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9292_ _0241_ clknet_leaf_69_wb_clk_i as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8243_ _3245_ as2650.stack\[5\]\[5\] as2650.stack\[4\]\[5\] _0385_ _3407_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ as2650.holding_reg\[6\] _4162_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_62_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8174_ _3168_ _3306_ _3339_ _3214_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5386_ _0714_ _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7125_ _2328_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7828__I1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7453__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8650__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7056_ _4251_ _2224_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6256__A3 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8663__I _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ _0634_ _1262_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_74_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7205__A2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8953__A2 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6183__I _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7958_ _4121_ _3119_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _2122_ _2123_ _4252_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5231__A4 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7889_ _3065_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7508__A3 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8705__A2 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5519__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7228__B _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6192__A2 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8469__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7141__A1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7692__A2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8059__B _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8641__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5455__A1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8573__I _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9213__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8944__A2 _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A2 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7132__A1 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _0566_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6268__I _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5171_ _0375_ _0505_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7435__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8632__A1 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7986__A3 _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8930_ _1607_ _1420_ _1398_ _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5997__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8416__C _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8861_ _3939_ _3944_ _3946_ _3752_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6217__B _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8935__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7812_ _1388_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8792_ _3893_ _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5749__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7743_ _2150_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4955_ _0293_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8699__A1 _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7674_ _2830_ _2834_ _2866_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4886_ _4466_ _4467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8151__C _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6625_ as2650.stack\[0\]\[11\] _1873_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7371__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6556_ _1766_ _1818_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5507_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9275_ _0224_ clknet_leaf_54_wb_clk_i as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6487_ as2650.r0\[2\] _1752_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8226_ _2476_ _3388_ _3389_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8871__A1 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5438_ _0314_ _0768_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5685__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8157_ _2596_ _3321_ _3322_ _1443_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5369_ as2650.stack\[6\]\[12\] _4473_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7108_ _2221_ _1188_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7426__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8623__A1 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8088_ _2245_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9236__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8393__I _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7039_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6906__I _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8326__C _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8926__A2 _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__A1 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__A3 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__I1 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4715__A3 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8568__I _4409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__A1 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8311__B1 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7665__A2 _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8862__A1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6468__A3 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7417__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8614__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8517__B _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8009__S _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5720__I _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8236__C _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8917__A2 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6928__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7647__I _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__A1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6943__A4 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _4259_ _4306_ _4318_ _4320_ _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4671_ _4192_ _4119_ _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7353__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6156__A2 _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6410_ _1672_ _1666_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9109__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7390_ _2571_ _2589_ _2374_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _0861_ _1624_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9060_ _0009_ clknet_leaf_52_wb_clk_i as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6272_ _1550_ _1551_ _1553_ _1556_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8011_ _1057_ _2296_ _3179_ _4183_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__9259__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6864__B1 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5223_ _0557_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7408__A2 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8605__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5154_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7331__B _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__I _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5085_ _0422_ _0316_ _4523_ _0298_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_84_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8913_ as2650.stack\[2\]\[6\] _3982_ _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4642__A2 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9030__A1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8844_ _0845_ _3927_ _3928_ as2650.r123\[2\]\[6\] _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7041__B1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7592__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8775_ _3827_ _3871_ _3878_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5987_ _0543_ _1234_ _1195_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6395__A2 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4938_ _4502_ _4518_ _4519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7726_ _1324_ _2381_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7657_ _2815_ _2727_ _2850_ _2536_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7344__A1 _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ _4397_ _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6608_ as2650.stack\[5\]\[5\] _1863_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7588_ _2779_ _2782_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7895__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6539_ _0743_ _1038_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9327_ _0276_ clknet_leaf_12_wb_clk_i as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8844__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9258_ _0207_ clknet_leaf_38_wb_clk_i as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5658__A1 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8209_ _3196_ _3373_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9189_ _0138_ clknet_leaf_19_wb_clk_i net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6083__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5425__A4 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4633__A2 _4117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__S _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9021__A1 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__A2 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__I3 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8835__A1 _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6310__A2 _4182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__A2 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9012__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ _4394_ _1158_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6890_ _1894_ _2108_ _2111_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5841_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7574__A1 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7377__I _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8560_ _3710_ _3711_ _1535_ _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7511_ _2698_ _2707_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4723_ as2650.r123\[1\]\[0\] as2650.r123\[0\]\[0\] as2650.r123_2\[1\]\[0\] as2650.r123_2\[0\]\[0\]
+ _4146_ _4301_ _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_8491_ _1187_ _3209_ _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7442_ _2309_ _2640_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4654_ as2650.cycle\[7\] _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7877__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5888__A1 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9081__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7373_ _2572_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4585_ _4165_ _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6324_ as2650.psl\[7\] _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9112_ _0061_ clknet_leaf_51_wb_clk_i as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8826__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9043_ _4515_ _1402_ _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6255_ _0827_ _0640_ _0665_ _1539_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5206_ _0519_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6186_ _1441_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8054__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5137_ _0470_ _0472_ _0473_ _0324_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7801__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5068_ _0405_ _4253_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5812__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5663__I1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9003__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8827_ _3918_ _3920_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6191__I _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8758_ _1908_ _3862_ _3867_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7709_ _2352_ _2897_ _2900_ _2758_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7317__B2 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8620__B _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8689_ as2650.stack\[5\]\[11\] _3819_ _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7868__A2 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5879__A1 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6140__B _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7096__A3 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7750__I _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8067__B _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4854__A2 as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4606__A2 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8348__A3 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9329__D _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6359__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5031__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7308__A1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7925__I _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7859__A2 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A1 _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5414__S0 _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8520__A3 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8284__A2 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A1 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _0821_ _1175_ _1171_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5180__I _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7795__A1 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7991_ _2255_ _2262_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6942_ _1664_ _1463_ _2151_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_16_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7547__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6873_ _2061_ _2097_ _2086_ _0909_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__9239__D _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8612_ _3724_ _1024_ _3759_ _0695_ _3760_ _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5824_ _1132_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7011__A3 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5755_ _0506_ _1035_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8543_ _3689_ _3695_ _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8440__B _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ _4286_ _4287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8474_ _3263_ _3624_ _3628_ _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5686_ as2650.r123\[0\]\[4\] as2650.r123_2\[0\]\[4\] _4108_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7425_ _2623_ _0685_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4637_ _4140_ _4142_ _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5355__I _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7356_ _2549_ _2555_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4568_ as2650.ins_reg\[1\] _4149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6307_ _1588_ _1554_ _0676_ _1589_ _1590_ _0455_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7287_ _1076_ _2384_ _2488_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6286__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5089__A2 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9026_ _4357_ _4085_ _4087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6238_ _4251_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4836__A2 _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6169_ _0691_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7786__A1 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8615__B _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7538__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7710__A1 _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6513__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8266__A2 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6277__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8018__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7226__B1 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8525__B _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5627__I1 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7529__A1 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6752__A2 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _0871_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4763__A1 _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ _4313_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7701__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7210_ _4427_ _2334_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8190_ _3351_ _3354_ _4256_ _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7141_ _2216_ _2344_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8486__I _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8257__A2 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5903__I _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7072_ _1476_ _2264_ _2268_ _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_87_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4818__A2 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6023_ _1228_ _1309_ _1310_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__5124__B _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7768__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7974_ _1691_ _1413_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__A1 _4503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5243__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6925_ _4210_ _1661_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6856_ _2036_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8193__A1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5807_ as2650.stack\[0\]\[1\] _1121_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8170__B _4498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7940__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6743__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6787_ _2014_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8526_ _3677_ _3680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5738_ _1052_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8457_ _3598_ _3101_ _3287_ _3601_ _3612_ _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8496__A2 _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ _0998_ _0987_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7408_ _2593_ _2606_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8388_ _3535_ _3545_ _3546_ _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7339_ as2650.pc\[4\] _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__I _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8329__C _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9009_ _1383_ _3011_ _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7471__A3 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5482__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A2 _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_63 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8971__A3 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7774__A4 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_74 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_85 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8184__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8080__B _4497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A1 _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6498__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9142__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7143__C _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9292__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__A1 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _0284_ _0298_ _0308_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8962__A3 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _1785_ _1939_ _1940_ _1842_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7690_ _1488_ _2870_ _2876_ _2882_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8175__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6641_ as2650.r123\[3\]\[4\] _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7922__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ as2650.r123\[0\]\[7\] as2650.r123_2\[0\]\[7\] _4108_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8311_ _0918_ as2650.stack\[3\]\[7\] as2650.stack\[2\]\[7\] _3200_ _3241_ _3473_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_5523_ _0512_ _0845_ _0856_ _4285_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9291_ _0240_ clknet_leaf_68_wb_clk_i as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8478__A2 _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6489__A1 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5454_ as2650.r123\[0\]\[6\] _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8242_ _1590_ as2650.stack\[3\]\[5\] as2650.stack\[2\]\[5\] _3199_ _4487_ _3406_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_69_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5161__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8173_ _3307_ _3338_ _3251_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5385_ _0718_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7124_ _2137_ _2327_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7989__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7055_ _1441_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8650__A2 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6661__A1 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5464__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _0643_ _1253_ _1295_ _1262_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__A1 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7957_ _1682_ _3128_ _2918_ _2922_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6908_ _4239_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7888_ _1658_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8166__A1 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8166__B2 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6839_ _2055_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4712__I _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9165__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6132__C _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8509_ _4243_ _4244_ _4426_ _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_109_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7141__A2 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5152__A1 _4499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8641__A2 _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7898__C _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8157__A1 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__A1 _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7132__A2 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5143__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5694__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5170_ _0506_ _0507_ _4516_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8632__A2 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7601__C _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5997__A3 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8860_ net41 _3945_ _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7811_ _2996_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8935__A3 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8791_ _3887_ _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7742_ _2303_ _2932_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8148__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4954_ _4154_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7673_ _2814_ _2649_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8699__A2 _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5628__I _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4885_ _4465_ _4466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4532__I _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6624_ _1001_ _1870_ _1875_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7371__A2 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5382__A1 _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6555_ _1768_ _1790_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5506_ _0567_ _0753_ _0816_ _0470_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_119_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9274_ _0223_ clknet_leaf_54_wb_clk_i as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6486_ _0994_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8225_ _1410_ _2475_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5134__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5437_ _4350_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5363__I _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5685__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8156_ _1555_ _3280_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5368_ _0585_ as2650.stack\[5\]\[12\] as2650.stack\[4\]\[12\] _0393_ _0704_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7107_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8087_ _1068_ _3167_ _3253_ _3254_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5299_ _4457_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8623__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5437__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7038_ _1523_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8387__A1 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8387__B2 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8989_ _1669_ _2195_ _4040_ _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8139__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5212__I2 as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5373__A1 _4467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7114__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8311__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8311__B2 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5125__A1 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6322__B1 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6468__A4 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5273__I _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6873__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6873__B2 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8614__A2 _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5428__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__I _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8378__A1 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9330__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8533__B _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5649__S _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6928__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7050__A1 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4939__A1 _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__A2 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5448__I _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4670_ _4250_ _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7353__A2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8550__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6156__A3 _4340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5364__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6340_ _1388_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8302__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6271_ _1555_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8010_ _2296_ _3177_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5222_ _0347_ _0461_ _0558_ _4212_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6864__B2 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8066__B1 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8494__I _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5153_ _0381_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8605__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5911__I _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5084_ _4161_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8912_ _3981_ _1100_ _3984_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8369__A1 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8843_ _3930_ _3931_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7041__A1 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7041__B2 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8774_ as2650.stack\[7\]\[13\] _3869_ _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _0348_ _1235_ _1276_ _1212_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7592__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7725_ _2379_ _2915_ _2916_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4937_ _4503_ _4510_ _4517_ _4518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ _2828_ _2836_ _2844_ _2849_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4868_ _4442_ _4257_ _4445_ _4448_ _4449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__7344__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _1093_ _1862_ _1864_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7587_ _2780_ _2781_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\] _4375_ _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9326_ _0275_ clknet_leaf_42_wb_clk_i as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6538_ _1778_ _1787_ _1801_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9203__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9257_ _0206_ clknet_leaf_37_wb_clk_i as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6469_ _0343_ _0983_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8844__A2 _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8208_ _1582_ as2650.stack\[1\]\[4\] as2650.stack\[0\]\[4\] _3238_ _3373_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9188_ _0137_ clknet_leaf_19_wb_clk_i net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8618__B _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8139_ as2650.pc\[2\] as2650.pc\[1\] as2650.pc\[0\] _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_87_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6607__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6083__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9021__A2 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7032__A1 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6652__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5969__I0 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8780__A1 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8532__A1 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5346__A1 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6543__B1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7099__A1 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8296__B1 _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8835__A2 _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5731__I _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8599__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__B _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5821__A2 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9012__A2 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7658__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7023__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5840_ _1140_ _1049_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7574__A2 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8771__A1 _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5771_ _1090_ _1091_ _1009_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7510_ _2647_ _1525_ _2668_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _4173_ as2650.ins_reg\[1\] _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_8490_ _3639_ _4347_ _3641_ _3643_ _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8523__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7441_ _2595_ _2438_ _2533_ _2616_ _2639_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__9226__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ _4233_ _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5906__I _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5888__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7372_ _2209_ _1415_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4584_ _4148_ _4164_ _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9111_ _0060_ clknet_leaf_51_wb_clk_i as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6323_ as2650.psl\[3\] _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8826__A2 _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9042_ _3018_ _4096_ as2650.psu\[4\] _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _0754_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5205_ _4349_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6185_ _1468_ _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8157__C _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _4436_ _0347_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _0404_ _4404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9003__A2 _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8173__B _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8826_ _1953_ _3919_ _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8757_ as2650.stack\[7\]\[7\] _3863_ _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5969_ _0476_ _1260_ _1195_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7708_ _2364_ _2899_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8688_ _1011_ _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7639_ _2757_ _2789_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5879__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9309_ _0258_ clknet_leaf_17_wb_clk_i net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8817__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5500__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5551__I _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7253__A1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6382__I _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7005__A1 _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7556__A2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8753__A1 as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9249__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7308__A2 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8505__A1 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6516__B1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A2 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__S1 _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8808__A2 _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A2 _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7244__A1 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7990_ _2267_ _3154_ _3156_ _3158_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7795__A2 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8992__A1 _4503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7388__I _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6292__I _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6872_ _0909_ _2082_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8744__A1 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8611_ _4507_ _3410_ _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5823_ as2650.r123_2\[3\]\[0\] _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8542_ _3652_ _0367_ _3691_ _3694_ _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_56_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_56_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5754_ _1076_ _1009_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_37_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7337__B _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4705_ _4285_ _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8473_ _3266_ _3620_ _3627_ _2960_ _3628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5685_ _0958_ _1012_ _1013_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7424_ net10 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4636_ _4198_ _4217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7355_ _1558_ _2395_ _2554_ _2399_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4567_ _4147_ _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6306_ _4486_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7286_ _2308_ _2487_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6467__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9025_ _3016_ _4082_ _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6286__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7072__B _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6168_ _1451_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7235__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8682__I _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5119_ _4395_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ _4192_ _4404_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7786__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8983__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8735__A1 _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5549__A1 _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8809_ _0690_ _3893_ _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5549__B2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7710__A2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7474__A1 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8806__B _4517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7226__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5237__B1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8974__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9071__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4625__I _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7001__I _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7529__A2 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8726__A1 as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8260__C _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4763__A2 _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ _0802_ _0803_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7140_ _1663_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7465__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7071_ _1671_ _2269_ _2271_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6022_ _0736_ _1227_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8965__A1 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7768__A2 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5779__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7973_ as2650.psu\[7\] _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4535__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6924_ _1512_ _1394_ _2135_ _1675_ _2138_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__6440__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _2058_ _2064_ _2080_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8193__A2 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout48 net13 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5806_ _1062_ _1120_ _1122_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6786_ _4359_ _1006_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7940__A2 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8525_ _0368_ _2373_ _3678_ _3679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5737_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5951__A1 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8456_ _3069_ _3603_ _3605_ _3611_ _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5668_ _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7407_ net1 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5703__A1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _4197_ _4199_ _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8677__I _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8387_ _2348_ _3540_ _3532_ _3128_ _3191_ _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_117_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5599_ _4389_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7338_ _2307_ _2537_ _2538_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7269_ _2439_ _2458_ _2465_ _2470_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_78_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9008_ _0871_ _0872_ _0883_ _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5034__C _4449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8405__B1 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8345__C _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__A1 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_64 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_75 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8708__A1 _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_86 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_109_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8184__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7931__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5276__I _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_1_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7447__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4681__A1 _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4970_ _4218_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8271__B _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8175__A2 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ _1883_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6186__A1 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7922__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6571_ as2650.r0\[7\] _0959_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5933__A1 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8310_ _3196_ _3471_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5522_ _0375_ _0854_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9290_ _0239_ clknet_leaf_9_wb_clk_i as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7615__B _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6489__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8241_ _3199_ _3404_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5453_ _0645_ _0603_ _0787_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5914__I _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8172_ _3325_ _3326_ _3337_ _3210_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5384_ as2650.holding_reg\[5\] _4130_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7438__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7123_ _0939_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7054_ _2251_ _2255_ _2257_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8446__B _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6005_ _1287_ _1293_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4672__A1 _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6413__A2 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7956_ _3127_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ as2650.cycle\[6\] _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7887_ _1661_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _2058_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6177__A1 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4727__A2 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6769_ _1996_ _1967_ _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8508_ _3646_ _1576_ _3660_ _3661_ _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_40_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7677__A1 _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8439_ _3343_ _3578_ _3595_ _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8929__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7601__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4966__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8157__A2 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4903__I _4483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7904__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6963__I0 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5143__A2 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6891__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8093__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7840__A1 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 io_in[33] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7810_ _2996_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8790_ as2650.r123\[1\]\[0\] _3889_ _3891_ _1701_ _3892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7741_ _2290_ _2931_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4953_ _4315_ _4329_ _4339_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4957__A2 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8148__A2 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5909__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7329__C _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7672_ _1008_ _1596_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6159__A1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4884_ _4168_ _4465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6623_ as2650.stack\[0\]\[10\] _1873_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _1768_ _1790_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5382__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7659__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5505_ _0571_ _0818_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9273_ _0222_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6485_ _0545_ _0960_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8224_ _0758_ _0652_ _3387_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5436_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6331__A1 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6331__B2 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8155_ _1554_ _0446_ _3320_ _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6882__A2 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5367_ _4495_ as2650.stack\[3\]\[12\] as2650.stack\[2\]\[12\] _4474_ _0502_ _0703_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7106_ _1056_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8086_ _2436_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5298_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ _1461_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7831__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8387__A2 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6398__A1 _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9132__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8988_ _4053_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6937__A3 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A2 _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7939_ _2222_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8139__A2 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7898__A1 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9282__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__I3 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5373__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6322__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4723__I2 as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6625__A2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8378__A2 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7050__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4939__A2 _4463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__I _4503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__C _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8550__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8302__A2 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6270_ _1554_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5221_ _4378_ _4382_ _0341_ _0345_ _4305_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_130_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__A1 _4455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8066__A1 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8066__B2 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5152_ _4499_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7813__A1 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9155__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8911_ as2650.stack\[2\]\[5\] _3982_ _3984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8369__A2 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8842_ _2091_ _3891_ _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9030__A3 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4971__C _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7041__A2 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8773_ _3825_ _3871_ _3877_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5985_ _1272_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5639__I _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5052__A1 as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7724_ net51 _2306_ _2852_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4936_ _4516_ _4517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7329__B1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7655_ _2815_ _2348_ _2848_ _2223_ _2772_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_127_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ _4271_ _4447_ _4448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_123_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8541__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6606_ as2650.stack\[5\]\[4\] _1863_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7586_ net36 _2746_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4798_ as2650.r0\[1\] _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9325_ _0274_ clknet_leaf_42_wb_clk_i as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6537_ _1782_ _1786_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5107__A2 _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9256_ _0205_ clknet_leaf_36_wb_clk_i as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6468_ _0342_ _1734_ _0982_ _0995_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8207_ as2650.stack\[6\]\[4\] _3200_ _3243_ as2650.stack\[7\]\[4\] _4497_ _3372_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_133_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8685__I _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5419_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9187_ _0136_ clknet_leaf_19_wb_clk_i net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6399_ _1674_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8057__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8618__C _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8138_ _3301_ _3304_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4718__I as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8069_ _2313_ _3226_ _3236_ _3190_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__A1 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7032__A2 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8532__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5346__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6543__B2 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8296__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7099__A2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8296__B2 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9178__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6310__A4 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8048__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6329__B _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4609__A1 as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7271__A2 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7939__I _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8263__C _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7023__A2 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8220__A1 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_opt_1_0_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8771__A2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ as2650.pc\[4\] _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_76_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\] _4301_ _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7440_ _2617_ _2621_ _2638_ _2439_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6534__A1 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4652_ _4232_ _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7371_ _2542_ _2556_ _2570_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4583_ _4149_ _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9110_ _0059_ clknet_leaf_52_wb_clk_i as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8287__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6322_ _1604_ _0350_ _1597_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5127__C _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9041_ _4097_ _4099_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6253_ _1535_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4848__A1 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8039__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5204_ _0436_ _0514_ _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_130_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6184_ _4154_ _4225_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5135_ _0346_ _0460_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5066_ _4236_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8825_ _3890_ _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8756_ _1906_ _3862_ _3866_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5968_ _1254_ _1196_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7707_ net51 _2898_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4919_ _4495_ as2650.stack\[3\]\[8\] as2650.stack\[2\]\[8\] _4474_ _4499_ _4500_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7584__I _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8687_ _3821_ _3815_ _3822_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5899_ _1175_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8514__A2 _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7638_ _2831_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7569_ _2754_ _2764_ _2751_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9308_ _0257_ clknet_leaf_16_wb_clk_i net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8278__A1 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9320__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8629__B _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9239_ _0188_ clknet_leaf_67_wb_clk_i as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8450__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8202__A1 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7005__A2 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5279__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5016__A1 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8505__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7713__B1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6516__B2 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8269__A1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7443__B _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5742__I as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8441__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7795__A3 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8992__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6940_ _1476_ _2153_ _2154_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6871_ _2094_ _2090_ _2095_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5007__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5822_ _1115_ _1126_ _1131_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8610_ _1602_ _3720_ _3758_ _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5753_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8541_ _4507_ _3249_ _3693_ _1376_ _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_124_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4704_ _4127_ _4170_ _4283_ _4284_ _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_8472_ _2182_ _2335_ _3357_ _3618_ _3626_ _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5684_ as2650.stack\[2\]\[11\] _0991_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7423_ _2606_ _0740_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4635_ _4128_ _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7180__A1 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7354_ _2395_ _2553_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_25_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _4146_ _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6305_ as2650.psu\[4\] _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7285_ _1076_ _2438_ _2471_ _2486_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5652__I _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9024_ _3015_ _4080_ _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6236_ _1369_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7483__A2 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8680__A1 _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6167_ _0935_ _1372_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8432__A1 _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5118_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7800__C _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6098_ _4191_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5246__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7786__A3 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8983__A2 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5049_ _0384_ as2650.stack\[5\]\[9\] as2650.stack\[4\]\[9\] _0387_ _0388_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6994__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8196__B1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8808_ as2650.r123\[1\]\[4\] _3889_ _3905_ _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8739_ _3855_ _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8499__A1 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7171__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7474__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5485__A1 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7710__C _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7226__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8423__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5237__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6434__B1 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6393__I _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8974__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8726__A2 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6737__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8541__C _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7438__B _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5737__I _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4641__I _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8113__I _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8269__B _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8662__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7070_ _4514_ _2273_ _1386_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5476__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ _0771_ _1287_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8414__A1 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4816__I _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8965__A2 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7972_ _4443_ _3032_ _3142_ _1031_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_94_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _0970_ _2137_ _1660_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6854_ _2060_ _2063_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout49 net25 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_5805_ as2650.stack\[0\]\[0\] _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6785_ _1981_ _2013_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5400__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7940__A3 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4551__I _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5736_ _1054_ _1035_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8524_ _3677_ _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5667_ as2650.pc\[10\] _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8455_ _3266_ _3601_ _3607_ _3310_ _3610_ _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7406_ _2604_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4618_ _4153_ _4198_ _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8386_ _3347_ _3532_ _3544_ _1639_ _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6900__A1 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5703__A2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5598_ _0921_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7337_ net53 _2377_ _1425_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4549_ _4129_ _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7268_ _2466_ _2469_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5467__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6219_ _0623_ _1502_ _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9007_ _3991_ _3996_ _4003_ _4069_ _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_89_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7199_ _2124_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8405__A1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7530__C _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8405__B2 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4690__A2 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_65 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8169__B1 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8708__A2 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_76 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_87 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7392__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9029__I _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8892__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6388__I _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7440__C _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4636__I _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6958__A1 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8271__C _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7168__B _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7383__A1 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__B _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8580__B1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7922__A3 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6570_ _1734_ _1037_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5521_ _0823_ _0507_ _4516_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8240_ _3205_ as2650.stack\[1\]\[5\] as2650.stack\[0\]\[5\] _3245_ _3404_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_121_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5452_ _0512_ _0774_ _0786_ _4285_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7615__C _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8883__A1 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8171_ _3330_ _3332_ _3336_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5383_ _0716_ _4276_ _0717_ _4162_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7122_ _2324_ _2325_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7438__A2 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8635__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7053_ _1359_ _2256_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5930__I _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8446__C _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6004_ _0686_ _1279_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6949__A1 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7955_ _4187_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7857__I _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5621__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6906_ _4235_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_54_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7886_ _3062_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _2060_ _2063_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5377__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6177__A2 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6768_ _0644_ _1024_ _1965_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8688__I _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8507_ _1435_ _2202_ _1468_ _1380_ _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_137_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5719_ _0978_ _1043_ _1044_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6699_ _1798_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7525__C _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8438_ _3593_ _3594_ _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9061__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8369_ _3343_ _3512_ _3527_ _3528_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8626__A1 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8929__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7601__A2 _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6963__I1 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8617__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8547__B _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8093__A2 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5750__I as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7840__A2 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput6 io_in[5] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9042__A1 _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4952_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7740_ _2268_ _2925_ _2930_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_91_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7671_ _2365_ _2859_ _2863_ _2368_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_71_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4883_ _4118_ _4224_ _4464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6159__A2 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _0990_ _1870_ _1874_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6553_ _1771_ _1816_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5504_ _0823_ _0337_ _0836_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7659__A2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6316__C1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6484_ _1731_ _1732_ _1738_ _1730_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9272_ _0221_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8223_ _3385_ _3354_ _3386_ _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5435_ _0635_ _0663_ _0737_ _0578_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6331__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8154_ _3275_ _3278_ _3319_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5366_ _0392_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_82_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7105_ _2308_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8085_ _3168_ _3217_ _3252_ _3214_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5297_ _0619_ _0627_ _0632_ _0628_ _0436_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_87_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6095__A1 _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7036_ _2209_ _1422_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7831__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9033__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7595__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8987_ _2231_ _4052_ _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6398__A2 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7938_ _2332_ _0409_ _1660_ _2947_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8139__A3 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7347__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7869_ _2209_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6570__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6307__C1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6322__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5771__S _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8367__B _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4723__I3 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6666__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9024__A1 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7586__A1 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6389__A2 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4914__I _4494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A2 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7338__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6849__B1 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7510__A1 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5220_ _0517_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__A2 _4452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ as2650.stack\[7\]\[10\] _0392_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8066__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6077__A1 _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5082_ _0418_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7813__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8910_ _3981_ _1093_ _3983_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9015__A1 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8841_ _0774_ _3927_ _3928_ as2650.r123\[2\]\[5\] _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7577__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__I _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7200__I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8772_ as2650.stack\[7\]\[12\] _3873_ _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7041__A3 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5984_ _0553_ _1255_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5052__A2 _4484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7723_ _2886_ _2384_ _2914_ _2724_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_75_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7329__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4935_ _4464_ _4515_ _4516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7329__B2 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7654_ _2322_ _2846_ _2847_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ _4446_ _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6605_ _1855_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7585_ net37 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5655__I _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4797_ _4377_ _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8829__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9324_ _0273_ clknet_leaf_42_wb_clk_i as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4563__A1 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6536_ _1797_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9255_ _0204_ clknet_leaf_37_wb_clk_i as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7501__A1 as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6467_ as2650.r0\[1\] _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8206_ _3196_ _3370_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7803__C _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5418_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9186_ _0135_ clknet_leaf_27_wb_clk_i net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6398_ _4184_ _4225_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8057__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8137_ _1076_ _3303_ _3033_ _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5349_ _0567_ _0552_ _0637_ _0324_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8068_ _3137_ _3217_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__A2 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9006__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7019_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8634__C _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6543__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7740__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8876__I _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7780__I _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6396__I _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__I _4489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6059__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6329__C _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4609__A2 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8544__C _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8220__A2 _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7020__I _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5034__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6231__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8560__B _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7955__I _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4720_ _4110_ _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _4137_ _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8523__A3 _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7731__A1 _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7370_ _2557_ _2569_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4582_ _4162_ _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6321_ _1429_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8287__A2 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9122__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9040_ _2231_ _4098_ _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6252_ _0815_ _1516_ _1518_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_143_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5203_ _0528_ _0530_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8039__A2 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6183_ _4294_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5134_ _0458_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7798__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9272__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5065_ as2650.r123\[0\]\[2\] _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4554__I _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8824_ _4463_ _3915_ _3917_ as2650.r123\[2\]\[0\] _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8755_ as2650.stack\[7\]\[6\] _3863_ _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5967_ _1200_ _1199_ _1258_ _1233_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7865__I _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7970__A1 _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7706_ net39 _2858_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4918_ _4498_ _4499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8686_ as2650.stack\[5\]\[10\] _3819_ _3822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5898_ _1171_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8514__A3 _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7637_ _2777_ as2650.pc\[8\] _2649_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7722__A1 _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4849_ _4420_ _4422_ _4429_ _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7568_ _2608_ _2581_ _2618_ _2752_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9307_ _0256_ clknet_leaf_16_wb_clk_i net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ as2650.r0\[1\] _1015_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7499_ _2578_ _2692_ _2693_ _2695_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9238_ _0187_ clknet_leaf_0_wb_clk_i as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4729__I _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9169_ _0118_ clknet_leaf_55_wb_clk_i as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7105__I _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7789__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7789__B2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6944__I _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8450__A2 _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6461__A1 _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5264__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7005__A3 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__A1 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7961__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4775__A1 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7713__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6516__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7713__B2 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9145__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7724__B _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8269__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9295__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5244__B _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__I _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8441__A2 _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8992__A3 _4467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _2079_ _2089_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5007__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6204__A1 _4347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ as2650.stack\[0\]\[7\] _1127_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8290__B _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8540_ _3328_ _2956_ _3692_ _4507_ _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4766__A1 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4703_ net5 _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8471_ _1350_ _3625_ _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7704__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5683_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7422_ _2618_ _2620_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4634_ _4206_ _4207_ _4214_ _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_135_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7180__A2 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7634__B _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7353_ _1288_ _0686_ _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4565_ as2650.ins_reg\[0\] _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8449__C _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6304_ as2650.psu\[3\] _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7284_ _1395_ _2479_ _2485_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9023_ _4081_ _4083_ _4084_ _3118_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4549__I _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6235_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8680__A2 _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_65_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_65_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6166_ _1450_ _0945_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6097_ _0693_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5246__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6443__B2 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5048_ _0386_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6994__A2 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8196__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8196__B2 as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8807_ _1761_ _3904_ _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6999_ _2129_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6746__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9168__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8738_ _1889_ _1854_ _1051_ _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8669_ as2650.stack\[6\]\[6\] _3806_ _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8499__A2 _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7171__A2 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8671__A2 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8423__A2 _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5237__A2 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6434__A1 as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6434__B2 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4996__A1 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8187__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6737__A2 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4922__I _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7701__A4 _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__I _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ _0741_ _1279_ _1302_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_98_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7870__B1 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8414__A2 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5228__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8965__A3 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7971_ _3138_ _3126_ _3140_ _3141_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4987__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6922_ _1682_ _2136_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9310__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6853_ _2078_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5804_ _1119_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6784_ _0715_ _0648_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6252__C _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5400__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5149__B _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8523_ _2265_ _3658_ _3669_ _3676_ _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5735_ _1058_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8454_ _3608_ _3609_ _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5666_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8350__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7405_ _1581_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4617_ _4136_ _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8385_ _3536_ _3538_ _3543_ _3183_ _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5597_ _0926_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7336_ _2492_ _2493_ _2535_ _2536_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4911__A1 _4477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4911__B2 _4478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4548_ as2650.ins_reg\[2\] _4128_ _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8102__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7267_ _2467_ _2468_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_78_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6664__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5467__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9006_ _1553_ _1524_ _1433_ _3997_ _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6218_ _0621_ _0722_ _0801_ _1493_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_77_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7198_ _2393_ _2400_ _2352_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8405__A2 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6149_ _4186_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6416__A1 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4978__A1 _4451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_55 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_66 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_77 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_88 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4742__I _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5927__B1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7392__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6195__A3 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8341__A1 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6655__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4917__I _4497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6407__A1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9333__CLK clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8947__A3 _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7080__A1 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__A1 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7907__A1 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__I _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7383__A2 _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8580__A1 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8580__B2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7922__A4 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _0850_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5146__B2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5451_ _4510_ _0781_ _0785_ _0698_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6894__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8170_ as2650.stack\[7\]\[3\] _3202_ _4498_ _3335_ _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5382_ _4276_ _0661_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7121_ _2310_ _1549_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7438__A3 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7052_ _1379_ _1670_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6003_ _0699_ _1234_ _1195_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8399__A1 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6949__A2 _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7071__A1 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7954_ _2917_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6905_ _1203_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7885_ _2221_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6836_ _2061_ _2062_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_126_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _0612_ _1023_ _1965_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8506_ _0333_ _4392_ _4514_ _1362_ _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_143_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5718_ as2650.stack\[2\]\[14\] _0957_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7126__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6698_ _1700_ _1927_ _1928_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7094__B _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8437_ _0708_ _3369_ _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9206__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5137__B2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5649_ as2650.r123\[0\]\[1\] as2650.r123_2\[0\]\[1\] _4108_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8874__A2 _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8368_ _3302_ _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7319_ _2459_ _2481_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8626__A2 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8299_ _3459_ _3430_ _3460_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_46_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7113__I _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__A1 _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5568__I _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8562__A1 _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6399__I _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8865__A2 _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6876__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8078__B1 as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8617__A2 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6628__A1 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5300__A1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5851__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput7 io_in[6] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__9042__A2 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7053__A1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6800__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _0284_ _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7670_ _2173_ _2825_ _2862_ _2719_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4882_ _4290_ _4347_ _4462_ _4463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6621_ as2650.stack\[0\]\[9\] _1873_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5367__A1 _4495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8789__I _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5367__B2 _4474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6552_ _1796_ _1815_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8305__A1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7108__A2 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8305__B2 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5503_ _4215_ _0665_ _0369_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6316__B1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9271_ _0220_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6316__C2 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6483_ _0329_ _1004_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8222_ _0674_ _0547_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6102__I _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5434_ _0483_ _0738_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7642__B _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8153_ _0453_ _0340_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5365_ _0592_ as2650.stack\[1\]\[12\] as2650.stack\[0\]\[12\] _0496_ _0701_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8608__A2 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5941__I _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6619__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7104_ _2242_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8084_ _3219_ _3250_ _3251_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5296_ _0306_ _0621_ _0631_ _0311_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6095__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ _2239_ _2225_ _1474_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9033__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__A1 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8986_ _1046_ _4043_ _4051_ _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7595__A2 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7937_ _3110_ _3111_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7868_ _2339_ _2190_ _3045_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7347__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8544__A1 _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6819_ _2026_ _2027_ _2045_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5358__A1 _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7799_ _4452_ _2986_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6307__B1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6307__C2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__I as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6947__I _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5530__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7283__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9024__A2 _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8383__B _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7035__A1 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5298__I _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5349__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5349__B2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6010__A2 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7018__I _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6849__A1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7510__A2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8558__B _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5521__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5150_ _0410_ _0437_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8066__A3 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6077__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5081_ _0412_ _0417_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_42_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9015__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6592__I _4495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8840_ _2071_ _3904_ _3929_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7577__A2 _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8771_ _3823_ _3870_ _3876_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9051__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5983_ _0556_ _1205_ _1273_ _1209_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7722_ _2902_ _2913_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4934_ _4169_ _4514_ _4515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_19_wb_clk_i clknet_opt_2_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7329__A2 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7637__B _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7653_ net52 _2768_ _2423_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4865_ _4260_ _4446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4840__I _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6604_ _1855_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _2778_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4796_ _4303_ _4376_ _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9323_ _0272_ clknet_leaf_5_wb_clk_i as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6535_ _1749_ _1798_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8829__A2 _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4563__A2 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9254_ _0203_ clknet_leaf_36_wb_clk_i as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6466_ _1731_ _1732_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7501__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8205_ _1582_ as2650.stack\[5\]\[4\] as2650.stack\[4\]\[4\] _3238_ _3370_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5512__A1 as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9185_ _0134_ clknet_leaf_17_wb_clk_i net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5671__I _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6397_ _1667_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8136_ _3302_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5348_ _0638_ _0568_ _0640_ _0356_ _0325_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_47_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8067_ _3230_ _3234_ _2971_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5279_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5815__A2 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7018_ _1670_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9006__A2 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7598__I _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7568__A2 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8969_ _2221_ _3182_ _0941_ _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8517__A1 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8650__C _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6528__B1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__I _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7740__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5503__A1 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8453__B1 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9074__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9002__B _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7559__A2 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8756__A1 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6231__A2 _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8508__A1 _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5756__I _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4650_ _4223_ _4230_ _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7731__A2 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 io_in[9] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4581_ _4161_ _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6320_ as2650.psl\[1\] _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7495__A1 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6251_ _1520_ _1534_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5491__I _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5202_ _4341_ _0523_ _0535_ _0536_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6182_ _1349_ _4513_ _0655_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7247__A1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7920__B _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5133_ _0315_ _4378_ _4382_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7798__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8995__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5064_ _4521_ _4287_ _0402_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6470__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4835__I _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8747__A1 as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8823_ _3916_ _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8754_ _1904_ _3862_ _3865_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _0452_ _1255_ _1202_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7705_ _2361_ _2894_ _2896_ _2388_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4917_ _4497_ _4498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8685_ _1000_ _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5666__I _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _1054_ _4501_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7636_ _2829_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4848_ _4425_ _4428_ _4429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7567_ _0409_ _2747_ _2762_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4536__A2 _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _4359_ _4176_ _4360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7881__I _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9306_ _0255_ clknet_leaf_16_wb_clk_i net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _0544_ _0981_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7498_ _2694_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9237_ _0186_ clknet_leaf_5_wb_clk_i as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _0994_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9168_ _0117_ clknet_leaf_54_wb_clk_i as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9097__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8119_ _3063_ _3285_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9099_ _0048_ clknet_leaf_65_wb_clk_i as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8986__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__A2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6960__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7961__A2 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7277__B _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5972__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5576__I _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__C _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7713__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7229__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8977__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7031__I _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8992__A4 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8729__A1 _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6204__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5820_ _1108_ _1126_ _1130_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _4171_ _4282_ _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8470_ as2650.pc\[14\] _1620_ _2420_ _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7165__B1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5682_ _1007_ _0965_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7421_ _2619_ _2561_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5715__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4633_ _4184_ _4117_ _4213_ _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7352_ _2550_ _2551_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7634__C _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4564_ _4138_ _4144_ _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7468__A1 _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6303_ _1582_ _4387_ _0832_ _1583_ _1586_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7283_ _1075_ _2419_ _2422_ _2484_ _1675_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9022_ _4442_ _4081_ _4084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6110__I _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6234_ _4213_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6140__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _4233_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8968__A1 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _0294_ _4420_ _4218_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6443__A2 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5047_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8196__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8806_ _3880_ _3887_ _4517_ _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6998_ _2142_ _1453_ _2196_ _2198_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8737_ _3829_ _3846_ _3854_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5954__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5949_ _0330_ _1234_ _1194_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_43_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8668_ _1904_ _3805_ _3808_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7619_ _2646_ _2812_ _2813_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8599_ _2176_ _3688_ _3746_ _3748_ _2411_ _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7116__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8959__A1 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6434__A2 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4996__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8187__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6198__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9112__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7934__A2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9262__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6370__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7026__I _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6122__A1 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8566__B _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7870__A1 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7870__B2 _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8285__C _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A1 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7970_ _4443_ _3132_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _4195_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4987__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6852_ _2076_ _2077_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5210__S _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5803_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _2004_ _2011_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8522_ _3670_ _3673_ _3674_ _3675_ _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5734_ _0973_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7689__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8453_ _2180_ _2335_ _3360_ _3604_ _2960_ _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5665_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5944__I _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7404_ _2179_ _2413_ _2599_ _2602_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4616_ as2650.ins_reg\[2\] _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8384_ _3419_ _3540_ _3531_ _2961_ _3542_ _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6361__A1 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5596_ _4238_ _0927_ _0404_ _4190_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7335_ _2382_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4547_ as2650.ins_reg\[3\] _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7266_ net29 net54 _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6113__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9005_ _1602_ _4060_ _4068_ _3970_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6217_ _0526_ _1501_ _0532_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7197_ _1551_ _2395_ _2398_ _2399_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6148_ _1368_ _1397_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6416__A2 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6079_ _4405_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9135__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4978__A2 _4453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_56 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8169__A2 _4475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_67 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_78 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_89 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9285__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8341__A2 _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6104__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7604__A1 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7080__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5091__A1 _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7907__A2 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8580__A2 _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6591__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5450_ _0784_ _0507_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5146__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5381_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7120_ _2323_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6595__I _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7843__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7051_ _2252_ _2254_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9158__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6002_ _0452_ _1235_ _1291_ _1212_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5432__C _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7953_ _3123_ _3125_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6904_ _1908_ _2114_ _2119_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7884_ _3058_ _1522_ _3060_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8020__A1 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6835_ _0716_ _2036_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6766_ _1961_ _1986_ _1994_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5717_ _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8505_ _1485_ _2125_ _2923_ _4265_ _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6697_ _1833_ _1837_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8050__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8436_ _3347_ _3578_ _3592_ _2245_ _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5137__A2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5648_ _0958_ _0977_ _0979_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8367_ _3515_ _3524_ _3525_ _3526_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _4352_ _0894_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7318_ _1084_ _2419_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8087__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8298_ _2649_ _0747_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7834__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _0454_ _0475_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4648__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7062__A2 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4753__I _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A3 _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__A1 _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8011__A1 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8562__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6573__A1 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5376__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7285__B _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5128__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6876__A2 _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8078__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9300__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8078__B2 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4928__I _4508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4639__A1 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5300__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput8 io_in[7] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5439__I0 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8563__C _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8250__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4663__I as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6800__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _0285_ _0287_ _0288_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4811__A1 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4881_ _4348_ _4461_ _4462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6620_ _1868_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6551_ _1800_ _1814_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8305__A2 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5502_ _0338_ _0827_ _0835_ _0365_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_9270_ _0219_ clknet_leaf_51_wb_clk_i as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6316__A1 _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6482_ _1714_ _1720_ _1747_ _1740_ _1728_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__6316__B2 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8221_ _0674_ _0547_ _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5433_ _4352_ _0741_ _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7923__B _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8152_ _2934_ _3311_ _3313_ _3317_ _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__8069__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5364_ _0699_ _4509_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7103_ _2306_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6619__A2 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7816__A1 _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8083_ _2244_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5295_ _0628_ _0614_ _0630_ _0309_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7034_ _4410_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9033__A3 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8473__C _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5055__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8985_ _4043_ _4050_ _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5055__B2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4573__I _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7936_ _1573_ _2264_ _2200_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4802__A1 _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7867_ _3043_ _2412_ _3044_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8544__A2 _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6818_ _2026_ _2027_ _2045_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7798_ _2180_ _2309_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6749_ _1835_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6307__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9323__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8419_ _2854_ _3553_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6858__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5530__A2 _4467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7807__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7283__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8480__A1 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5294__A1 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8232__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7035__A2 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7794__I _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5349__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6203__I _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6849__A2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7034__I _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8471__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5080_ _0412_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_97_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8293__C _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5037__A1 _4468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5489__I _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6785__A1 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5588__A2 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8770_ as2650.stack\[7\]\[11\] _3873_ _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5982_ _0560_ _1237_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7721_ _1513_ _2907_ _2912_ _1477_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4933_ _4513_ _4505_ _4514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7652_ _2830_ _2845_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4864_ _4443_ _4444_ _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6603_ _1087_ _1856_ _1861_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7583_ _2334_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ as2650.r123\[1\]\[1\] as2650.r123\[0\]\[1\] as2650.r123_2\[1\]\[1\] as2650.r123_2\[0\]\[1\]
+ _4173_ _4375_ _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_59_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6534_ _0443_ _0648_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9322_ _0271_ clknet_leaf_12_wb_clk_i as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7653__B _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6465_ _0343_ _0286_ _0983_ _0996_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_9253_ _0202_ clknet_leaf_37_wb_clk_i as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8204_ _3100_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5416_ _0746_ _0748_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_9184_ _0133_ clknet_3_3__leaf_wb_clk_i net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5512__A2 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6396_ _1671_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8135_ _3159_ _3164_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5347_ _0644_ _0337_ _0680_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8462__A1 as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8066_ _3068_ _3231_ _3232_ _3233_ _3217_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_87_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5278_ _0607_ _4130_ _0610_ _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_101_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7017_ _2222_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8214__A1 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7568__A3 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5579__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8968_ _3068_ _0952_ _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7919_ _2939_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8899_ as2650.stack\[2\]\[0\] _3976_ _3977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8517__A2 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6528__A1 as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7119__I _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5200__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8150__B1 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6700__A1 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7256__A2 _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8453__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4609__A4 as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8205__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8205__B2 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5019__A1 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6216__B1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5102__I _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8508__A2 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6519__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6361__C _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _4160_ _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5772__I _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6250_ _1359_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5201_ _0537_ _0531_ _0532_ _4338_ _4297_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6181_ _1465_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8444__A1 as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5132_ _4435_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_112_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5258__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _4288_ _0374_ _0400_ _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6108__I _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8822_ _3880_ _3914_ _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5012__I _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8753_ as2650.stack\[7\]\[5\] _3863_ _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5965_ _0456_ _1205_ _1256_ _1165_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4851__I as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7704_ _2177_ _2895_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4916_ _4496_ _4497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5896_ _1187_ _1189_ _1156_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8684_ _3818_ _3815_ _3820_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7635_ _0997_ _0830_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4847_ _4427_ _4245_ _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7566_ _2744_ _2341_ _2577_ _2162_ _2345_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4778_ _4358_ _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9305_ _0254_ clknet_leaf_16_wb_clk_i net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6517_ _1718_ _1779_ _1781_ _1754_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_134_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7497_ _1658_ _0940_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8198__C _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9236_ _0185_ clknet_leaf_33_wb_clk_i as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6448_ _0286_ _0983_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9167_ _0116_ clknet_leaf_4_wb_clk_i as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6379_ as2650.stack\[6\]\[14\] _1646_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8118_ _3262_ _3284_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8435__A1 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9098_ _0047_ clknet_leaf_65_wb_clk_i as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8049_ _3216_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7402__I _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6997__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7558__B _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7410__A2 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7174__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8910__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A2 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8674__A1 _4495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8426__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8977__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6356__C _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8729__A2 _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6204__A3 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ as2650.pc\[2\] _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _4205_ _4215_ _4231_ _4281_ _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5681_ _1008_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7165__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7165__B2 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8362__B1 _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8901__A2 _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7420_ _2539_ net10 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4632_ _4210_ _4212_ _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5715__A2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7351_ _2543_ _0574_ _2450_ _2451_ _2505_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4563_ _4141_ _4143_ _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6302_ _4477_ _1236_ _1585_ as2650.psu\[5\] _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7282_ _2323_ _2482_ _2483_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7468__A2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9021_ _3019_ _4082_ _4083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6233_ _1517_ _0792_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7931__B _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8417__A1 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _1400_ _1446_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5115_ net8 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6095_ _4210_ _1206_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_85_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5046_ _0379_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4782__S _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8481__C _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8805_ _3902_ _3903_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5677__I _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6997_ _2201_ _2203_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5403__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8736_ as2650.stack\[3\]\[14\] _3844_ _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5948_ _0368_ _1235_ _1240_ _1212_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_94_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7156__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7892__I _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8667_ as2650.stack\[6\]\[5\] _3806_ _3808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5879_ _4250_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7618_ _2780_ _2643_ _2644_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6903__A1 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5706__A2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8598_ _1575_ _3747_ _1515_ _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9064__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7549_ net35 _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7459__A2 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8656__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9219_ _0168_ clknet_leaf_22_wb_clk_i as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8408__A1 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8959__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5890__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8391__C _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__I _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7934__A3 _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8898__I _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8895__A1 _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6370__A2 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5005__S0 _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8566__C _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5881__A1 _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A2 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8582__B _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6920_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7198__B _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6851_ _2053_ _2066_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5497__I _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6189__A2 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _1046_ _1048_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6782_ _2005_ _2010_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8521_ _4141_ _1197_ _0969_ _2148_ _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__7138__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ _1057_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8886__A1 _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7689__A2 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8452_ _3357_ _3600_ _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5664_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7403_ _2600_ _0936_ _2344_ _2601_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_129_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4615_ _4142_ _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8383_ _3281_ _3541_ _2601_ _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5595_ _4189_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7217__I _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7334_ _1084_ _2239_ _1488_ _2518_ _2534_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8638__A1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5165__C _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4546_ _4118_ _4126_ _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7265_ net30 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7310__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6113__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5960__I _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8476__C _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9004_ _2215_ _4064_ _4060_ _4067_ _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6216_ _0432_ _0419_ _0423_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7196_ _2134_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6147_ _1430_ _1431_ _1380_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_100_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ _1361_ _1363_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_85_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7887__I _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5029_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_57 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_68 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_79 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5927__A2 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7836__B _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8719_ _0920_ _1049_ _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8326__B1 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8629__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5560__B1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__I as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7301__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6104__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5870__I _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A2 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5863__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7368__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6591__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7540__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6343__A2 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7037__I _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5380_ _0650_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8577__B _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5780__I _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7050_ _2253_ _1404_ _0944_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7843__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A1 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ _1272_ _1290_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9045__A1 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7952_ _4121_ _3124_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5082__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6903_ as2650.stack\[4\]\[7\] _2115_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7359__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7883_ _2748_ _3059_ _3052_ _2942_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8020__A2 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6834_ _1803_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6031__A1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _1964_ _1985_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8308__B1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8504_ _2280_ _2497_ _2288_ _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_52_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4593__A1 _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ _1030_ _1035_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6696_ _4358_ _1835_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8435_ _2970_ _3590_ _3591_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5647_ as2650.stack\[2\]\[8\] _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8366_ _0398_ _3100_ _3077_ _3511_ _2939_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5578_ _0337_ _0908_ _0910_ _4351_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7391__B _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7317_ _2496_ _2511_ _2517_ _2153_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8087__A2 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4529_ _4109_ _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8297_ _1596_ _0747_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7248_ _2448_ _2396_ _2449_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_85_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5845__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4648__A2 _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9036__A1 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7179_ _2381_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8795__B1 _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9252__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8011__A2 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6573__A2 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4584__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5086__B _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A1 _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9005__C _3970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A2 _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7589__A1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 io_in[8] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8250__A2 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6800__A3 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4811__A2 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4880_ _4440_ _4460_ _4461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6013__A1 _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7761__A1 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4575__A1 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6550_ _1802_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5501_ _0666_ _0829_ _0834_ _0363_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6316__A2 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6481_ _1730_ _1739_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8220_ _3065_ _3182_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9125__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5432_ _0651_ _4355_ _0766_ _4351_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7923__C _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8151_ _2418_ _3312_ _3315_ _3085_ _3316_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8069__A2 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5363_ _0644_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7102_ _2305_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8082_ _3235_ _3237_ _3249_ _3210_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5294_ _4310_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9275__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9018__A1 _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7033_ _2233_ _2235_ _2237_ _1437_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_45_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5015__I _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8984_ _3114_ _0492_ _4049_ _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6252__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7935_ _3107_ _3108_ _3109_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A2 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7866_ _0926_ _1422_ _1402_ _1399_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6004__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _2030_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7752__A1 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7797_ _2233_ _2985_ _2285_ _2220_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__6555__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6748_ _1975_ _1977_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6679_ _1367_ _1177_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6307__A2 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8418_ _3574_ _3575_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6858__A3 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8349_ _0966_ _3479_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7405__I _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7807__A2 _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5818__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9009__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6491__A1 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8232__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7140__I _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6243__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8783__A3 _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7991__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4557__A1 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9298__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9016__B _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8574__C _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8223__A2 _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__A2 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5981_ _1198_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7982__A1 _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7720_ net51 _2793_ _2795_ _2911_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4796__A1 _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4932_ _4309_ _4512_ _4513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5993__B1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7651_ _2765_ _2788_ _2831_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4863_ _4241_ _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4623__B _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7734__A1 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ as2650.stack\[5\]\[3\] _1857_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7582_ as2650.pc\[9\] _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4794_ _4109_ _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9321_ _0270_ clknet_leaf_63_wb_clk_i as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6533_ _0519_ _1005_ _0649_ _0329_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9252_ _0201_ clknet_leaf_43_wb_clk_i as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6464_ _0286_ _4316_ _0982_ _0996_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8203_ _3347_ _3346_ _3367_ _2245_ _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5415_ _4365_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9183_ _0132_ clknet_leaf_15_wb_clk_i as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6395_ _1442_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8134_ _3255_ _3257_ _3286_ _3298_ _3300_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_47_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5346_ _4215_ _0681_ _0369_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8462__A2 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8065_ _3035_ _3037_ _3065_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ _0612_ _4259_ _4323_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7016_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8056__I _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8214__A2 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6225__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6225__B2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7568__A4 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8967_ _0408_ _3182_ _2142_ _2694_ _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_70_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7918_ _3087_ _3090_ _3093_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8898_ _3974_ _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7849_ _3028_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7725__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__C _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5200__A2 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8150__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8150__B2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7135__I _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6700__A2 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8453__A2 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8394__C _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__A2 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6216__B2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6923__B _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7964__A1 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7738__C _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7716__A1 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6519__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5258__C _4489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8141__A1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__I _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8692__A2 _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5200_ _0294_ _4218_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4702__A1 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _4222_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8585__B _3735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5131_ _0439_ _4355_ _0468_ _4351_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5062_ _4285_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9313__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8821_ _3914_ _3915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8752_ _1900_ _3862_ _3864_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7648__C _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ _0463_ _1237_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7703_ as2650.addr_buff\[3\] _2740_ _2821_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5430__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4915_ as2650.psu\[2\] _4482_ _4496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8683_ as2650.stack\[5\]\[9\] _3819_ _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7707__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5895_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6124__I _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7634_ _2402_ _2818_ _2827_ _2758_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4846_ _4426_ _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8380__A1 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7565_ _2757_ _2760_ _2386_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4777_ as2650.r0\[7\] _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8479__C _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9304_ _0253_ clknet_leaf_2_wb_clk_i as2650.r123\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6516_ _0342_ _1717_ _1780_ as2650.r0\[0\] _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7496_ _2690_ _2526_ _2474_ _2321_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9235_ _0184_ clknet_leaf_33_wb_clk_i as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__I _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6447_ _4379_ _4316_ _0982_ _0995_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__8683__A2 _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9166_ _0115_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6378_ _1028_ _1648_ _1655_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8117_ _3034_ _3272_ _3283_ _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5329_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9097_ _0046_ clknet_leaf_65_wb_clk_i as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6446__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8048_ _2380_ _1056_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6997__A2 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7946__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7558__C _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7174__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8371__A1 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6969__I _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5185__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4932__A1 _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5113__I _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7937__A1 _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4952__I _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _4249_ _4266_ _4280_ _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5680_ _0964_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8362__A1 _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8362__B2 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4631_ as2650.alu_op\[0\] _4211_ _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5783__I _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5715__A3 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7350_ _2543_ _0574_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4923__A1 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4562_ _4142_ _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8114__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7281_ _2467_ _2426_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8665__A2 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9020_ _3058_ _1383_ _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7873__B1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6232_ _1360_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8417__A2 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6163_ _4124_ _4202_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5114_ _0451_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__C _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5045_ _0383_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7659__B _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8804_ _0583_ _3894_ _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6996_ _1435_ _1466_ _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5403__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8735_ _3827_ _3846_ _3853_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5947_ _0459_ _1201_ _1202_ _1239_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_40_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8666_ _1900_ _3805_ _3807_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8353__A1 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5878_ _4166_ _1169_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7617_ _2777_ _2727_ _2811_ _2536_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_107_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9209__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4829_ _4216_ _4232_ _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5693__I _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8597_ _0665_ _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6903__A2 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_43_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_43_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7548_ net36 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8105__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7479_ _2236_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9218_ _0167_ clknet_3_7__leaf_wb_clk_i as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8408__A2 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9149_ _0098_ clknet_leaf_66_wb_clk_i as2650.r123\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6419__A1 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5890__A2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A1 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6029__I as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7569__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__I _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__A3 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5089__B _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8344__A1 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8895__A2 _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5005__S1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6658__A1 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4947__I _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__A1 _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5881__A2 _4446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A3 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7083__A1 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6830__A1 _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4682__I _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _2055_ _2065_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5801_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_63_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5397__A1 _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6781_ _2008_ _2009_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5397__B2 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8520_ _1252_ _4278_ _1453_ _3674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5732_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7138__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8335__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8451_ _1025_ _3606_ _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5663_ as2650.r123\[0\]\[2\] as2650.r123_2\[0\]\[2\] as2650.psl\[4\] _0993_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8886__A2 _3965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7402_ _2136_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _4191_ _4194_ _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8382_ _2168_ _2236_ _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5594_ _4404_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7333_ _2519_ _2532_ _2533_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8638__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4545_ _4125_ _4126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5018__I _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7264_ _2364_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9003_ _0634_ _4065_ _4066_ _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6215_ _0301_ _0290_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7195_ _2395_ _2397_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7233__I _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6146_ _0930_ _1388_ _0696_ _1389_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6077_ _4200_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5028_ _0357_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input10_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5688__I _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8023__B1 _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_58 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_69 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8574__A1 _4508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ _4427_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8718_ _3829_ _3834_ _3842_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8326__A1 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8326__B2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8649_ _1636_ _2373_ _3795_ _2438_ _3678_ _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_103_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6888__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9181__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8629__A2 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5560__B2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4767__I _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5863__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6982__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7065__A1 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6812__A1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5615__A2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5598__I _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7368__A2 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8565__A1 _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8317__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7540__A2 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8577__C _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7481__C _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__A1 _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6000_ _0664_ _1255_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5854__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9045__A2 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8593__B _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7056__A1 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7951_ _3119_ _3120_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9054__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _1906_ _2114_ _2118_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7882_ _2282_ _2283_ _3051_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_78_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7359__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8556__A1 as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _1973_ _2056_ _2059_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_1_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _1957_ _1988_ _1992_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_56_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8308__B2 as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8503_ _3063_ _4399_ _3656_ _1632_ _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5715_ _1031_ _1040_ _1033_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__6319__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6695_ _1831_ _1847_ _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8434_ _3137_ _3578_ _3585_ _2572_ _2837_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_137_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5646_ _0957_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8365_ _3138_ _3512_ _3521_ _2573_ _2838_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5542__A1 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5577_ _0909_ _0369_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7316_ _2514_ _2516_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4528_ _4108_ _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8296_ _1189_ _3455_ _3457_ _3310_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7247_ _2440_ _0327_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__A3 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7178_ _2281_ _2282_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7047__A1 _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ _1387_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5412__S _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__C _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6977__I _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__A1 _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7286__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__A2 _4514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9077__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7038__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7589__A2 _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8786__A1 _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5121__I _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8538__A1 _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7210__A1 _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5221__B1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__A2 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5500_ _0833_ _0457_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6480_ _1727_ _1741_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8710__A1 _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5431_ _0440_ _0742_ _0765_ _4416_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6572__I0 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8150_ _1555_ _2340_ _2197_ _2172_ _1465_ _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5362_ _4127_ _0697_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7101_ _2304_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7277__A1 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8081_ _3240_ _3242_ _3248_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5293_ _0628_ _0614_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7032_ _1459_ _2236_ _1373_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7029__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8777__A1 _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8983_ _0492_ _2192_ _4048_ _3062_ _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6252__A2 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6127__I _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7934_ _2186_ _2941_ _2748_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7865_ _3039_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7201__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4870__I as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _2033_ _2043_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8342__I _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7796_ _2587_ _2984_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7752__A2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6747_ _1810_ _1976_ _1943_ _1944_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5763__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ _1908_ _1901_ _1909_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7504__A2 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8417_ _2856_ _3303_ _3033_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5629_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8348_ as2650.pc\[9\] as2650.pc\[8\] _3479_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7268__A1 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8279_ _0918_ as2650.stack\[3\]\[6\] as2650.stack\[2\]\[6\] _3331_ _4488_ _3442_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_65_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5818__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8945__C _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8961__B _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7440__A1 _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6243__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7991__A2 _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7577__B _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4780__I _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5754__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4557__A2 _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5506__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5116__I _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4955__I _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7431__A1 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5980_ _4457_ _0451_ _0570_ _0578_ _1270_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_64_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7982__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4931_ _4511_ _4512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5993__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4796__A2 _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8162__I _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7650_ _2839_ _2843_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4862_ _4423_ _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8931__A1 _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7734__A2 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6601_ _1079_ _1856_ _1860_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7581_ _2646_ _2775_ _2776_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4548__A2 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5745__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _4373_ _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9320_ _0269_ clknet_leaf_61_wb_clk_i as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6532_ _1772_ _1773_ _1789_ _1795_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_53_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9251_ _0200_ clknet_leaf_42_wb_clk_i as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6463_ _0444_ _0961_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__9242__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8202_ _2970_ _3365_ _3366_ _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5414_ as2650.r123\[1\]\[6\] as2650.r123\[0\]\[6\] as2650.r123_2\[1\]\[6\] as2650.r123_2\[0\]\[6\]
+ _4366_ _4112_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9182_ _0131_ clknet_leaf_14_wb_clk_i as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6394_ _0943_ _1384_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8133_ _3299_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _0452_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8998__A1 _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8064_ _1068_ _3176_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5276_ _0611_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_68_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_68_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4865__I _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7015_ _2191_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7670__A1 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5897__S _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7422__A1 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6225__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8966_ _2274_ _4029_ _4030_ _4032_ _4033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_102_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7917_ _0406_ _3092_ _2527_ _3089_ _3047_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5696__I _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5984__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8897_ _3974_ _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7848_ _3027_ as2650.holding_reg\[7\] _3007_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8922__A1 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7779_ net49 _2967_ _2968_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7489__A1 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7416__I _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8150__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8989__A1 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6464__A2 _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7413__A1 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6990__I _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6216__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5019__A3 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7964__A2 _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8508__A4 _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8913__A1 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9265__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6924__B1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7326__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8141__A2 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6230__I _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6152__A1 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4702__A2 _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8585__C _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5130_ _0440_ _0441_ _0467_ _4416_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5061_ _0375_ _0398_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7404__A1 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8820_ _3885_ _1367_ _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8751_ as2650.stack\[7\]\[4\] _3863_ _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5966__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5963_ _1164_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7702_ _2177_ _2893_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4914_ _4494_ _4495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6405__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8682_ _3813_ _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5894_ _0945_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8904__A1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7633_ _2542_ _2826_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4845_ as2650.addr_buff\[7\] _4426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8380__A2 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7564_ _2758_ _2759_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ as2650.psl\[3\] _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6515_ _1014_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9303_ _0252_ clknet_leaf_2_wb_clk_i as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7495_ _2690_ _2691_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7236__I _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9234_ _0183_ clknet_leaf_32_wb_clk_i as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6446_ _0414_ _0962_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9165_ _0114_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6377_ as2650.stack\[6\]\[13\] _1646_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8116_ _3274_ _3257_ _3282_ _3069_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5328_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9096_ _0045_ clknet_leaf_54_wb_clk_i as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4595__I _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7643__A1 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8047_ _1058_ _3167_ _3215_ _2982_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6446__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5259_ as2650.stack\[3\]\[11\] _4485_ _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9138__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8199__A2 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8949_ _3638_ _4016_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9288__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6315__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8530__I _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7574__C _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5185__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5375__B _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4932__A2 _4512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7146__I _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6685__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6985__I _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7882__A1 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7634__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7937__A2 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5948__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4620__A1 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7765__B _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8362__A2 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ _4139_ as2650.alu_op\[2\] as2650.ins_reg\[4\] _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4561_ as2650.alu_op\[2\] _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8114__A2 _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6300_ _0755_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7280_ _2463_ _2481_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6895__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6231_ _1360_ _4371_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7873__A1 _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7873__B2 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4687__A1 _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _4372_ _4406_ _0335_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7625__A1 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6428__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5113_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6093_ _1368_ _4181_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5304__I _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _0378_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8803_ as2650.r123\[1\]\[3\] _3901_ _3898_ _1743_ _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5939__A1 _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6995_ _4200_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8734_ as2650.stack\[3\]\[13\] _3844_ _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _1236_ _1238_ _1208_ _0361_ _1165_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_55_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8665_ as2650.stack\[6\]\[4\] _3806_ _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5877_ _1168_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8353__A2 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7616_ _1573_ _2787_ _2796_ _2797_ _2810_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4828_ _4210_ _4408_ _4409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8596_ _3744_ _3745_ _1538_ _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7547_ _2362_ _2734_ _2742_ _2354_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4759_ _4153_ _4291_ _4340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8105__A2 _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6116__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7478_ _2542_ _2663_ _2675_ _2386_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7864__A1 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9217_ _0166_ clknet_leaf_40_wb_clk_i as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7864__B2 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6429_ _1698_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_wb_clk_i clknet_3_3__leaf_wb_clk_i clknet_leaf_12_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9148_ _0097_ clknet_leaf_60_wb_clk_i as2650.r123\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7616__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7616__B2 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9079_ _0028_ clknet_leaf_46_wb_clk_i as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8959__A4 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8592__A2 _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4602__A1 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9303__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5330__A2 _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7607__A1 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7083__A2 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6830__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4841__A1 _4421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8032__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8032__B2 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8583__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5800_ _0955_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6780_ _2006_ _2007_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5731_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8335__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8450_ _1018_ _3579_ _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5662_ _0958_ _0990_ _0992_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6346__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7401_ net33 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4613_ _4192_ _4193_ _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8381_ _2426_ _2846_ _3539_ _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6897__A2 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5593_ _0922_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7332_ _1676_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4544_ _4119_ _4124_ _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7263_ _2405_ _2462_ _2464_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6214_ _0866_ _1494_ _1498_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9002_ _0633_ _4065_ _2587_ _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7194_ _0351_ _0328_ _2396_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6145_ _1365_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8271__A1 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ _4209_ _4157_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5085__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5027_ _0338_ _0348_ _0364_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7389__C _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4832__A1 _4403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8023__A1 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8023__B2 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_59 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8574__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6978_ _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8717_ as2650.stack\[4\]\[14\] _3832_ _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ as2650.r123_2\[0\]\[1\] _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8326__A2 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9326__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8648_ _1515_ _3793_ _3794_ _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8579_ _3728_ _3729_ _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4899__A1 _4476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5560__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7424__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8964__B _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8262__A1 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6812__A2 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8565__A2 _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6576__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5379__A2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8317__A2 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__A1 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5119__I _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5563__B _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5303__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7056__A2 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__I _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5067__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4693__I _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8165__I _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7950_ _3122_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__A1 _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8005__A1 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6901_ as2650.stack\[4\]\[6\] _2115_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7881_ _2991_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8556__A2 _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6832_ _2037_ _2038_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6567__A1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _1959_ _1987_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_108_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8308__A2 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8502_ _1669_ _1548_ _3655_ _3062_ _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6319__A1 _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5714_ _1039_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6319__B2 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6694_ _1832_ _1846_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8433_ _3088_ _3231_ _3580_ _3589_ _1638_ _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5645_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5029__I _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8364_ _3038_ _3512_ _3518_ _3523_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _0860_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7315_ _2515_ _2462_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4527_ as2650.psl\[4\] _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7819__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8295_ _2689_ _3456_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7295__A2 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7246_ _2440_ _0327_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7177_ _1066_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8244__A1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6128_ as2650.psu\[5\] _1411_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7047__A2 _4169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A1 as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8795__A2 _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8075__I _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6059_ _0883_ _1228_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__A2 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6323__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5367__C _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7863__B _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6730__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4778__I _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8483__A1 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5297__B2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8235__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7038__A2 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5049__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_4__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8538__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5221__A1 _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5221__B2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8710__A2 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5430_ _0363_ _0754_ _0764_ _4414_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5524__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6572__I1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6389__B _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4688__I _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5361_ _0695_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7100_ _2291_ _2303_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7277__A2 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8474__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8080_ as2650.stack\[7\]\[1\] _3243_ _4497_ _3247_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5292_ _0606_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7031_ _2206_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__A1 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7029__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8777__A2 _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7013__B _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6408__I _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5312__I _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8982_ _4044_ _4047_ _2192_ _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9171__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout53_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7933_ _4444_ _2941_ _2922_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5460__A1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7864_ _3036_ _3038_ _3040_ _3041_ _2527_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _2035_ _2042_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7795_ _2983_ _1633_ _2132_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6143__I _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6746_ _0743_ _1016_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7683__B _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__S _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6677_ as2650.stack\[3\]\[7\] _1902_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8416_ _3255_ _3555_ _3564_ _3573_ _3300_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5628_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5515__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8347_ _3506_ _3507_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5559_ _0325_ _0888_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7268__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8278_ _3327_ _3440_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7229_ _2374_ _2431_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8217__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8768__A2 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6243__A3 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__A1 _4510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__I _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5754__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6988__I _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5892__I _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5506__A2 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7900__B1 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8201__C _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8456__A1 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9194__CLK clknet_opt_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8208__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8208__B2 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6228__I _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7768__B _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5442__A1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7487__C _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4930_ _4198_ _4312_ _4511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _4441_ _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_61_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6600_ as2650.stack\[5\]\[2\] _1857_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7734__A3 _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7580_ _2744_ _2643_ _2644_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4792_ _4220_ _4372_ _4127_ _4373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6942__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6531_ _1777_ _1788_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9250_ _0199_ clknet_leaf_43_wb_clk_i as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6462_ _0414_ _0961_ _1715_ _1719_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8201_ _3137_ _3346_ _3359_ _2572_ _2837_ _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5413_ _4362_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9181_ _0130_ clknet_leaf_15_wb_clk_i as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6393_ _1550_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5307__I _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8447__A1 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8132_ _3165_ _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5344_ _0338_ _0665_ _0679_ _0365_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8998__A2 _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8063_ _2299_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5275_ _0545_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7522__I _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7014_ _2199_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7670__A2 _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5681__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6138__I _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8965_ _3724_ _2344_ _1383_ _4031_ _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_110_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7916_ _3091_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_37_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8896_ _1889_ _1048_ _1118_ _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7847_ _2186_ _1417_ _1625_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8922__A2 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6933__A1 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7778_ _2333_ _0929_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6729_ _1924_ _1950_ _1958_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8302__B _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7489__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9379_ net48 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5217__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8989__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7110__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6464__A3 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7413__A2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8610__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5887__I _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4791__I _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6924__A1 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6924__B2 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9027__C _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6152__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8429__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5571__B _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5060_ _0331_ _4510_ _4517_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7404__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8601__A1 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5797__I _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8750_ _3855_ _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5962_ _0438_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7701_ as2650.addr_buff\[3\] _2729_ _2732_ _2820_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4913_ as2650.psu\[2\] _4494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8681_ _0989_ _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8365__B1 _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5893_ _4168_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8904__A2 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7632_ _2169_ _2819_ _2825_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4844_ _4424_ _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6915__A1 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5718__A2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7563_ _2751_ _2756_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4775_ _4222_ _4207_ _4214_ _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9302_ _0251_ clknet_leaf_3_wb_clk_i as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6514_ as2650.r0\[2\] _1015_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8668__A1 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7494_ net34 net33 _2597_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9233_ _0182_ clknet_leaf_33_wb_clk_i as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6445_ _1712_ _1713_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9164_ _0113_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6376_ _1021_ _1648_ _1654_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8115_ _2596_ _3279_ _3281_ _3273_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5327_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9095_ _0044_ clknet_leaf_53_wb_clk_i as2650.stack\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7643__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8046_ _1058_ _3168_ _3213_ _3214_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5258_ _0584_ _0593_ _0594_ _4489_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ _0412_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8948_ as2650.carry _4005_ _4015_ _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8879_ _0699_ _3958_ _3960_ _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7159__B2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7882__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4786__I _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7162__I _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8831__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7398__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5410__I _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6070__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4620__A2 _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9038__B _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7570__A1 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6373__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4560_ _4140_ _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4923__A3 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6230_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7873__A2 _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4687__A2 _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5884__A1 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4696__I _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6161_ _1445_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _0445_ _0447_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_97_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8822__A1 _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6092_ _4114_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _0381_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7389__A1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7389__B2 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8802_ _3888_ _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6994_ _2199_ _2200_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8733_ _3825_ _3846_ _3852_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8889__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8664_ _3798_ _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7615_ _2542_ _2806_ _2809_ _2385_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4827_ _4407_ _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7561__A1 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8595_ _1517_ _0557_ _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7546_ _2735_ _2741_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4758_ _4308_ _4321_ _4324_ _4339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7477_ _2668_ _2670_ _2674_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6116__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4689_ _4117_ _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9105__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9216_ _0165_ clknet_leaf_40_wb_clk_i as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ _1693_ _1694_ _1697_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_88_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7864__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5875__A1 _4403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9147_ _0096_ clknet_leaf_60_wb_clk_i as2650.r123\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6359_ _1608_ _1483_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9078_ _0027_ clknet_leaf_45_wb_clk_i as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9255__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8029_ _3196_ _3197_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_52_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7092__A3 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5230__I _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6052__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4602__A2 _4182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7304__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6010__B _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8804__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5618__A1 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7083__A3 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7620__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6236__I _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7791__A1 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ as2650.pc\[0\] _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ as2650.stack\[2\]\[9\] _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7543__A1 _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7400_ _2596_ _2598_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9128__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ as2650.cycle\[0\] _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8380_ _2814_ _2320_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5592_ _4390_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7331_ _2525_ _2530_ _2531_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ as2650.cycle\[1\] _4123_ _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7262_ _2460_ _2407_ _2463_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7846__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9001_ _4334_ _0621_ _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9048__A1 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9278__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6213_ _1493_ _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7193_ _1203_ _4437_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5315__I _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ as2650.psl\[6\] _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _1359_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5085__A2 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6282__A1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5026_ _4414_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8023__A2 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6034__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7782__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8716_ _3827_ _3834_ _3841_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5928_ _1153_ _1181_ _1221_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8647_ _1547_ _3794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5859_ as2650.r123_2\[0\]\[0\] _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8578_ _2171_ _1548_ _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7529_ _2690_ _2434_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7837__A2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5848__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9039__A1 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6812__A3 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6576__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7773__A1 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4587__A1 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7525__A1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5839__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__A3 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__A2 _4404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4814__A2 _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _1904_ _2114_ _2117_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8005__A2 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7880_ _2993_ _3032_ _3057_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6016__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ _2056_ _2057_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6567__A2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8181__I _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6762_ _1265_ _1911_ _1913_ as2650.r123_2\[2\]\[2\] _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8501_ _1538_ _0441_ _3654_ _1546_ _3655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5713_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7516__A1 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6319__A2 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6693_ _1770_ _1828_ _1923_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8432_ _3583_ _3588_ _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5644_ _0962_ _0965_ _0975_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8363_ _3519_ _3522_ _3010_ _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5575_ _0440_ _0906_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7314_ _1073_ _0453_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4526_ as2650.r123\[0\]\[0\] _4107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7819__A2 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4750__A1 _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8294_ _1104_ _3424_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7245_ _1553_ _2389_ _2127_ _2446_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_49_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5045__I _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__I0 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7176_ _2305_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A2 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6255__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _1227_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7755__A1 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6604__I _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7507__A1 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8180__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6730__A2 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7170__I _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7994__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8215__B _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7746__A1 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5221__A2 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4980__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4732__A1 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ _4145_ _4167_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5291_ _0620_ _0625_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6485__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7030_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8176__I _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8226__A2 _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9316__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7013__C _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8981_ _4466_ _0491_ _4046_ _1624_ _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7985__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7932_ _3105_ _3106_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5460__A2 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout46_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7863_ _3039_ _4254_ _3036_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _2041_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7794_ _2629_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6745_ _1939_ _1972_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6676_ _1114_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8415_ _0597_ _3101_ _3571_ _3114_ _3572_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5627_ as2650.r123\[0\]\[0\] as2650.r123_2\[0\]\[0\] _4109_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8346_ _0968_ _3303_ _3033_ _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5558_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5771__I0 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8277_ _0494_ as2650.stack\[1\]\[6\] as2650.stack\[0\]\[6\] _3328_ _3440_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5489_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7228_ _2386_ _2401_ _2410_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_132_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8086__I _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7159_ _2354_ _2356_ _2360_ _2362_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8019__C _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7976__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5451__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7874__B _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8153__A1 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7900__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7900__B2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4714__A1 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_7_wb_clk_i clknet_3_3__leaf_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__B _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7719__A1 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ _4113_ _4441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _4166_ _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6942__A2 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8599__C _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _1793_ _1794_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4953__A1 _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8144__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6461_ _4317_ _1005_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8695__A2 _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8200_ _3088_ _3231_ _3348_ _3364_ _1416_ _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5412_ as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\] _0657_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9180_ _0129_ clknet_leaf_15_wb_clk_i as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6392_ _1667_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8131_ _3287_ _3258_ _3297_ _3101_ _2940_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5343_ _0666_ _0673_ _0678_ _0338_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8447__A2 _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8062_ _3036_ _3223_ _3229_ _1577_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5274_ _4275_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7013_ _2189_ _2214_ _2219_ _1644_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5681__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8964_ _1188_ _2292_ _2242_ _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6630__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5433__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7915_ _2344_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8895_ _3957_ _3972_ _3973_ _3970_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7846_ _2997_ _3024_ _3025_ _3026_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_58_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7777_ _1456_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4989_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6933__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _1926_ _1949_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4944__A1 _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8135__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8302__C _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6659_ _1078_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8686__A2 _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9378_ net46 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8329_ _2615_ _3484_ _3489_ _3064_ _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8438__A2 _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7110__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6464__A4 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5672__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5424__A2 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6064__I _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8374__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6999__I _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A1 _4464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8126__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8126__B2 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5408__I as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9161__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5360__A1 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6860__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4982__I _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8601__A2 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6612__A1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5415__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _1229_ _1230_ _1252_ _4279_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7700_ _2890_ _2891_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4912_ _4474_ _4492_ _4493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8680_ _3811_ _3815_ _3817_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5892_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8365__A1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8365__B2 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7631_ _2821_ _2824_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4843_ _4423_ _4267_ _4424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6915__A2 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7562_ _2563_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8117__A1 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _4230_ _4355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9301_ _0250_ clknet_leaf_1_wb_clk_i as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6513_ _0715_ _0961_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7493_ net35 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9232_ _0181_ clknet_leaf_29_wb_clk_i as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6679__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6444_ _1247_ _1705_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9163_ _0112_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6375_ as2650.stack\[6\]\[12\] _1650_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8114_ _1552_ _3280_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5326_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9094_ _0043_ clknet_leaf_53_wb_clk_i as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8045_ _3165_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5257_ as2650.stack\[2\]\[11\] _4476_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8840__A2 _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5053__I _4483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7689__B _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _0417_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6603__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8947_ _4010_ _4014_ _4005_ _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8356__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8878_ _0553_ _3959_ _3960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7829_ _3013_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9184__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8108__A1 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8032__C _4488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8659__A2 _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7882__A3 _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7095__A1 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8292__B1 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5898__I _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7398__A2 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8207__C _4497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8595__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5138__I _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6678__B _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4977__I _4522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5333__A1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5884__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6160_ _4233_ _4126_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5111_ _4365_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7086__A1 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _4206_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6833__A1 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5042_ _0377_ _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5601__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7389__A2 _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8586__A1 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8801_ _3899_ _3900_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6993_ _0334_ _1381_ _2143_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_129_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6061__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8732_ as2650.stack\[3\]\[12\] _3848_ _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5944_ _1204_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8338__A1 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8663_ _3798_ _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5875_ _4403_ _4117_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6432__I _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7614_ _2758_ _2808_ _2782_ _2402_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4826_ as2650.alu_op\[0\] _4261_ _4407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8594_ _3705_ _1016_ _3743_ _1520_ _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7545_ _2740_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4757_ _4295_ _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5048__I _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7476_ _2466_ _2673_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ _4268_ _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8510__A1 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8510__B2 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6427_ _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5324__A1 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9215_ _0164_ clknet_leaf_39_wb_clk_i as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9146_ _0095_ clknet_leaf_57_wb_clk_i as2650.r123\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5875__A2 _4117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6358_ _1630_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ as2650.r123\[0\]\[5\] _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8274__B1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9077_ _0026_ clknet_leaf_46_wb_clk_i as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6289_ _1572_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8028_ _0383_ as2650.stack\[1\]\[0\] as2650.stack\[0\]\[0\] _0386_ _3197_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8577__A1 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8329__A1 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5563__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7304__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_2_0_wb_clk_i_I clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__I _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7173__I _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6010__C _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7068__A1 _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8804__A2 _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7901__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5421__I _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7240__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5296__C _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ _0956_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4611_ as2650.cycle\[1\] _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5554__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5591_ _4512_ _4362_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7330_ _1155_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4542_ as2650.cycle\[3\] _4120_ _4122_ _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_50_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7261_ _1073_ _2167_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7846__A3 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9000_ _3718_ _1539_ _4063_ _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6212_ _0802_ _1495_ _1496_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7192_ _2394_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9048__A2 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7059__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6143_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8907__I _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7811__I _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5609__A2 _4182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6074_ _0921_ _0670_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8128__B _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7032__B _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6427__I _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5025_ _0353_ _0354_ _0362_ _0363_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_73_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8559__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6976_ _1581_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7782__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8715_ as2650.stack\[4\]\[13\] _3832_ _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5927_ _1186_ _1191_ _1217_ _1219_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ _1043_ _1144_ _1152_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8646_ _3713_ _0905_ _1518_ _3792_ _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8731__A1 _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _4128_ _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5789_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8577_ _3718_ _0742_ _3727_ _1574_ _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7528_ _2689_ _2384_ _2723_ _2724_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7207__B _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7459_ _0756_ _0770_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__9222__CLK clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5848__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9039__A2 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8247__B1 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9129_ _0078_ clknet_leaf_55_wb_clk_i as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6337__I _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8980__C _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6025__A2 _4510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8970__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4587__A2 _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5536__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7289__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5839__A2 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5303__A4 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8238__B1 _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7213__A1 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4990__I _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6830_ _4358_ _0649_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6761_ _1955_ _1990_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4578__A2 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7078__I _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5712_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8500_ _1516_ _3653_ _1535_ _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _0612_ _1006_ _1829_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7516__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8431_ _3357_ _3577_ _3585_ _3224_ _3587_ _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5643_ _0968_ _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__9245__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7806__I _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8362_ _2784_ _3222_ _3521_ _3419_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5574_ _4356_ _0754_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7313_ _2512_ _2513_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4525_ net50 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8293_ _2574_ _3450_ _3453_ _3454_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4750__A2 _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5326__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7244_ _2443_ _2444_ _2445_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7175_ _2307_ _2376_ _2378_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ _1230_ _1382_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7452__A1 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6157__I _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6255__A2 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6057_ _0891_ _1253_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5008_ _0346_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5996__I _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7204__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8305__C _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7755__A2 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8952__A1 _4494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6959_ _1556_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7507__A2 _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5518__A1 _4494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8629_ _1575_ _4370_ _3776_ _3688_ _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5518__B2 _4473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8180__A2 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6620__I _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7691__A1 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7691__B2 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7451__I _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7443__A1 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6067__I _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9118__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7994__A2 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7746__A2 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9268__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4980__A2 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6182__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4732__A2 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5290_ _0616_ _0624_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7682__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7682__B2 _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8980_ _0382_ _0971_ _4045_ _1187_ _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7985__A2 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7931_ _0927_ _2283_ _4188_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8192__I _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7862_ _3039_ _1659_ _2476_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8934__A1 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8934__B2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6813_ _2039_ _2040_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7793_ _2966_ _2980_ _2981_ _2982_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _1843_ _1973_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _1906_ _1901_ _1907_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4971__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8414_ _3503_ _3555_ _3342_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5626_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8345_ _3255_ _3481_ _3502_ _3505_ _3300_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5557_ _0825_ _0635_ _0886_ _4454_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5920__A1 _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5771__I1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8276_ _0381_ _3438_ _4498_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5488_ _0745_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7673__A1 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4895__I _4475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7227_ _1068_ _2411_ _2416_ _2429_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7158_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8217__A3 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7425__A1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6109_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7089_ _0663_ _0761_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7976__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5987__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8316__B _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6615__I _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8925__A1 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5739__A1 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8153__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6350__I _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6164__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7900__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4714__A2 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__A1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9090__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7719__A2 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4650__A1 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8740__I _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _4357_ _4370_ _4336_ _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6942__A3 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8144__A2 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6260__I _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6460_ _1707_ _1721_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5411_ _0745_ _4176_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6391_ _1666_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8130_ _3296_ _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5342_ _0677_ _0457_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7655__A1 _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8061_ _3224_ _3226_ _3228_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7655__B2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5273_ _0608_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7012_ _2215_ _2217_ _2218_ _2214_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7024__C _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5130__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8080__A1 as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8963_ _4393_ _2253_ _3992_ _1474_ _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7914_ _3043_ _2145_ _3089_ _3086_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5479__C _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8894_ net21 _3962_ _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7845_ as2650.holding_reg\[6\] _2998_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6394__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7776_ _2303_ _2965_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4988_ _0315_ _4522_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_71_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6727_ _1918_ _1952_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4944__A2 _4522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8135__A2 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6170__I _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6146__A1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ _1894_ _1891_ _1895_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7894__A1 _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5609_ _0293_ _4182_ _4261_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_9377_ net46 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6589_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8328_ _3085_ _3486_ _3487_ _3488_ _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7646__A1 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8259_ _3420_ _3421_ _2601_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8825__I _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8071__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8071__B2 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6621__A2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A1 _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A1 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6924__A3 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__A2 _4515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__B1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__A2 _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7637__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5112__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6860__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8062__A1 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6612__A2 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5960_ _4268_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_80_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4623__A1 _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4911_ _4477_ as2650.stack\[1\]\[8\] as2650.stack\[0\]\[8\] _4478_ _4492_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5891_ _1182_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8365__A2 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7630_ _2822_ _2823_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4842_ _4235_ _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5179__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6376__A1 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8403__C _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7561_ _2751_ _2756_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4773_ _4353_ _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9300_ _0249_ clknet_leaf_1_wb_clk_i as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6512_ _1751_ _1775_ _1776_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6128__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7492_ _1110_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9231_ _0180_ clknet_leaf_30_wb_clk_i as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7876__A1 _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6679__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6443_ as2650.r123_2\[1\]\[1\] _1699_ _1711_ _1703_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9162_ _0111_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6374_ _1012_ _1647_ _1653_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5351__A2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7628__A1 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8113_ _0407_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5325_ _0660_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7035__B _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9093_ _0042_ clknet_leaf_53_wb_clk_i as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8044_ _3193_ _3211_ _3212_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5256_ _0592_ as2650.stack\[1\]\[11\] as2650.stack\[0\]\[11\] _0586_ _0593_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ _0522_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8053__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6165__I _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7800__A1 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8946_ _3718_ _4398_ _4013_ _2317_ _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4614__A1 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8877_ _3940_ _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8356__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7828_ _3012_ as2650.holding_reg\[2\] _3007_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6367__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9329__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7759_ _2948_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8108__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6119__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7867__A1 _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7619__A1 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8983__C _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8292__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7095__A2 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8292__B2 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8044__A1 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8595__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8504__B _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6358__A1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5419__I _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7570__A3 _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5581__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5333__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5154__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ as2650.r123\[1\]\[3\] as2650.r123\[0\]\[3\] as2650.r123_2\[1\]\[3\] as2650.r123_2\[0\]\[3\]
+ _4366_ _4111_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_48_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8283__A1 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _0694_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5097__B2 _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _0378_ _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4993__I _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8586__A2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8800_ _0488_ _3894_ _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6597__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6992_ _4114_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8731_ _3823_ _3845_ _3851_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5943_ _0350_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8414__B _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8338__A2 _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8662_ _1898_ _3799_ _3804_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5874_ _0935_ _1166_ _1167_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7613_ _2789_ _2807_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _4404_ _4405_ _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8593_ _3740_ _3741_ _3647_ _3742_ _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5021__A1 _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5329__I _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7544_ _2737_ _2739_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4756_ _4336_ _4330_ _4337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7475_ _2671_ _2672_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4687_ _4235_ _4267_ _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8510__A2 _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9214_ _0163_ clknet_leaf_39_wb_clk_i as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6426_ _1695_ _1177_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5324__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9145_ _0094_ clknet_leaf_59_wb_clk_i as2650.r123\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6357_ _1632_ _1635_ _1640_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5308_ _0612_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _1512_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9076_ _0025_ clknet_leaf_56_wb_clk_i as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8027_ _3195_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5239_ _4431_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8308__C _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6037__B1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8577__A2 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8929_ _1378_ _1477_ _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_61_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6760__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8501__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8265__A1 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7068__A2 _4504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7403__B _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__A1 as2650.alu_op\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8017__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8234__B _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4610_ _4188_ _4189_ _4190_ _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5590_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6751__A1 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5554__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4541_ as2650.cycle\[7\] as2650.cycle\[6\] _4121_ as2650.cycle\[4\] _4122_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7260_ _2459_ _2461_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5306__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6503__A1 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6211_ _0799_ _0797_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7191_ _4428_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _4284_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7059__A2 _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4937__B _4517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8195__I _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _0921_ _4291_ _4138_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_97_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _4373_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8559__A2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ _2183_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7539__I _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5242__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8714_ _3825_ _3834_ _3840_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5926_ _1179_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7983__B _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8645_ _1576_ _3791_ _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5857_ as2650.stack\[1\]\[14\] _1142_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8731__A2 _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _4193_ _4388_ _4389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6742__A1 _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8576_ _3719_ _3690_ _3725_ _3726_ _3713_ _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5788_ _1102_ _1081_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7527_ _2382_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4739_ _4319_ _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7274__I _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8495__A1 _4478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7458_ _1596_ _0820_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ _1553_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7389_ _2541_ _2575_ _2585_ _2586_ _2588_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8247__A1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9128_ _0077_ clknet_leaf_2_wb_clk_i as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8247__B2 _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9059_ _0008_ clknet_leaf_48_wb_clk_i as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4808__A1 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7470__A2 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5481__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7449__I _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8054__B _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__A1 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8970__A2 _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5397__C _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6981__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8989__B _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A2 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8501__C _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7184__I _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__I _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7912__I _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8238__A1 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8238__B2 _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8410__A1 _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7213__A2 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6263__I _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6760_ _1915_ _1989_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6972__A1 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5775__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5711_ _4110_ _0788_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6691_ _1920_ _1921_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8713__A2 _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8430_ _2216_ _3586_ _2150_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5642_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8361_ _1621_ _2792_ _3520_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _0899_ _0903_ _0905_ _4223_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7312_ _2491_ net9 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8477__A1 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8292_ _1544_ _2335_ _2197_ _2187_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7243_ _2443_ _2444_ _4278_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8229__A1 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7174_ _2337_ _2377_ _1425_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6125_ _1410_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6255__A3 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7452__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6056_ _1175_ _1341_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8653__I _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5007_ _0341_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_113_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8401__A1 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7204__A2 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6173__I _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8952__A2 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _2167_ _2159_ _2170_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5766__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ net6 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6889_ as2650.stack\[4\]\[1\] _2109_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8704__A2 _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8628_ _1520_ _3747_ _3772_ _3775_ _3713_ _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_8559_ _1517_ _1200_ _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8468__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7691__A2 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7443__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7179__I _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8943__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5757__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6706__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8459__A1 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7682__A2 _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6258__I _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8631__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5445__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7930_ _4238_ _4120_ _0943_ _3039_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7861_ _1442_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7198__A1 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9212__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8934__A2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7737__A3 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6812_ _0793_ _1843_ _1973_ _2005_ _2010_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_7792_ _2436_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5748__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ as2650.r0\[7\] _1015_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7817__I _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ as2650.stack\[3\]\[6\] _1902_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8413_ _3567_ _3570_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7370__A1 _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8344_ _2940_ _3504_ _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5556_ _0317_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7122__A1 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8275_ as2650.stack\[5\]\[6\] as2650.stack\[4\]\[6\] _4468_ _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7552__I _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5487_ _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7226_ _2380_ _2419_ _2423_ _2428_ _1676_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7673__A2 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7157_ _2134_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7425__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6108_ _4206_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7088_ _2191_ _0923_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _0841_ _1243_ _1302_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_73_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8386__B1 _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8925__A2 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5739__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6936__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7361__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5247__I _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__A2 _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5675__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8613__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8507__B _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9235__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6027__B _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8916__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4650__A2 _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__I _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6155__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5410_ _0744_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6390_ _4270_ _1416_ _1657_ _1665_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5341_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4961__I0 _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7655__A2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8060_ _0352_ _2338_ _2417_ _3216_ _3227_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_86_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8852__A1 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5272_ _0546_ _0548_ _0550_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_86_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7011_ _4193_ _4250_ _0928_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8604__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8417__B _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8080__A2 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8962_ _1624_ _1381_ _1357_ _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6091__A1 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout51_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7913_ _3088_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8893_ _0862_ _3958_ _3971_ _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7844_ _1102_ _1634_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6918__A1 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7775_ _2964_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7591__A1 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ _0315_ _0324_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6394__A2 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6726_ _1922_ _1951_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4795__I3 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6657_ as2650.stack\[3\]\[1\] _1892_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6146__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9108__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5608_ _4185_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9376_ net46 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7894__A2 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6588_ _1824_ _1826_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_139_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8327_ _2315_ _3480_ _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5539_ _0866_ _0870_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8258_ _2182_ _3280_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5657__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9258__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7209_ _1658_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_15_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8189_ _3352_ _3320_ _3353_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8046__C _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A2 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9020__A1 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A1 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A2 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8997__B _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6137__A2 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7334__B2 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5896__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4699__A2 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8288__I _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7192__I _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5705__I _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7637__A2 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8834__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6860__A3 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8237__B _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8062__A2 _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6073__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4623__A2 _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9011__A1 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4910_ as2650.stack\[7\]\[8\] _4485_ _4490_ _4491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5890_ _1170_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4841_ _4421_ _4207_ _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7573__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6376__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6271__I _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ _2754_ _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5584__B1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4772_ _4317_ _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6511_ _1735_ _1756_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7491_ _2646_ _2687_ _2688_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6128__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9230_ _0179_ clknet_3_7__leaf_wb_clk_i as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6442_ _1707_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5336__B1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7876__A2 _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9161_ _0110_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6373_ as2650.stack\[6\]\[11\] _1650_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8112_ _3275_ _3278_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5324_ _4151_ _0649_ _0654_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_138_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9092_ _0041_ clknet_leaf_52_wb_clk_i as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8043_ _2244_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5255_ _0384_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7830__I _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5186_ _0514_ _0521_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8053__A2 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5350__I _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8945_ _3719_ _1636_ _4011_ _4012_ _1575_ _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9002__A1 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8876_ _3940_ _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8356__A3 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7827_ _2167_ _3009_ _3011_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7564__A1 _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6367__A2 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6181__I _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7758_ _2292_ _2418_ _2947_ _0940_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _1806_ _1843_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6119__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7689_ _2857_ _2186_ _1676_ _2881_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_137_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7867__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5878__A1 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9080__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5525__I as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8292__A2 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6055__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8571__I _4506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7555__A1 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__I _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7307__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7915__I _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6040__B _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5333__A3 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__A1 as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8807__A1 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7086__A3 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6294__A1 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5097__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ _4470_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6266__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6991_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8730_ as2650.stack\[3\]\[11\] _3848_ _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5942_ _1202_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8661_ as2650.stack\[6\]\[3\] _3800_ _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7546__A1 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5873_ _4233_ _4227_ _4372_ _4277_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__9229__D _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7612_ _2790_ _2757_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5557__B1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4824_ _4388_ _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8592_ _3722_ _3376_ _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7543_ _4277_ _2738_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4755_ as2650.psl\[3\] _4335_ _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8430__B _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7474_ _2600_ _2597_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4686_ _4237_ _4240_ _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9213_ _0162_ clknet_3_7__leaf_wb_clk_i as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6425_ _1454_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5345__I _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9144_ _0093_ clknet_leaf_59_wb_clk_i as2650.r123\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6356_ _0861_ _1565_ _1637_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5307_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9075_ _0024_ clknet_leaf_56_wb_clk_i as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8274__A2 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6287_ _1428_ _1484_ _1571_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5088__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6285__A1 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8026_ _3194_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5238_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _4508_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6037__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6037__B2 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7785__A1 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8928_ _3992_ _3993_ _2921_ _3995_ _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8859_ _3938_ _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6760__A2 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5255__I _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8265__A2 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7068__A3 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6276__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7403__C _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6086__I _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8234__C _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7528__A1 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7528__B2 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6200__A1 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7645__I _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6751__A2 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5554__A3 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ as2650.cycle\[5\] _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6210_ _0721_ _0723_ _0806_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7190_ _1551_ _2387_ _2388_ _2392_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _1409_ _1423_ _1426_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _1348_ _1357_ _0930_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8008__A2 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ _0354_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5490__A2 _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6974_ _1689_ _2182_ _2158_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5242__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8713_ as2650.stack\[4\]\[12\] _3836_ _3840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7519__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8644_ _3787_ _3790_ _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ _1028_ _1144_ _1151_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7983__C _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _4236_ _4191_ _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8575_ _3705_ _1007_ _3719_ _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5787_ _1105_ _0974_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6742__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7526_ _2317_ _2697_ _2706_ _2722_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_120_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4738_ _4159_ _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7457_ _1560_ _2358_ _2654_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4669_ _4181_ _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6408_ _0938_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7388_ _2587_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9127_ _0076_ clknet_leaf_0_wb_clk_i as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8247__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6339_ _1578_ _1618_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7290__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5803__I _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9058_ _0007_ clknet_leaf_8_wb_clk_i as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A2 _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8009_ _3177_ _2310_ _2297_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7758__A1 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7758__B2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6430__A1 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6981__A2 _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8183__A1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7930__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6497__A1 as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8238__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5713__I _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5472__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7213__A3 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6421__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5224__A2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5710_ _4109_ as2650.r123_2\[0\]\[6\] _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6690_ _1799_ _1849_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8174__A1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5641_ _4270_ _0970_ _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4999__I _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8360_ _0986_ _3171_ _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7308__C _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5572_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7311_ _2491_ net9 _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8291_ _3224_ _3452_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7242_ _0455_ _0485_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9141__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4948__B _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__A1 as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7173_ _2304_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8229__A2 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_1__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6124_ _0758_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7988__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9291__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _0894_ _1243_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6255__A4 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5006_ _0343_ _4175_ _4365_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__5463__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8401__A2 _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6412__A1 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7994__B _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6957_ _2169_ _2163_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4974__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5908_ _1198_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6888_ _1888_ _2108_ _2110_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4974__B2 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8627_ _4508_ _3443_ _3774_ _3724_ _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5839_ _0496_ _0919_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8558_ _3705_ _0996_ _3709_ _3652_ _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7509_ _2322_ _2703_ _2705_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8489_ _3139_ _4459_ _2370_ _3642_ _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7979__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8640__A2 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8065__B _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6403__A1 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5201__C _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8156__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6706__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9164__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6182__A3 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5142__A1 _4455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6890__A1 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7434__A3 _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8631__A2 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5445__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6274__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7860_ _3037_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7198__A2 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8395__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _1973_ _2037_ _2038_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7791_ net49 _2966_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6742_ _4358_ _0995_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4956__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8147__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6673_ _1107_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8698__A2 _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8412_ _3064_ _3310_ _3569_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5624_ _0920_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7370__A2 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8343_ _4501_ _3444_ _3503_ _3481_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5555_ _0824_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8274_ as2650.stack\[6\]\[6\] _3331_ _3202_ as2650.stack\[7\]\[6\] _3437_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5486_ _0635_ _0752_ _0816_ _0578_ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7122__A2 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _2323_ _2425_ _2427_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5133__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8870__A2 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5684__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7156_ _2120_ _2359_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7989__B _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _1365_ _1374_ _1392_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_100_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8664__I _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8622__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7087_ _2278_ _2290_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6038_ _1323_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8386__A1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8386__B2 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7989_ _1357_ _3157_ _2287_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6936__A2 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6912__I _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8689__A2 _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5528__I _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7361__A2 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5372__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7743__I _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7649__B1 _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8310__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5124__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8861__A2 _3944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5675__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6872__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8613__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6624__A1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8507__C _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6094__I _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8377__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8749__I _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5340_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8301__A1 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__I1 _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6269__I _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5271_ as2650.holding_reg\[4\] _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8852__A2 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7010_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8484__I _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8604__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8961_ _4026_ _4027_ _2222_ _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_95_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5122__B _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6091__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7912_ _3035_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8892_ _1636_ _3959_ _3971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7843_ _1689_ _1417_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6918__A2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4986_ _4243_ _4432_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7774_ _2258_ _2263_ _2955_ _2963_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_51_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7591__A2 _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6725_ _1247_ _1911_ _1913_ as2650.r123_2\[2\]\[1\] _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _1070_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8540__A1 _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6146__A3 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _0938_ _0924_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6587_ _1799_ _1849_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8326_ _2162_ _2677_ _2198_ _1550_ _1577_ _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_121_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _0866_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8257_ _1525_ _2236_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _0731_ _0727_ _0730_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6303__B1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7208_ _4410_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8188_ _0554_ _0446_ _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7139_ _2337_ _2339_ _2342_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6907__I as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_55_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8359__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9020__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8062__C _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5593__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8997__C _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7334__A2 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8569__I _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7473__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__A2 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7098__A1 _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9202__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8598__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6073__A2 _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5820__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9011__A2 _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7022__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ _4172_ _4421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7573__A2 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _4351_ _4352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5584__B2 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5168__I _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6510_ _1735_ _1756_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7490_ _2671_ _2643_ _2644_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6441_ _1708_ _1709_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6533__B1 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5336__B2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9160_ _0109_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _1001_ _1647_ _1652_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8111_ _3220_ _3276_ _3277_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7089__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5323_ _0655_ _0656_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_9091_ _0040_ clknet_leaf_53_wb_clk_i as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8042_ _1058_ _3077_ _3209_ _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6836__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5254_ as2650.stack\[7\]\[11\] _4485_ _4490_ _0590_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5185_ _0514_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5631__I _4421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8589__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7261__A1 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8944_ _4354_ _3010_ _1578_ _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9002__A2 _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8875_ _3938_ _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8210__B1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7826_ _0439_ _3010_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5414__I2 as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7757_ _1616_ _2420_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4969_ _4310_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6708_ _0650_ _1780_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7688_ _2423_ _2880_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8513__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9225__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ as2650.r123\[3\]\[3\] _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7226__C _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8309_ _1582_ as2650.stack\[1\]\[7\] as2650.stack\[0\]\[7\] _3238_ _3471_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9289_ _0238_ clknet_leaf_9_wb_clk_i as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8338__B _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7252__A1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5802__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7004__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8201__B1 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5566__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5110__S0 _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7307__A2 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8504__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5318__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A2 _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4541__A2 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8807__A2 _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8248__B _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7491__A1 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6294__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7243__A1 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6046__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6990_ _2130_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8991__A1 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7378__I _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_0_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8660_ _1896_ _3799_ _3803_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5872_ _4263_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8743__A1 as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7611_ _2799_ _2800_ _2805_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4823_ _4119_ _4404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5557__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9248__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8591_ as2650.psu\[4\] _3707_ _4465_ _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7542_ _1599_ _0890_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4754_ as2650.carry _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7473_ net34 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4685_ _4118_ _4265_ _4266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5626__I _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8002__I _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9212_ _0161_ clknet_leaf_41_wb_clk_i as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6424_ _1156_ _1375_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6355_ _1638_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9143_ _0092_ clknet_leaf_54_wb_clk_i as2650.stack\[0\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5306_ _0635_ _0552_ _0637_ _4454_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6809__A1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9074_ _0023_ clknet_leaf_46_wb_clk_i as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ _1488_ _1510_ _1570_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8158__B _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5237_ _0567_ _0451_ _0570_ _0470_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_103_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8025_ _4471_ _4483_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ _0439_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6037__A2 _4429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8431__B1 _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5099_ _0426_ _0429_ _0435_ _0412_ _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7785__A2 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6588__A3 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8927_ _4202_ _3994_ _1478_ _1463_ _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_25_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8858_ _1054_ _3941_ _3943_ _3944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7809_ _2991_ _4228_ _2992_ _2995_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5548__A1 _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5548__B2 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8789_ _3890_ _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8340__C _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8847__I _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7848__I0 _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6276__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5271__I as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7225__A1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7776__A2 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8973__A1 _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5787__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7528__A2 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5539__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6200__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8250__C _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5554__A4 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4762__A2 _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7661__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6140_ as2650.psu\[5\] _1409_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7464__A1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6071_ _4157_ _1353_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5022_ _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7216__A1 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8964__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5778__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6973_ _4243_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9070__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8712_ _3823_ _3833_ _3839_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ _1178_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7519__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8716__A1 _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8643_ _1376_ _2082_ _3789_ _0695_ _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5855_ as2650.stack\[1\]\[13\] _1142_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _4386_ _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8574_ _4508_ _3337_ _3723_ _3724_ _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5786_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8160__C _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7057__B _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7525_ _2153_ _2708_ _2721_ _2385_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4737_ _4317_ _4258_ _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5950__A1 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7456_ _2650_ _2652_ _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4668_ _4234_ _4180_ _4248_ _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_79_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6407_ _0692_ _1668_ _1681_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5702__A1 as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4599_ _4179_ _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7387_ _1631_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9126_ _0075_ clknet_leaf_0_wb_clk_i as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ _1619_ _1621_ _1578_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_88_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6269_ _0555_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9057_ _0006_ clknet_leaf_8_wb_clk_i as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8008_ _3174_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7207__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5481__A3 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7758__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8955__A1 _4466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8183__A2 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5266__I as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6497__A2 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7414__C _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7446__A1 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6249__A2 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8245__C _4497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8946__A1 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4680__A1 as2650.alu_op\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4983__A2 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8174__A2 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6185__A1 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5571_ _4357_ _4398_ _4336_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5932__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7310_ _2497_ _2510_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ _1112_ _2604_ _3451_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6488__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__B _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7241_ _2390_ _2441_ _2442_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_132_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7172_ _2309_ _2372_ _2375_ _2311_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7324__C _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5160__A2 _4476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7437__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ _1348_ _1352_ _1407_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_124_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7988__A2 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _0909_ _1196_ _1194_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_61_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5999__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5999__B2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5005_ as2650.r123\[1\]\[2\] as2650.r123\[0\]\[2\] as2650.r123_2\[1\]\[2\] as2650.r123_2\[0\]\[2\]
+ _4366_ _0339_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_113_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6660__A2 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7994__C _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6956_ _2168_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5907_ _1164_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6887_ as2650.stack\[4\]\[0\] _2109_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6176__A1 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8626_ _1583_ _2957_ _3773_ _3722_ _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5838_ _1139_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8557_ _1187_ _3297_ _3706_ _3708_ _3647_ _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5923__A1 _4347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _0699_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7508_ _2222_ _1572_ _2423_ _2704_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_8488_ _2362_ _4438_ _3642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7676__A1 _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7439_ _2402_ _2598_ _2637_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5814__I _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5151__A2 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9109_ _0058_ clknet_leaf_52_wb_clk_i as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7979__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6100__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8346__B _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7600__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4965__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8156__A2 _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9309__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5142__A2 _4452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7419__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8919__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6810_ _0715_ _1040_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7790_ _2724_ _2979_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__B1 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6741_ _1969_ _1970_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__A2 _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7386__I _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__I _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4803__I _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6672_ _1904_ _1901_ _1905_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8411_ _2856_ _3568_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5623_ _4478_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8342_ _2241_ _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5554_ _0356_ _0639_ _0661_ _0751_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_8273_ _3092_ _3427_ _3434_ _3435_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_117_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5485_ _0483_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5634__I as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7224_ _2403_ _2426_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6330__A1 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__A2 _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7155_ _2358_ _4438_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6106_ _1375_ _1377_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7086_ _2208_ _2286_ _2287_ _2289_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_115_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6037_ _1324_ _4429_ _1172_ _1233_ _0822_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_100_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7988_ _1350_ _1521_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6939_ _1511_ _2142_ _1671_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6149__A1 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8609_ as2650.psu\[5\] _3648_ _3758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7897__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7649__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7245__B _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__B2 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8855__I _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6872__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4883__A1 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8074__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8074__B2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6624__A2 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8377__A2 _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9131__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5060__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9281__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6560__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5270_ _4162_ _0551_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8765__I _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8065__A1 _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8960_ _1365_ _1390_ _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7911_ _3079_ _2935_ _3085_ _3086_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8891_ _3957_ _3968_ _3969_ _3970_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_64_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7842_ _3023_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6918__A3 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7773_ _2238_ _2958_ _2959_ _2962_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4985_ _4433_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5051__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6724_ _1914_ _1954_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7879__A1 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6655_ _1888_ _1891_ _1893_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6146__A4 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5606_ _4209_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5354__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _1827_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8325_ _0967_ _2605_ _3485_ _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5537_ _0868_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8256_ _3360_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6303__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5468_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6303__B2 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7207_ _2402_ _2404_ _2409_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8187_ _0554_ _0446_ _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5399_ _0536_ _0728_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7138_ _2337_ _2341_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7803__A1 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6606__A2 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9154__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8359__A2 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5967__C _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6909__A3 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5593__A2 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5896__A3 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8295__A1 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4856__A1 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8047__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8518__C _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8598__A2 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7929__I _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7022__A2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5449__I _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8770__A2 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5584__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _4249_ _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6440_ _4503_ _0984_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5336__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6533__B2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6371_ as2650.stack\[6\]\[10\] _1650_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8110_ _2440_ _4380_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8286__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5322_ _0657_ as2650.r123\[1\]\[5\] _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9090_ _0039_ clknet_leaf_50_wb_clk_i as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8041_ _3100_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5253_ _0584_ _0587_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5912__I _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4847__A1 _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9177__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5184_ _0515_ _4130_ _0518_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8589__A2 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4528__I _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7261__A2 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8943_ _3719_ _3001_ _4011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8874_ _3939_ _3955_ _3956_ _3953_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_36_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7013__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8210__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7825_ _1394_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8210__B2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7756_ _2933_ _2945_ _2946_ _2437_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5414__I3 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _0284_ _0298_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6707_ _1936_ _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7687_ _2768_ _2879_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4899_ _4476_ _4479_ _4480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _1882_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6569_ _1808_ _1811_ _1812_ _1805_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8277__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8308_ as2650.stack\[6\]\[7\] _3200_ _3202_ as2650.stack\[7\]\[7\] _0501_ _3470_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__8277__B2 _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9288_ _0237_ clknet_leaf_38_wb_clk_i as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8619__B _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7523__B _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8239_ _3401_ _3402_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8338__C _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8029__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8201__A1 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7004__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8201__B2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5110__S1 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5566__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8504__A2 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5318__A2 _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5869__A3 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8268__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A1 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8440__A1 _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _1159_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5006__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5006__B2 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7610_ _2802_ _2804_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4822_ _4111_ _4403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8590_ _1229_ _2957_ _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7541_ _2656_ _2659_ _2736_ _2714_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4753_ _4333_ _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7472_ _2368_ _2669_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4684_ _4251_ _4256_ _4264_ _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_105_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9211_ _0160_ clknet_leaf_6_wb_clk_i as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6423_ _4284_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8259__A1 _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9142_ _0091_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6354_ _1415_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5305_ _0638_ _0568_ _0640_ _0367_ _0317_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6809__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9073_ _0022_ clknet_leaf_45_wb_clk_i as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6285_ _1563_ _1569_ _1483_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8158__C _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8024_ _3189_ _3192_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7482__A2 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5236_ _0571_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6285__A3 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _0490_ _0499_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_96_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8431__A1 _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6037__A3 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8431__B2 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5098_ _4297_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_44_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8926_ _1155_ _3647_ _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6993__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8857_ _0368_ _3942_ _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7808_ _1352_ _1565_ _2992_ _2993_ _2994_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8788_ _0698_ _3888_ _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7739_ _2255_ _2262_ _2926_ _2929_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_33_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7848__I1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6276__A3 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8670__A1 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7225__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8084__B _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7479__I _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__A1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8489__A1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8259__B _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8661__A1 as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6070_ _1354_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input9_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ _4384_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7216__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9215__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4806__I _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8964__A2 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6972_ _2179_ _2159_ _2181_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8711_ as2650.stack\[4\]\[11\] _3836_ _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5923_ _4347_ _1192_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7519__A3 _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8716__A2 _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8642_ _1619_ _3720_ _3788_ _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6727__A1 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5854_ _1021_ _1144_ _1150_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8441__C _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4805_ net6 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8573_ _1376_ _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5785_ _1103_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6242__B _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5637__I _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7524_ _2466_ _2692_ _2720_ _2405_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8013__I _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4736_ _4316_ _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7455_ _2650_ _2652_ _2394_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7152__A1 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4667_ _4247_ _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ _1680_ _1672_ _1673_ _1678_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7386_ _2573_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5702__A2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _4172_ _4178_ _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9125_ _0074_ clknet_leaf_69_wb_clk_i as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6337_ _1620_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5305__C _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9056_ _0005_ clknet_leaf_8_wb_clk_i as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6268_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8007_ _1055_ _4197_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5219_ _0555_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6199_ _1429_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8616__C _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7207__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8404__A1 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8404__B2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8955__A2 _4499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8909_ as2650.stack\[2\]\[4\] _3982_ _3983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8707__A2 _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7391__A1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6194__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7930__A3 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4744__A3 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__A1 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8891__A1 _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8643__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5209__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4680__A2 as2650.alu_op\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8946__A2 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6957__A1 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7002__I _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5885__C _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7382__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ _0902_ _0354_ _4223_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7240_ _0350_ _0319_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8882__A1 _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6288__I _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7171_ _2373_ _2374_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _4391_ _1361_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7437__A2 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6053_ _0753_ _1272_ _1339_ _1233_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5004_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8937__A2 _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4671__A2 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ as2650.addr_buff\[2\] _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5906_ _4384_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6886_ _2107_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8625_ _1429_ _3720_ _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5837_ as2650.r123_2\[3\]\[7\] _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6176__A2 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8556_ as2650.psu\[2\] _3707_ _4465_ _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5768_ _1052_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7507_ _2690_ _2605_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _4146_ _4149_ _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8678__I _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8487_ _3640_ _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5699_ _1025_ _0974_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7438_ _2351_ _2630_ _2636_ _2497_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_107_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_100_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7369_ _2561_ _2565_ _2568_ _2466_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9108_ _0057_ clknet_leaf_50_wb_clk_i as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8625__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9039_ _3024_ _4096_ _1583_ _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7979__A3 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6926__I _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6100__A2 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6147__B _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8928__A2 _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6939__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__A2 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8400__I1 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7364__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__A2 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7492__I _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8313__B1 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9060__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7419__A2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8616__A1 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8092__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8919__A2 _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5602__B2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6740_ _1938_ _1946_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6671_ as2650.stack\[3\]\[5\] _1902_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7355__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8410_ _2815_ _3533_ _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5622_ _0942_ _0947_ _0953_ _4421_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_108_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8341_ _3063_ _3490_ _3499_ _3501_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__8498__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5553_ _4370_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5915__I _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8272_ _3128_ _3416_ _3418_ _2873_ _3191_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5484_ _0817_ _0791_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5669__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7223_ _1620_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5133__A3 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7154_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8607__A1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8447__B _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6105_ _1378_ _1380_ _1383_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5650__I _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7085_ _1523_ _1373_ _2288_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8166__C _4488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6036_ _4420_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9032__A1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7987_ _1390_ _2256_ _2474_ _2141_ _3155_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6938_ _2122_ _2152_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_41_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _2079_ _2089_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6149__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8608_ _1538_ _0792_ _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7526__B _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8539_ _1492_ _2956_ _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7649__A2 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__B1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4883__A2 _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6656__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4904__I _4484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6391__I _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5001__S _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5060__A2 _4510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7337__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5348__B1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7436__B _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6560__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4571__A1 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7950__I _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__A1 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9014__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7910_ _3080_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8890_ _3551_ _3970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7841_ _3022_ as2650.holding_reg\[5\] _3007_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7397__I _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7772_ _2960_ _2961_ _1378_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4984_ _4430_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6723_ _1915_ _1953_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7328__A1 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6654_ as2650.stack\[3\]\[0\] _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7879__A2 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6000__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5605_ _0293_ _0925_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6585_ _1831_ _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5645__I _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8324_ _2605_ _2767_ _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8021__I _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8828__A1 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ as2650.holding_reg\[7\] _4131_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8255_ _1621_ _2681_ _3417_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _0798_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7500__A1 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6303__A2 _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7206_ _2405_ _2407_ _2408_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8186_ _0676_ _0547_ _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ _0306_ _0722_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7081__B _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7137_ _2332_ _2340_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6476__I _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5380__I _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7068_ _4226_ _4504_ _0655_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_115_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8691__I _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6019_ _1234_ _1306_ _1307_ _1279_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__9005__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5290__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6542__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8819__A1 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8295__A2 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7770__I _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4856__A2 _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8047__A2 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7558__A1 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8106__I _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7010__I _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7022__A3 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7945__I as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6533__A2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__A1 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4544__A1 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _0990_ _1647_ _1651_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5321_ _4110_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7680__I _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8286__A2 _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8040_ _3198_ _3201_ _3208_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5252_ as2650.stack\[6\]\[11\] _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4847__A2 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__I _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5183_ _0519_ _4259_ _4323_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__A1 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8942_ _2588_ _4298_ _4009_ _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_3_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5272__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8873_ net44 _3945_ _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7824_ _1577_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7755_ net50 _2933_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4967_ _4338_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7855__I _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6706_ _1769_ _1038_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4783__A1 _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7686_ _2865_ _2878_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5980__B1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4898_ _4477_ as2650.stack\[5\]\[8\] as2650.stack\[4\]\[8\] _4478_ _4479_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8513__A3 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6637_ as2650.r123\[3\]\[2\] _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7721__A1 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7721__B2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6568_ _1829_ _1830_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8307_ _3327_ _3468_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5519_ _0584_ _0851_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9287_ _0236_ clknet_leaf_38_wb_clk_i as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6499_ _1763_ _1764_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8238_ _3127_ _3383_ _3394_ _2873_ _3190_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_106_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9121__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8169_ _3333_ _4475_ _3327_ _3334_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7788__A1 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7788__B2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9271__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8201__A2 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7960__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7712__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8268__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4541__A4 as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A2 _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4629__I _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7779__A1 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8440__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5254__A2 _4485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5006__A2 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4821_ _4385_ _4401_ _4402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7540_ _0900_ _0890_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4765__A1 _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4752_ _4332_ _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7471_ _2667_ _2664_ _2666_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4683_ _4133_ _4257_ _4260_ _4263_ _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__7703__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9210_ _0159_ clknet_leaf_3_wb_clk_i as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6422_ _4196_ _1673_ _1692_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9144__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9141_ _0090_ clknet_leaf_54_wb_clk_i as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8259__A2 _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6353_ _1636_ _1565_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ _0639_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9072_ _0021_ clknet_leaf_46_wb_clk_i as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6284_ _1564_ _1568_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8023_ _2311_ _3127_ _2873_ _3173_ _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__9294__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5235_ _0558_ _0517_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7482__A3 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5166_ _0492_ _0500_ _0503_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ _0430_ _0419_ _0421_ _4338_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__8174__C _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6442__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8925_ _1486_ _2198_ _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6993__A2 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8856_ _3940_ _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7807_ _1659_ _4271_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8190__B _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7585__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7942__A1 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8787_ _3888_ _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5999_ _1288_ _1205_ _1208_ _0673_ _1209_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4756__A1 _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7738_ _1657_ _1664_ _2917_ _2719_ _2928_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7669_ _2135_ _2860_ _2861_ _2127_ _2172_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5484__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6681__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8422__A2 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5236__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8973__A3 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8186__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7933__A1 _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A1 _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9167__CLK clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8489__A2 _4459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5172__A1 _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5743__I _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8110__A1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8661__A2 _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6672__A1 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5475__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5020_ _0355_ _0356_ _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6424__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6971_ _2180_ _2174_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8710_ _3821_ _3833_ _3838_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _4459_ _1193_ _1215_ _1192_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8177__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ as2650.stack\[1\]\[12\] _1146_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8641_ as2650.psu\[7\] _3648_ _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5918__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4822__I _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ _4373_ _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5784_ as2650.pc\[6\] _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8572_ _1588_ _2957_ _3721_ _3722_ _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7523_ _2713_ _2718_ _2719_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4735_ _4299_ _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7454_ _2622_ _2626_ _2651_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_135_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _4242_ _4246_ _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6405_ _0353_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6749__I _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7385_ _2576_ _2579_ _2584_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5653__I _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4597_ _4113_ _4177_ _4178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6336_ _1336_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9124_ _0073_ clknet_leaf_69_wb_clk_i as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8101__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9055_ _0004_ clknet_leaf_9_wb_clk_i as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _0456_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5218_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8006_ _1682_ _3173_ _3174_ _1456_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6198_ _1432_ _1440_ _1444_ _1482_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_85_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8404__A2 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ _0478_ _0486_ _0410_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8908_ _3974_ _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8168__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8632__C _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8168__B2 _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8839_ _0690_ _3927_ _3928_ as2650.r123\[2\]\[4\] _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8204__I _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7391__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7930__A4 _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7143__A2 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8340__A1 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6659__I _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8891__A2 _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8643__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5457__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5209__A2 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6406__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6957__A2 _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8159__A1 _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7439__B _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6709__A2 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7906__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5738__I _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7382__A2 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5393__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6590__B1 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8331__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7174__B _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8882__A2 _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7170_ _2308_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6121_ _1358_ _1393_ _1406_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6052_ _1198_ _1338_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5003_ as2650.r0\[2\] _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__I _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8398__A1 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9332__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7070__A1 _4514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _1609_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__A2 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5905_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6885_ _2107_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4552__I _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8624_ _3705_ _1040_ _3652_ _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5836_ _1138_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8570__A1 _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5384__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5767_ _1053_ _1087_ _1088_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8555_ _1400_ _1348_ _1403_ _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7506_ _2698_ _2702_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4718_ as2650.r0\[0\] _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5698_ as2650.pc\[13\] _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8486_ _2207_ _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__A1 _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7437_ _2389_ _2634_ _2635_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4649_ _4224_ _4180_ _4229_ _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _2566_ _2567_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9107_ _0056_ clknet_leaf_7_wb_clk_i as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6319_ _4335_ _4386_ _0757_ _1602_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7299_ _1609_ _0479_ _0484_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_104_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8627__C _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9038_ _4091_ _4092_ _4096_ _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7103__I _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8928__A3 _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6939__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7061__A1 _4126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5558__I _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6163__B _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7364__A2 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8869__I _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5494__S _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8313__A1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8313__B2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5127__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9205__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8616__A2 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7441__C _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7052__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8272__C _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5602__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6670_ _1099_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5621_ _0948_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5366__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8340_ _3097_ _3481_ _3500_ _3092_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5552_ _0817_ _0791_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7616__C _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8304__A1 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8271_ _3066_ _3415_ _3433_ _2935_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6299__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5483_ _0669_ _0660_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6866__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7222_ _2424_ _2406_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7632__B _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7153_ _4246_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8607__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5931__I _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ _1388_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7084_ _4115_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4547__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6035_ _1199_ _1321_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9032__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7858__I _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7986_ _2251_ _2271_ _2921_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6937_ _2121_ _2123_ _1460_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_74_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6868_ _1332_ _2072_ _2073_ as2650.r123_2\[2\]\[6\] _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7346__A2 _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8543__A1 _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8607_ _2779_ _0736_ _3640_ _3755_ _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5357__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5819_ as2650.stack\[0\]\[6\] _1127_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6799_ _1998_ _2018_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7526__C _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8538_ _3646_ _0984_ _1519_ _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__A1 _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8469_ _1030_ _3623_ _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6857__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8638__B _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5841__I _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6609__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7282__A1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8782__A1 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5596__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7337__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5348__B2 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4571__A2 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7008__I _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6848__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8548__B _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5751__I _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6076__A2 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9014__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7840_ _2179_ _1624_ _3021_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8773__A1 _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7771_ _2314_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _0314_ _0320_ _0321_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ _1918_ _1952_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7328__A2 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8525__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6653_ _1890_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5604_ _4426_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6584_ _1832_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8323_ _3480_ _3483_ _2298_ _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5535_ _4359_ _4277_ _0867_ _4163_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8254_ _1103_ _3171_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5466_ _0799_ _0795_ _0796_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7500__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7205_ _2310_ _1550_ _2406_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_8185_ _2144_ _3349_ _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5397_ _4341_ _0730_ _0731_ _0431_ _0433_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_67_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7136_ _2206_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7067_ _2270_ _2233_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _0783_ _1196_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9005__A2 _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5610__B _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__A2 _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8764__A1 _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7969_ _3004_ _3139_ _2748_ _3126_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8516__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_33_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_33_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6667__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8087__C _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7498__I _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7007__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7558__A2 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8323__S _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8507__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4792__A2 _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7730__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4544__A2 _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5320_ _4403_ as2650.r123_2\[1\]\[5\] _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7494__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ _4475_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _0444_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7246__A1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8792__I _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8994__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8941_ _0620_ _4007_ _4008_ _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9073__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8872_ _0598_ _3941_ _3954_ _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8746__A1 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7823_ _3008_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6221__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7754_ _1677_ _2937_ _2938_ _2944_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4966_ _0299_ _0303_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_71_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6705_ _1734_ _1835_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7685_ _2830_ _2877_ _2866_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4783__A2 _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__B2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _4468_ _4478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6636_ _1881_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8513__A4 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6567_ _0611_ _1005_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8306_ _0386_ as2650.stack\[5\]\[7\] as2650.stack\[4\]\[7\] _0383_ _3468_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_105_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5518_ _4494_ as2650.stack\[3\]\[14\] as2650.stack\[2\]\[14\] _4473_ _4498_ _0852_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_9286_ _0235_ clknet_leaf_49_wb_clk_i as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6498_ _1297_ _1697_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7485__A1 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__B _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8237_ _3233_ _3383_ _3400_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5449_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8168_ _0383_ as2650.stack\[5\]\[3\] as2650.stack\[4\]\[3\] _3328_ _3334_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7119_ _0902_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8434__B1 _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8099_ _3037_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6460__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4735__I _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7111__I _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8737__A1 _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7960__A2 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5971__A1 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7712__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8877__I _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7781__I _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7714__C _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7476__A1 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9096__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7228__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__B _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7779__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8976__A1 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8545__C _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6451__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4645__I _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7956__I _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7400__A1 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _4387_ _4396_ _4400_ _4401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _4309_ _4293_ _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7470_ _2664_ _2666_ _2667_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4682_ _4262_ _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8900__A1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6421_ _1691_ _1684_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9140_ _0089_ clknet_leaf_53_wb_clk_i as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6352_ _0827_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7467__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ _4383_ _0458_ _0516_ _0608_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_9071_ _0020_ clknet_leaf_45_wb_clk_i as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6283_ _1566_ _1567_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8022_ _3190_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _4434_ _4244_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7219__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5165_ _4494_ as2650.stack\[3\]\[10\] as2650.stack\[2\]\[10\] _4476_ _0502_ _0503_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_68_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8967__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5096_ _0431_ _0432_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_56_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6442__A2 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8027__I _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8924_ _1435_ _2270_ _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6993__A3 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8855_ _3940_ _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7806_ _0926_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8786_ _3880_ _3887_ _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _0675_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4756__A2 _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5953__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7737_ _2243_ _2927_ _2292_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4949_ as2650.holding_reg\[1\] _4129_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7668_ _2741_ _2821_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6619_ _0977_ _1870_ _1872_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8697__I _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7599_ _2780_ _2793_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5181__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7458__A1 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5335__B _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9269_ _0218_ clknet_leaf_50_wb_clk_i as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8365__C _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4692__A1 as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8958__A1 _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4995__A2 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8186__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7709__C _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7933__A2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8110__A2 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8556__B _4465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4683__A1 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8949__A1 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6970_ _4244_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _4438_ _1195_ _1193_ _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_46_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8177__A2 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8640_ _3722_ _3474_ _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ _1012_ _1143_ _1149_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6188__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9111__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ _4383_ _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8571_ _4506_ _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5783_ _0823_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7522_ _2497_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4734_ _4314_ _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7688__A1 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7453_ _0756_ _0741_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4665_ as2650.addr_buff\[7\] _4245_ _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__9261__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _4148_ _1668_ _1679_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7384_ _2566_ _2324_ _2329_ _2583_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4596_ _4176_ _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9123_ _0072_ clknet_leaf_68_wb_clk_i as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6335_ _1608_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4910__A2 _4485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8101__A2 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9054_ _0003_ clknet_leaf_9_wb_clk_i as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6266_ _0353_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _1057_ _0938_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5217_ net9 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6663__A2 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5466__A3 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4674__A1 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6197_ _1464_ _1481_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ _4449_ _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5079_ _0413_ _0415_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_44_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8907_ _3974_ _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8838_ _3916_ _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6974__I0 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8769_ _3821_ _3870_ _3875_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7679__A1 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8340__A2 _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6351__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4901__A2 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6103__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8376__B _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6654__A2 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7851__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8095__C _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4665__A1 as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8890__I _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7603__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9134__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7906__A2 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5917__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9284__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6590__A1 as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7455__B _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8331__A2 _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6342__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6893__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8095__A1 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ _1395_ _1363_ _1399_ _1405_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7190__B _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6051_ _0904_ _1209_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _4361_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_85_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7070__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6953_ _1236_ _2159_ _2166_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__I as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5081__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4833__I _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5904_ _4441_ _1197_ _4221_ _4214_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_81_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6884_ _1045_ _1854_ _1118_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_74_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8623_ _3079_ _0814_ _2208_ _3770_ _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5835_ as2650.r123_2\[3\]\[6\] _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8554_ as2650.overflow _3648_ _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5766_ as2650.stack\[1\]\[3\] _1063_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7505_ _2699_ _2701_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4717_ _4297_ _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5664__I _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8485_ _2779_ _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5697_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8322__A2 _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7436_ _1585_ _4447_ _2126_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5136__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4648_ _4225_ _4227_ _4228_ _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_107_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7367_ _2523_ _2494_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4579_ _4159_ _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9106_ _0055_ clknet_leaf_11_wb_clk_i as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ as2650.psl\[5\] _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7298_ _0479_ _0484_ _1609_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_104_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9037_ _4093_ _4095_ _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6249_ _1528_ _1533_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4647__A1 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9157__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_58_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_58_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7061__A2 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A1 _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8010__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5375__A2 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8313__A2 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5523__B _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6627__A2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4918__I _4498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A1 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5686__I0 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7052__A2 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5063__A1 _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4653__I _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8001__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8552__A2 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5620_ _0293_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8270_ _2677_ _3431_ _3432_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5482_ _0815_ _0791_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7221_ _1055_ net6 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6866__A2 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4877__A1 _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8068__A1 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7152_ _1549_ _2355_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ _0922_ _4181_ _4294_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_119_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7083_ _4234_ _1459_ _0939_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_112_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6248__C _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _0664_ _1272_ _1160_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7579__B1 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8240__A1 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7043__A2 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8240__B2 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7985_ _1523_ _3151_ _3153_ _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5659__I _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _1188_ _2150_ _0950_ _4421_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6867_ _2075_ _2092_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8543__A2 _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8606_ _2557_ _3753_ _3754_ _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5818_ _1100_ _1126_ _1129_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5357__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6798_ _2001_ _2017_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8537_ _0348_ _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5749_ _1053_ _1071_ _1072_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8468_ _1025_ _3606_ _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7419_ _1096_ _0755_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_124_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8399_ _2173_ _3556_ _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_2_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__A1 _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8059__A1 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4738__I _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7282__A2 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8231__A1 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5569__I _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8782__A2 _4464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6793__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8534__A2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6545__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8298__A1 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4571__A3 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9322__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7733__B _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8548__C _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5284__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8222__A1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8773__A2 _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7770_ _0924_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6784__A1 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _4289_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6721_ _1922_ _1951_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7694__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_3_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8525__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _1890_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6536__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7879__A4 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _4255_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6583_ _1838_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8322_ _0967_ _3482_ _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8289__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ _4276_ _0825_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8253_ _3415_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _0790_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7204_ _1055_ _4386_ _2406_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8184_ _1288_ _0407_ _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5511__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _0729_ _0720_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7135_ _2338_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6974__S _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4558__I as2650.alu_op\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8461__A1 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7066_ _4227_ _4199_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7869__I _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _0742_ _1235_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5610__C _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8764__A2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7968_ _2361_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _4425_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7899_ _1632_ _3061_ _3075_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8516__A2 _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7109__I _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5057__C _4489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7553__B _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6948__I _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5502__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8452__A1 _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7007__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8507__A2 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6351__C _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__A3 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7019__I _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5762__I _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7494__A2 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5250_ _0585_ as2650.stack\[5\]\[11\] as2650.stack\[4\]\[11\] _0586_ _0587_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5181_ _4275_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8443__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9218__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8940_ _0879_ _0875_ _0872_ _0536_ _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8871_ _0681_ _3942_ _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7822_ _3006_ as2650.holding_reg\[1\] _3007_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7753_ _2940_ _2943_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6221__A3 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4965_ _0299_ _0303_ _4333_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5937__I _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6704_ _1933_ _1934_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7684_ _2845_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5980__A2 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4896_ as2650.psu\[1\] _4477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6635_ as2650.r123\[3\]\[1\] _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6566_ _1770_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8305_ _3138_ _3449_ _3452_ _2586_ _2839_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_106_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5517_ _0592_ as2650.stack\[1\]\[14\] as2650.stack\[0\]\[14\] _0586_ _0851_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9285_ _0234_ clknet_leaf_36_wb_clk_i as2650.stack\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8131__B1 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6497_ as2650.r123_2\[1\]\[4\] _1699_ _1762_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8236_ _3384_ _3390_ _3399_ _2934_ _3091_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7485__A2 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5448_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8167_ as2650.stack\[6\]\[3\] _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5379_ _0712_ _0662_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7118_ _2321_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8434__A1 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8434__B2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8098_ _1075_ _3264_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7049_ _1400_ _4158_ _1353_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5799__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6996__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8198__B1 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6008__I _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5971__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7476__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7228__A2 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8425__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7779__A3 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4926__I _4506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6987__A1 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8728__A2 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7400__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8133__I _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _4315_ _4330_ _4331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4681_ _4134_ _4261_ _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6420_ _1545_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8900__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6911__A1 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _1166_ _0883_ _1507_ _1634_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5492__I _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5302_ _0609_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9070_ _0019_ clknet_leaf_45_wb_clk_i as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6282_ _1531_ _1470_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5478__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8021_ _0940_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5233_ _0568_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_130_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7219__A2 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8416__A1 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5164_ _0501_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8967__A2 _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ _4292_ _4293_ _4295_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_84_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8923_ _1189_ _0696_ _3990_ _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8719__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8854_ _1572_ _4245_ _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7805_ _2259_ _2261_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8785_ _3886_ _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5667__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5997_ _4442_ _1230_ _1252_ _4279_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7736_ _2281_ _2284_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4948_ _0286_ _4273_ _4319_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5953__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7667_ _2730_ _2732_ _2821_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7155__A1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _4449_ _4459_ _4460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5005__I1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6618_ as2650.stack\[0\]\[8\] _1871_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7598_ _2185_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6902__A1 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8199__B _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6549_ _1805_ _1812_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5108__S _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7458__A2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9268_ _0217_ clknet_leaf_36_wb_clk_i as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8219_ _1097_ _3381_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9199_ _0148_ clknet_leaf_26_wb_clk_i net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8646__C _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8407__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4692__A2 as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5641__A1 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6961__I _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7933__A3 _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7792__I _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8343__B1 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8894__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9063__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6201__I _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8646__A1 _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4683__A2 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5880__A1 _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7967__I _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5632__A1 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5920_ _4354_ _1196_ _1194_ _1213_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ as2650.stack\[1\]\[11\] _1146_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5487__I _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6188__A2 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ _4378_ _4382_ _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8570_ _4357_ _3720_ _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5782_ _1089_ _1100_ _1101_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7521_ _2498_ _2716_ _2717_ _2353_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8798__I _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4733_ as2650.psl\[3\] as2650.carry _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7137__A1 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7452_ _2649_ _0840_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8885__A1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4664_ _4243_ _4244_ _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5699__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6403_ _1669_ _1672_ _1673_ _1678_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7383_ _2321_ _2582_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4595_ _4175_ _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9122_ _0071_ clknet_leaf_68_wb_clk_i as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6334_ _1615_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9053_ _0002_ clknet_leaf_9_wb_clk_i as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _1549_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8004_ _1544_ _2325_ _3172_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5216_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6196_ _1466_ _1467_ _1472_ _0335_ _1480_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4566__I _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5147_ _0479_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ as2650.holding_reg\[2\] _4323_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5623__A1 _4478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8906_ _3975_ _1087_ _3980_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8837_ _3914_ _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7376__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6179__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8768_ as2650.stack\[7\]\[10\] _3873_ _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6974__I1 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7719_ _2793_ _2910_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8699_ _3829_ _3816_ _3830_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7679__A2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7117__I _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6351__A2 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8628__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8628__B2 _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6956__I _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7300__A1 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6103__A2 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6177__B _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4665__A2 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5862__A1 _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7603__A2 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8800__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A1 _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8564__B1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5100__I _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8867__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6342__A2 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8619__A1 _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8095__A2 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5770__I as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _1336_ _1237_ _1207_ _0898_ _1164_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input7_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A2 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9044__A1 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5605__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _2165_ _2163_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__A2 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5903_ _4166_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7358__A1 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6883_ _1346_ _2102_ _2105_ _1298_ _2106_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_34_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8622_ _3701_ _0821_ _2385_ _3769_ _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5834_ _1137_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5010__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6030__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5765_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8553_ _3646_ _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7504_ _2700_ _2680_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4716_ _4296_ _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8858__A1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8484_ _2436_ _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5696_ _0649_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7435_ _0757_ _0771_ _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _4155_ _4134_ _4143_ _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7530__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7366_ net32 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4578_ as2650.ins_reg\[2\] as2650.ins_reg\[3\] _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6317_ _1593_ _1594_ _1598_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_9105_ _0054_ clknet_leaf_41_wb_clk_i as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7297_ _4278_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9036_ _4078_ _4094_ _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7833__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ _0793_ _1401_ _1532_ _1419_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4647__A2 _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9035__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6179_ _1449_ _1453_ _1457_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_131_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_opt_3_0_wb_clk_i_I clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7061__A3 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7349__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__A1 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_27_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8849__A1 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8849__B2 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5590__I _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6088__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5686__I1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9026__A1 _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7588__A1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9251__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5063__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4810__A2 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5765__I _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7760__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _0866_ _0882_ _0311_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5481_ _0357_ _0639_ _0661_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_144_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7512__A1 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7220_ _2422_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7151_ _4447_ _4459_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8068__A2 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6079__A1 _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7815__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7082_ _1252_ _2279_ _2280_ _2285_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9017__A1 _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6033_ _0826_ _1201_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7579__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7579__B2 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7984_ _1511_ _3152_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6251__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _0948_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6866_ _1703_ _2091_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7376__B _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8605_ _2648_ _0771_ _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5817_ as2650.stack\[0\]\[5\] _1127_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6797_ _1993_ _2020_ _2024_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7751__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6554__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5748_ as2650.stack\[1\]\[1\] _1063_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8536_ _1396_ _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7503__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5679_ as2650.pc\[11\] _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8467_ _3128_ _3620_ _3621_ _3191_ _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7418_ _2366_ _2152_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__9124__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8398_ _2169_ _3537_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4868__A2 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8059__A2 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7349_ _1558_ _2387_ _2354_ _2548_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9274__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9019_ _3018_ _4080_ _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__A2 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8231__A2 _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7130__I _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8782__A3 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7990__A1 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5596__A3 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5585__I _4477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5518__C _4498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8298__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9006__B _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8470__A2 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5284__A2 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8564__C _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8136__I _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8222__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6233__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4981_ _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6720_ _1924_ _1950_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_44_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6651_ _1889_ _1047_ _1051_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7733__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5602_ _0925_ _0929_ _0932_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6582_ _1841_ _1844_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8321_ _2689_ _3456_ _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5533_ _4226_ _0826_ _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8252_ _1105_ _3414_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5464_ _0790_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7203_ as2650.pc\[1\] net7 _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9297__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4839__I _4182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8183_ _2541_ _3308_ _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5395_ _0729_ _0720_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7215__I _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7134_ _4256_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7065_ _2233_ _2234_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6016_ _0754_ _1201_ _1199_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8213__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7967_ _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7972__A1 _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7972__B2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _1486_ _2127_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7898_ _3063_ _3072_ _3074_ _2588_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_126_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8516__A3 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7724__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6849_ _1312_ _2072_ _2073_ as2650.r123_2\[2\]\[5\] _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8519_ _1197_ _3672_ _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8649__C _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7125__I _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4710__A1 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8384__C _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_42_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_42_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7963__A1 _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__B1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7715__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6518__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8140__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5264__B _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7494__A3 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_6__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5180_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6454__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5257__A2 _4476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8870_ _3939_ _3951_ _3952_ _3953_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_64_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6206__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7821_ _2996_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_64_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7752_ net50 _2941_ _2308_ _2942_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ _4336_ _0301_ _0302_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6703_ _1838_ _1845_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7706__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7683_ _2872_ _2875_ _2772_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6509__A2 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4895_ _4475_ _4476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6114__I _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6634_ _1880_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5193__A1 _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6565_ _1701_ _1803_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8304_ _3092_ _3465_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5516_ _4499_ _0846_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6496_ _1298_ _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9284_ _0233_ clknet_leaf_50_wb_clk_i as2650.stack\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8131__A1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8131__B2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8235_ _2299_ _3392_ _3395_ _3398_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5447_ _0716_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8166_ _0919_ as2650.stack\[3\]\[3\] as2650.stack\[2\]\[3\] _3331_ _4488_ _3332_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5378_ as2650.holding_reg\[5\] _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7117_ _2320_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8434__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8097_ _1067_ _3176_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7048_ _4185_ _1519_ _2224_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6996__A2 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8198__A1 _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9312__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8198__B2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8999_ _3718_ _4062_ _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4759__A1 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8370__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6959__I _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5184__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7283__C _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8122__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8122__B2 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7228__A3 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8425__A2 _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6436__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5239__A2 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__A2 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5103__I _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7936__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5411__A2 _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ as2650.alu_op\[1\] as2650.alu_op\[2\] _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8361__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5773__I _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6911__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6350_ _1633_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5301_ _0609_ _0636_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6281_ _0827_ _0887_ _1565_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5478__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8020_ _2970_ _3184_ _3188_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5232_ _0459_ _0471_ _0557_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6675__A1 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5163_ _4496_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8416__A2 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8967__A3 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5094_ _0418_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8922_ _2601_ _1412_ _1432_ _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5013__I _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8853_ _3938_ _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7927__A1 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7804_ _1351_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8784_ _1695_ _3885_ _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _1180_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5402__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7735_ _1032_ _1375_ _2257_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _4379_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7666_ _2857_ _2858_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7155__A2 _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4878_ _4458_ _4459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7384__B _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6617_ _1869_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5166__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__I _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7597_ _2789_ _2791_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_101_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6548_ _1808_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8104__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8104__B2 _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8655__A2 _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9267_ _0216_ clknet_leaf_38_wb_clk_i as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6479_ _1744_ _1745_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8218_ _2594_ _3381_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9198_ _0147_ clknet_leaf_26_wb_clk_i net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8149_ _3171_ _2522_ _3314_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7091__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A2 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8591__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8343__A1 _4501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8343__B2 _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9208__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8646__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4683__A3 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7082__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5632__A2 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5768__I _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ _1001_ _1143_ _1148_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4801_ _4381_ _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5396__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5781_ as2650.stack\[1\]\[5\] _1094_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7520_ _2320_ _2498_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4732_ _4311_ _4312_ _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7137__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8334__A1 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5148__A1 _4449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7451_ _0830_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4663_ as2650.addr_buff\[5\] _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5699__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _1671_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7382_ _2558_ _2581_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4594_ _4174_ _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_122_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9121_ _0070_ clknet_leaf_68_wb_clk_i as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6333_ _1608_ _1616_ _1367_ _1382_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8637__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5008__I _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _4387_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9052_ _0001_ clknet_leaf_9_wb_clk_i as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8003_ _1057_ _3171_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5452__B _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5215_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5320__A1 _4403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _1422_ _1377_ _1474_ _1479_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7223__I _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ _0481_ _0459_ _0482_ _0483_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7073__A1 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _0414_ _4275_ _4320_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5623__A2 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8905_ as2650.stack\[2\]\[3\] _3976_ _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__I _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8836_ _3925_ _3926_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7376__A2 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6179__A3 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8767_ _3818_ _3870_ _3874_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ _0480_ _0572_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7718_ _2891_ _2909_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8698_ as2650.stack\[5\]\[14\] _3814_ _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7649_ _0998_ _2574_ _2840_ _2842_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9319_ _0268_ clknet_leaf_44_wb_clk_i as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8628__A2 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6103__A3 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5311__A1 _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4757__I _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7133__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5862__A2 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8800__A2 _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6811__A1 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5614__A2 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6193__B _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8564__A1 _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8564__B2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5378__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8316__A1 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6327__B1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9180__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7752__B _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4667__I _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5000_ _4375_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6951_ as2650.addr_buff\[1\] _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5498__I _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5902_ _1160_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6882_ as2650.r123_2\[2\]\[7\] _2073_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7358__A2 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8555__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8621_ _2399_ _0841_ _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5833_ as2650.r123_2\[3\]\[5\] _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7927__B _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8602__I _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8552_ _3639_ _0437_ _3641_ _3703_ _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8307__A1 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5764_ _0598_ _1081_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6581__A3 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7503_ as2650.pc\[6\] net2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4715_ _4292_ _4293_ _4295_ _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8483_ _3123_ _3637_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5695_ _0978_ _1021_ _1022_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7434_ _2544_ _2631_ _2545_ _2632_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4646_ _4226_ _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6333__A3 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5541__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7365_ _2563_ _2564_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4577_ _4154_ _4157_ _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9104_ _0053_ clknet_leaf_10_wb_clk_i as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6316_ _4387_ _0367_ _0441_ _0351_ _0826_ _1599_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7296_ _2121_ _2366_ _2123_ _1460_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7294__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6097__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9035_ _2199_ _1695_ _1468_ _4167_ _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_89_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6247_ _1401_ _1531_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4647__A3 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9035__A2 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6178_ _1462_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_40_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7046__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8243__B1 as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _4414_ _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7841__I0 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9053__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A3 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8546__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8940__C _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8819_ _3912_ _3886_ _3913_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_opt_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__A2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8849__A2 _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__B1 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_67_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_67_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5532__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8387__C _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6088__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7588__A2 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9011__C _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7747__B _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4810__A3 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7760__A2 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5480_ _0805_ _0810_ _0813_ _0790_ _4298_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__7512__A2 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7482__B _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7150_ _2353_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7276__A1 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6079__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6101_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7081_ _2281_ _2284_ _2132_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _0833_ _1238_ _1208_ _0829_ _1165_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9017__A2 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7579__A2 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8776__A1 as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7983_ _2143_ _2473_ _2191_ _0923_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6251__A2 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6934_ _0945_ _2147_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8528__A1 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _2079_ _2089_ _2090_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_62_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8604_ _2399_ _0741_ _3753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4860__I _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _1093_ _1126_ _1128_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6796_ _1995_ _2019_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7751__A2 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8535_ _1514_ _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5747_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8466_ _1030_ _2768_ _2573_ _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5678_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7503__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7392__B _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7417_ _1097_ _2419_ _2614_ _2615_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5514__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _4209_ _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8397_ _3554_ _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__A3 _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7348_ _2387_ _2547_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7267__A1 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7279_ _2424_ _2480_ _2460_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5817__A2 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9018_ _3043_ _4076_ _4079_ _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_89_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8767__A1 _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6242__A2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8519__A1 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5596__A4 _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7567__B _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__I _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7742__A2 _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5087__B _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9006__C _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9099__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7258__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5106__I _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8470__A3 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8207__B1 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8758__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__A2 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _0315_ _0316_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5441__B1 _4484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8580__C _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7981__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5992__A1 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6650_ _0917_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8930__A1 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7733__A2 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5601_ net3 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6581_ _1806_ _1842_ _1843_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_31_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8320_ _3480_ _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5532_ as2650.holding_reg\[7\] _4163_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8251_ _2594_ _3381_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5463_ _0795_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7202_ _2367_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6400__I _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5444__C _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8182_ _3233_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5394_ _0714_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7249__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7133_ net54 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7940__B _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8997__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7064_ _2266_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6015_ _0758_ _1238_ _1303_ _1255_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7966_ _1475_ _1350_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7972__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6917_ _0928_ _2130_ _2131_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_70_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5983__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7897_ _2223_ _3067_ _3073_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_39_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8516__A4 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6848_ _1298_ _2071_ _2074_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7724__A2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8921__A1 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5735__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _2006_ _2007_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6932__B1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8518_ _1154_ _1433_ _3671_ _4203_ _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7488__A1 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8449_ _3138_ _3600_ _3604_ _2572_ _2838_ _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7406__I _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6160__A1 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7850__B _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4710__A2 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5370__B _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7660__A1 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A2 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7963__A2 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7715__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_11_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8140__A2 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4701__A2 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8979__A1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4675__I _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7651__A1 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6454__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8591__B _4465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7403__A1 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7820_ _3003_ _3004_ _3005_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7751_ _1416_ _2264_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4963_ _0300_ _4321_ _4324_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5965__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6702_ _1841_ _1844_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7682_ _1008_ _2873_ _2874_ _2838_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4894_ _4471_ _4475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ as2650.r123\[3\]\[0\] _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9264__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6564_ _1802_ _1813_ _1814_ _1800_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6390__A1 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8303_ _3233_ _3450_ _3458_ _3069_ _3464_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5515_ as2650.stack\[6\]\[14\] _0588_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9283_ _0232_ clknet_leaf_36_wb_clk_i as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6495_ _1746_ _1760_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8131__A2 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6130__I _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8234_ _2418_ _3382_ _3397_ _1419_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ _0777_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7890__A1 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8165_ _0377_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5377_ _0422_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7116_ _1543_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8096_ _2299_ _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7642__A1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7047_ _4224_ _4169_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6996__A3 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8198__A2 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8998_ _3762_ _4061_ _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7949_ _1427_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4759__A2 _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6305__I as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5708__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8370__A2 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7136__I _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7633__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6436__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9137__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7936__A2 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A1 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9287__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8361__A2 _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6372__A1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _0558_ _0517_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6280_ _1468_ _1469_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6885__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7872__A1 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5231_ _0357_ _0316_ _0346_ _0450_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_102_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4686__A1 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ _0495_ as2650.stack\[1\]\[10\] as2650.stack\[0\]\[10\] _0496_ _0500_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5093_ _4342_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8967__A4 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8921_ _1513_ _2120_ _2991_ _1576_ _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_49_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8852_ _2213_ _2920_ _3670_ _3937_ _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_92_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7803_ _2986_ _2989_ _2990_ _2982_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8975__I1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5938__A1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8783_ _3883_ _4205_ _4430_ _3884_ _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ as2650.r123_2\[0\]\[4\] _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6125__I _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7734_ _2238_ _2920_ _2921_ _2924_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4946_ _4273_ _4377_ _4381_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4610__A1 _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7665_ _2816_ _2817_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4877_ _4450_ _4457_ _4458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5005__I3 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6616_ _1869_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7596_ _2790_ _2765_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6547_ _1779_ _1809_ _1810_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_134_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8104__A2 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6115__A1 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9266_ _0215_ clknet_leaf_37_wb_clk_i as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6478_ _1283_ _1705_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8496__B _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8217_ _1091_ _1082_ _3305_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7863__A1 _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5429_ _0758_ _0354_ _0763_ _4374_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_9197_ _0146_ clknet_leaf_27_wb_clk_i net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4677__A1 as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8148_ _1083_ _0902_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7615__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8079_ _3244_ _4471_ _3195_ _3246_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A3 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7379__B1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8591__A2 _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7575__B _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8343__A2 _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6106__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6657__A2 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A1 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7606__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4683__A4 _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5114__I _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7082__A2 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4800_ _4379_ _4174_ _4300_ _4380_ _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8582__A2 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5780_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6593__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7485__B _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _4139_ _4196_ _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5784__I as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7450_ _2629_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4662_ as2650.addr_buff\[6\] _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5148__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6345__A1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6401_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7381_ _2580_ _2521_ _2513_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _4173_ as2650.ins_reg\[1\] _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9120_ _0069_ clknet_3_2__leaf_wb_clk_i as2650.alu_op\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8098__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6332_ _0901_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9302__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9051_ _0000_ clknet_leaf_9_wb_clk_i as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7845__A1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6263_ _4392_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4659__A1 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8002_ _0901_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5214_ _0546_ _0548_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_69_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5320__A2 as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6194_ _1477_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5145_ _0480_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5024__I _4373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8270__A1 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7073__A2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5076_ _0343_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4863__I _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8904_ _3975_ _1079_ _3979_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4831__A1 _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8835_ _2049_ _3919_ _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6179__A4 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8766_ as2650.stack\[7\]\[9\] _3873_ _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5978_ _0597_ _1223_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7717_ _2908_ _2887_ _2889_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4929_ _4509_ _4510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8697_ _1042_ _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8325__A2 _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7648_ net52 _2472_ _2577_ _2169_ _2841_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5139__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6887__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7579_ _0968_ _2727_ _2774_ _2536_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_101_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__A1 _4477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8089__A1 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9318_ _0267_ clknet_leaf_44_wb_clk_i as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4898__B2 _4478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7836__A1 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9249_ _0198_ clknet_leaf_43_wb_clk_i as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7064__A2 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4773__I _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A3 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7289__C _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8564__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8316__A2 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__A1 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9325__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__B2 _4403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7752__C _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7827__A1 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8252__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6950_ _2120_ _2159_ _2164_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4813__A1 _4389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8004__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5901_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6881_ _2103_ _2098_ _2104_ _2084_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_81_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8555__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8620_ _0651_ _3683_ _3768_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5832_ _1136_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5369__A2 _4473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8551_ _3701_ _0476_ _2557_ _3702_ _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _1084_ _1059_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7502_ _1103_ _1595_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4714_ _4154_ _4294_ _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8482_ _1030_ _3528_ _3636_ _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5694_ as2650.stack\[2\]\[12\] _0991_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7433_ _2623_ _0642_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4645_ _4163_ _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6333__A4 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7364_ _2558_ _2560_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4576_ _4137_ _4156_ _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9103_ _0052_ clknet_leaf_10_wb_clk_i as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6315_ net3 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7295_ _2365_ _2495_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7234__I _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9034_ _3009_ _4515_ _1405_ _2300_ _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6246_ _1529_ _1530_ _0860_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8491__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ _1458_ _1372_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9035__A3 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8243__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _4374_ _0452_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8243__B2 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5689__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5057__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7841__I1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5059_ _0391_ _0397_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A4 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8546__A2 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8818_ as2650.r123\[1\]\[7\] _3901_ _3890_ _1852_ _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8749_ _3855_ _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6313__I _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6309__A1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__B2 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5532__A2 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7809__A1 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4768__I _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7144__I _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7285__A2 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8482__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6983__I _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4638__A4 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8234__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__I _4389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7747__C _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6548__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5523__A2 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4678__I _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6100_ _1384_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7276__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8473__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7080_ _2282_ _2283_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8594__B _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _0854_ _1223_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8225__A1 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7982_ _4443_ _2122_ _1455_ _2968_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5302__I _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _1662_ _1674_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8528__A2 _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _2046_ _2068_ _2069_ _2052_ _2067_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5815_ as2650.stack\[0\]\[4\] _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8603_ _1090_ _3682_ _3751_ _3752_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6795_ _1283_ _1911_ _1913_ as2650.r123_2\[2\]\[3\] _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5211__A1 _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6133__I _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8534_ _3639_ _0313_ _3640_ _3686_ _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _1065_ _1035_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8465_ _3619_ _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5677_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7416_ _1189_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4628_ _4208_ _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8396_ _2855_ _3553_ _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7347_ _1288_ _0643_ _2546_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4559_ _4139_ _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7278_ _1066_ _0349_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9017_ _4077_ _4078_ _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6229_ _4201_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8216__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8767__A2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6778__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9170__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5450__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5202__A1 _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5202__B2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6950__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6978__I _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7258__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8455__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8455__B2 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5269__A1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7602__I _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8207__B2 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8861__C _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5441__A1 as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7194__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8930__A2 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5600_ _0930_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6580_ _0650_ _0994_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5531_ _4517_ _0863_ _4286_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5792__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4910__B _4490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8250_ _1097_ _3167_ _3413_ _3254_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7497__A2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ as2650.holding_reg\[6\] _4131_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7201_ _2403_ _2319_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8181_ _3345_ _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5393_ _0722_ _0727_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7132_ _1549_ _2335_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7249__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8446__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8997__A2 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7063_ _1447_ _2218_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6014_ _0762_ _1238_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7965_ _3104_ _2562_ _3118_ _3136_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5432__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4871__I as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6916_ _2121_ _2123_ _1460_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7896_ _1633_ _3044_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _1297_ _2072_ _2073_ as2650.r123_2\[2\]\[4\] _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8921__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6778_ _0545_ _1039_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6932__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5729_ _4503_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8517_ _4269_ _4248_ _4234_ _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8448_ as2650.pc\[13\] _1620_ _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8011__C _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8379_ _2168_ _3537_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5207__I as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6160__A2 _4126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8946__C _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8437__A1 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4781__I _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8912__A2 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6923__A1 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_51_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_51_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5117__I _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6151__A2 _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8428__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7332__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7100__A1 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5662__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7488__B _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7403__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8600__A1 _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__I _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7750_ _4408_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4962_ _0300_ _4327_ _4328_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_75_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6701_ _1930_ _1931_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7681_ _2856_ _2574_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7167__A1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4893_ _4473_ _4474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8903__A2 _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6632_ _1043_ _1871_ _1879_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6914__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ _1771_ _1816_ _1825_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6390__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8302_ _1545_ _2578_ _3384_ _3463_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5514_ _0382_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9282_ _0231_ clknet_leaf_38_wb_clk_i as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6494_ _1748_ _1759_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8233_ _1585_ _3280_ _3396_ _1373_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5445_ _0584_ _0778_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7670__C _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8164_ _3327_ _3329_ _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5376_ _0602_ _0603_ _0711_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7890__A2 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7115_ net54 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4866__I _4446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8095_ _2615_ _3258_ _3261_ _3091_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7046_ _2231_ _2248_ _2250_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5405__A1 _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8997_ _1578_ _1421_ _3022_ _1520_ _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7948_ _3119_ _3120_ _3121_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8006__C _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7879_ _3033_ _1474_ _3050_ _3056_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5708__A2 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6321__I _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8658__A1 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4776__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6196__C _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5644__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6991__I _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7936__A3 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6940__B _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9028__B _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6372__A2 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7327__I _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8649__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8649__B2 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5230_ _4436_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5883__A1 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5161_ _0492_ _0497_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__A2 _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5092_ _4311_ _0309_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8920_ _1632_ _1687_ _3988_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8851_ _2154_ _2923_ _3658_ _3936_ _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7802_ _4451_ _2986_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ _1267_ _1181_ _1284_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5938__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8782_ _4257_ _4464_ _0335_ _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6060__A1 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4945_ _4524_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7733_ _1466_ _4170_ _2923_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8888__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7664_ net39 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4876_ _4454_ _4456_ _4457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_123_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7595_ _0966_ _0832_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7237__I _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6546_ _0544_ _1752_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9334_ _0283_ clknet_leaf_62_wb_clk_i as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7312__A1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6477_ as2650.r123_2\[1\]\[3\] _1726_ _1743_ _1723_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6115__A2 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9265_ _0214_ clknet_leaf_38_wb_clk_i as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8216_ _1091_ _3341_ _3379_ _3380_ _3122_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5428_ _4396_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9196_ _0145_ clknet_leaf_26_wb_clk_i net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4596__I _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4677__A2 as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5874__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8147_ _3266_ _3312_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5359_ _0694_ _4506_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7615__A2 _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8078_ _3245_ as2650.stack\[5\]\[1\] as2650.stack\[4\]\[1\] _0385_ _3246_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8812__A1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7029_ _1206_ _1389_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7379__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7379__B2 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8576__B1 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5220__I _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A1 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8531__I _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8879__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7551__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A1 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7606__A2 as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5617__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9254__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8706__I _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7082__A3 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6226__I _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A1 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4730_ _4310_ _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _4235_ _4241_ _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7542__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6400_ _1675_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7380_ _2512_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4592_ as2650.ins_reg\[0\] _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6896__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6331_ _1353_ _1371_ _1580_ _1592_ _1614_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_127_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8098__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9050_ _4105_ _4106_ _1428_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5305__B1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6262_ _1545_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4659__A2 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5856__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8001_ _2336_ _3169_ _3065_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5213_ _4303_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6193_ _4465_ _0971_ _1154_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_97_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5144_ _0458_ _0460_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5608__A1 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8270__A2 _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ _4274_ _0341_ _0345_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6281__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8903_ as2650.stack\[2\]\[2\] _3976_ _3979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4831__A2 _4409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__I _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8834_ _0583_ _3915_ _3917_ as2650.r123\[2\]\[3\] _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6033__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8765_ _3868_ _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5977_ _0598_ _1224_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7716_ _2765_ _2789_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ _4508_ _4509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8696_ _3827_ _3816_ _3828_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7647_ _1443_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4859_ _4350_ _4419_ _4439_ _4440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7578_ _2750_ _2761_ _2771_ _2773_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9317_ _0266_ clknet_leaf_44_wb_clk_i as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6529_ _1312_ _1697_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9248_ _0197_ clknet_leaf_54_wb_clk_i as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7836__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9277__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9179_ _0128_ clknet_leaf_15_wb_clk_i as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8954__C _4466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__I _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8261__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7430__I _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6272__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7772__A1 _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4586__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__A1 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7827__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7340__I _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4813__A2 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8004__A2 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5900_ _1174_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6880_ _2096_ _2099_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6015__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7212__B1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8555__A3 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ as2650.r123_2\[3\]\[4\] _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7763__A1 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4577__A1 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5762_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8550_ _2648_ _0485_ _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8104__C _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7501_ as2650.pc\[7\] net2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_6_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4713_ _4156_ _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8481_ _2940_ _3634_ _3635_ _3302_ _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5693_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7432_ _2623_ _0642_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _4217_ _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7363_ _2562_ _2351_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4575_ _4155_ _4142_ _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9102_ _0051_ clknet_leaf_10_wb_clk_i as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6314_ _0676_ _0553_ _0664_ _0757_ _0753_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7294_ net53 _2494_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _0822_ _0783_ _0644_ _0519_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_9033_ _1689_ _3058_ _1413_ _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8491__A2 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6176_ _1459_ _1460_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9035__A4 _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__I _4451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5127_ _0456_ _0457_ _0464_ _4385_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8243__A2 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5058_ as2650.stack\[3\]\[9\] _0392_ _0396_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6006__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8817_ _4290_ _0884_ _0915_ _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7754__A1 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8748_ _1898_ _3856_ _3861_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7506__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8679_ as2650.stack\[5\]\[8\] _3816_ _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7809__A2 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8482__A2 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6493__A1 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__A2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4784__I _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8256__I _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8234__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6245__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7745__A1 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8170__A1 as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4959__I _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7335__I _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8473__A2 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8594__C _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6030_ _0823_ _1224_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5287__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8225__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7981_ _3143_ _3032_ _3150_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7984__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6932_ _2141_ _1452_ _2143_ _2144_ _2146_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_70_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6863_ _2081_ _2087_ _2088_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7736__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6539__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8602_ _3551_ _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6414__I _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5814_ _1119_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6794_ _1991_ _2022_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5211__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8533_ _3139_ _0320_ _2439_ _3685_ _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5745_ _1068_ _1059_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8464_ _3618_ _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5676_ _1004_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5474__B _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7415_ _2603_ _2613_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8700__A3 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4869__I _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4627_ _4197_ _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8395_ _0997_ _3508_ _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_102_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6711__A2 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4722__A1 _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7346_ _2544_ _2545_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ as2650.alu_op\[1\] _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7277_ _2467_ _2472_ _2346_ _2478_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9016_ _2993_ _1371_ _2412_ _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6228_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8216__A2 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6159_ _4393_ _1441_ _1442_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9315__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7975__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5450__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7990__A4 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7727__A1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8152__A1 _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput40 net40 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__8455__A2 _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5269__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8207__A2 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7966__A1 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5441__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8391__A1 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7194__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _0862_ _4467_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8143__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4689__I _4117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5461_ _4260_ _0792_ _0794_ _0712_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7200_ net29 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4704__A1 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8180_ _2540_ _3344_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5392_ _0629_ _0618_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7131_ _2334_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8446__A2 _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7062_ _2232_ _2265_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _4445_ _4448_ _1231_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_41_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__I _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7957__A1 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7964_ _3126_ _3129_ _3135_ _3104_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6915_ _2129_ _4195_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7709__A1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7895_ _3064_ _3038_ _3067_ _3070_ _3071_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6846_ _1912_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8382__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8921__A3 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _0443_ _1979_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6932__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8516_ _1511_ _4405_ _4269_ _2279_ _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_5728_ _1052_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4943__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8134__A1 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8134__B2 _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4599__I _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8447_ _2841_ _3601_ _3602_ _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5659_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9107__D _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6696__A1 _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8378_ _2803_ _3496_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7329_ net53 _2526_ _2527_ _1556_ _2529_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8437__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__A1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5120__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6923__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4934__A1 _4169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8428__A2 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6439__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6229__I _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5662__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6611__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _4322_ _4397_ _4129_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _0716_ _1004_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7680_ _2312_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7167__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8364__A1 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4892_ _4472_ _4473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6631_ as2650.stack\[0\]\[14\] _1869_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4925__A1 _4504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6562_ _1796_ _1815_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8116__A1 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6390__A3 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8301_ _2528_ _3462_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5513_ _0384_ as2650.stack\[5\]\[14\] as2650.stack\[4\]\[14\] _0387_ _0847_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9281_ _0230_ clknet_leaf_43_wb_clk_i as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8667__A2 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6493_ _1749_ _1758_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5308__I _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6678__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8232_ _2180_ _0407_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9160__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5444_ as2650.stack\[2\]\[13\] _0588_ _4484_ as2650.stack\[3\]\[13\] _0502_ _0779_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8163_ _0494_ as2650.stack\[1\]\[3\] as2650.stack\[0\]\[3\] _3328_ _3329_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5375_ _0512_ _0690_ _0710_ _0401_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7114_ _2311_ _2316_ _2317_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8094_ _2531_ _3260_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6139__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7045_ net23 _2249_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5043__I _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8996_ _1411_ _1398_ _1524_ _4004_ _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_76_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__A2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7947_ _3119_ _3120_ _2852_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8355__A1 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7878_ _1634_ _1522_ _2260_ _3055_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6829_ _2037_ _2038_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5218__I _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8529__I _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7094__A1 _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6049__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6841__A1 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8346__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7608__I as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9183__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8649__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__I _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5332__A1 _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7343__I _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5160_ as2650.stack\[6\]\[10\] _4476_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5883__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7085__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8282__B1 _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5091_ _4313_ _0428_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8850_ _1512_ _4408_ _1415_ _1436_ _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8585__A1 _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7801_ _2182_ _2309_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5399__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8781_ _4385_ _3881_ _4413_ _3882_ _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5993_ _1185_ _1269_ _1283_ _1218_ _1179_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_52_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6060__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7732_ _4420_ _2922_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4944_ _4319_ _4522_ _4523_ _4524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8337__A1 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4610__A3 _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7663_ _2855_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4875_ _4455_ _4452_ _4456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6899__A1 as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6614_ _1140_ _1117_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7594_ _2788_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7560__A2 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9333_ _0282_ clknet_leaf_63_wb_clk_i as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6545_ as2650.r0\[5\] _0980_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5571__A1 _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9264_ _0213_ clknet_leaf_38_wb_clk_i as2650.stack\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6476_ _1742_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7312__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6115__A3 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8215_ _3078_ _3346_ _3166_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5323__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _0663_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9195_ _0144_ clknet_leaf_27_wb_clk_i net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5874__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8146_ _2492_ _3305_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5358_ _4227_ _4513_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7076__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8077_ _4469_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8812__A2 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5289_ _0621_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7028_ _2232_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9120__D _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7379__A2 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8979_ _0330_ _0971_ _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8328__A1 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7000__A1 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6332__I _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7591__C _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7303__A2 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8500__A1 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4668__A3 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5865__A2 _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7067__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7082__A4 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6042__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9039__B _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4660_ _4237_ _4240_ _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7542__A2 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5553__A1 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ as2650.halted net5 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _1601_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4697__I _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5305__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5305__B2 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6261_ _4392_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8000_ _2161_ _0408_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5212_ as2650.r123\[1\]\[4\] as2650.r123\[0\]\[4\] as2650.r123_2\[1\]\[4\] as2650.r123_2\[0\]\[4\]
+ _4146_ _0339_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5856__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _1475_ _1476_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_124_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9079__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7058__A1 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5143_ _0480_ _0317_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5608__A2 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5074_ _4161_ _0346_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_111_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8902_ _3975_ _1071_ _3978_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6281__A2 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6417__I _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7957__B _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8833_ _3923_ _3924_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7230__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8764_ _3811_ _3870_ _3872_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ as2650.r123_2\[0\]\[3\] _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7715_ _2886_ _2316_ _2906_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4927_ _4507_ _4508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8695_ as2650.stack\[5\]\[13\] _3814_ _3828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7646_ _2677_ _2818_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4858_ _4431_ _4438_ _4439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7692__B _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7577_ _0968_ _2575_ _2772_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4789_ _4360_ _4364_ _4369_ _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_101_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9316_ _0265_ clknet_leaf_47_wb_clk_i as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6528_ as2650.r123_2\[1\]\[5\] _1726_ _1792_ _1723_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9247_ _0196_ clknet_leaf_54_wb_clk_i as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6459_ _1698_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5847__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9178_ _0127_ clknet_leaf_15_wb_clk_i as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7049__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8129_ _3291_ _3295_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7711__I as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8261__A3 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6272__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A3 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7867__B _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7221__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6024__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7772__A2 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__A2 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7158__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6062__I _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__A2 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__A1 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8210__C _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7288__A1 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9221__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5406__I _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7621__I _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8788__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6237__I _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7212__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7212__B2 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ _1135_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8960__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7763__A2 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5761_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4577__A2 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7500_ _2689_ _2316_ _2696_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _4144_ _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8480_ _3212_ _3619_ _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5692_ _1016_ _0987_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8712__A1 _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7431_ _1410_ _2357_ _2627_ _2628_ _2629_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4643_ _4221_ _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7362_ _2366_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_128_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4574_ _4139_ _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9101_ _0050_ clknet_leaf_10_wb_clk_i as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6313_ _1596_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7293_ net30 net29 net54 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9032_ _0793_ _1417_ _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6244_ _0438_ _0330_ _4353_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6175_ _4252_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8779__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _4396_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5057_ _0382_ _0394_ _0395_ _4489_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7203__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6006__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8816_ _3910_ _3911_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8951__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8747_ as2650.stack\[7\]\[3\] _3857_ _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5959_ _0505_ _1223_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8678_ _3814_ _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7629_ _2353_ _2737_ _2739_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5517__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9244__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5517__B2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4740__A2 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7690__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8537__I _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8981__B _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7442__A1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__A2 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7993__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_45_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7745__A2 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8942__A1 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__A1 _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8170__A2 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4731__A2 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7681__A1 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4975__I _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7433__A1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7980_ _0963_ _3148_ _3149_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__9117__CLK clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5444__B1 _4484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7984__A2 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6931_ _0943_ _2145_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8182__I _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _2056_ _2057_ _2081_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_34_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8115__C _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7736__A2 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8933__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8601_ _0742_ _3684_ _3738_ _3750_ _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_34_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5813_ _1119_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6793_ _1915_ _2021_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9267__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8532_ _2983_ _0328_ _3685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5744_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8463_ as2650.pc\[14\] _3617_ _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5675_ _0657_ _0511_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_136_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7414_ _2605_ _2611_ _2612_ _2328_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6172__A1 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4626_ _4178_ _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8394_ _0998_ _3341_ _3550_ _3552_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7345_ _2543_ _1271_ _2443_ _2499_ _2500_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_2_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4557_ _4135_ _4137_ _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7276_ _2167_ _2474_ _2477_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9015_ _1695_ _1522_ _0655_ _2288_ _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4885__I _4465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7672__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6227_ _1511_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6158_ _4124_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5109_ _4361_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6089_ _4221_ _4514_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7975__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4789__A2 _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5986__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6605__I _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8924__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6340__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6163__A1 _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5910__A1 _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput30 net30 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7415__A1 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6218__A2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7966__A2 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5977__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6515__I _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8915__A1 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9047__B _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8143__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6250__I _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5460_ _0793_ _4260_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6154__A1 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7351__B1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4704__A2 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _4334_ _0724_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7130_ _2333_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7654__A1 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6457__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7061_ _4126_ _1379_ _1364_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_115_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6012_ as2650.r123_2\[0\]\[5\] _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
.ends

