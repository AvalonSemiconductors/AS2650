magic
tech gf180mcuD
magscale 1 10
timestamp 1701085154
<< metal1 >>
rect 3602 38558 3614 38610
rect 3666 38607 3678 38610
rect 6738 38607 6750 38610
rect 3666 38561 6750 38607
rect 3666 38558 3678 38561
rect 6738 38558 6750 38561
rect 6802 38558 6814 38610
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 6862 38274 6914 38286
rect 17166 38274 17218 38286
rect 7074 38222 7086 38274
rect 7138 38271 7150 38274
rect 8082 38271 8094 38274
rect 7138 38225 8094 38271
rect 7138 38222 7150 38225
rect 8082 38222 8094 38225
rect 8146 38222 8158 38274
rect 6862 38210 6914 38222
rect 17166 38210 17218 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 30046 38274 30098 38286
rect 30046 38210 30098 38222
rect 33854 38274 33906 38286
rect 33854 38210 33906 38222
rect 37326 38274 37378 38286
rect 37326 38210 37378 38222
rect 7758 38162 7810 38174
rect 7758 38098 7810 38110
rect 8878 38162 8930 38174
rect 11006 38162 11058 38174
rect 9874 38110 9886 38162
rect 9938 38110 9950 38162
rect 11778 38110 11790 38162
rect 11842 38110 11854 38162
rect 8878 38098 8930 38110
rect 11006 38098 11058 38110
rect 4286 38050 4338 38062
rect 7310 38050 7362 38062
rect 1810 37998 1822 38050
rect 1874 37998 1886 38050
rect 3378 37998 3390 38050
rect 3442 37998 3454 38050
rect 5954 37998 5966 38050
rect 6018 37998 6030 38050
rect 4286 37986 4338 37998
rect 7310 37986 7362 37998
rect 9438 38050 9490 38062
rect 14254 38050 14306 38062
rect 12338 37998 12350 38050
rect 12402 37998 12414 38050
rect 13122 37998 13134 38050
rect 13186 37998 13198 38050
rect 9438 37986 9490 37998
rect 14254 37986 14306 37998
rect 15038 38050 15090 38062
rect 19966 38050 20018 38062
rect 19506 37998 19518 38050
rect 19570 37998 19582 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 29026 37998 29038 38050
rect 29090 37998 29102 38050
rect 32834 37998 32846 38050
rect 32898 37998 32910 38050
rect 36418 37998 36430 38050
rect 36482 37998 36494 38050
rect 15038 37986 15090 37998
rect 19966 37986 20018 37998
rect 2382 37938 2434 37950
rect 4958 37938 5010 37950
rect 3602 37886 3614 37938
rect 3666 37886 3678 37938
rect 2382 37874 2434 37886
rect 4958 37874 5010 37886
rect 6526 37938 6578 37950
rect 6526 37874 6578 37886
rect 6750 37938 6802 37950
rect 6750 37874 6802 37886
rect 8206 37938 8258 37950
rect 8206 37874 8258 37886
rect 13358 37938 13410 37950
rect 13358 37874 13410 37886
rect 13470 37938 13522 37950
rect 13470 37874 13522 37886
rect 21310 37938 21362 37950
rect 21310 37874 21362 37886
rect 2046 37826 2098 37838
rect 2046 37762 2098 37774
rect 2718 37826 2770 37838
rect 2718 37762 2770 37774
rect 3950 37826 4002 37838
rect 3950 37762 4002 37774
rect 4622 37826 4674 37838
rect 10446 37826 10498 37838
rect 14590 37826 14642 37838
rect 6178 37774 6190 37826
rect 6242 37774 6254 37826
rect 13906 37774 13918 37826
rect 13970 37774 13982 37826
rect 4622 37762 4674 37774
rect 10446 37762 10498 37774
rect 14590 37762 14642 37774
rect 20974 37826 21026 37838
rect 20974 37762 21026 37774
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 3614 37490 3666 37502
rect 3614 37426 3666 37438
rect 14702 37490 14754 37502
rect 14702 37426 14754 37438
rect 23662 37490 23714 37502
rect 23662 37426 23714 37438
rect 27246 37490 27298 37502
rect 27246 37426 27298 37438
rect 6750 37378 6802 37390
rect 25902 37378 25954 37390
rect 10210 37326 10222 37378
rect 10274 37326 10286 37378
rect 11106 37326 11118 37378
rect 11170 37326 11182 37378
rect 39442 37326 39454 37378
rect 39506 37326 39518 37378
rect 6750 37314 6802 37326
rect 25902 37314 25954 37326
rect 5406 37266 5458 37278
rect 6414 37266 6466 37278
rect 12686 37266 12738 37278
rect 23326 37266 23378 37278
rect 2258 37214 2270 37266
rect 2322 37214 2334 37266
rect 4274 37214 4286 37266
rect 4338 37214 4350 37266
rect 5954 37214 5966 37266
rect 6018 37214 6030 37266
rect 7298 37214 7310 37266
rect 7362 37214 7374 37266
rect 8194 37214 8206 37266
rect 8258 37214 8270 37266
rect 10770 37214 10782 37266
rect 10834 37214 10846 37266
rect 13458 37214 13470 37266
rect 13522 37214 13534 37266
rect 13682 37214 13694 37266
rect 13746 37214 13758 37266
rect 21634 37214 21646 37266
rect 21698 37214 21710 37266
rect 25666 37214 25678 37266
rect 25730 37214 25742 37266
rect 26226 37214 26238 37266
rect 26290 37214 26302 37266
rect 37650 37214 37662 37266
rect 37714 37214 37726 37266
rect 5406 37202 5458 37214
rect 6414 37202 6466 37214
rect 12686 37202 12738 37214
rect 23326 37202 23378 37214
rect 1822 37154 1874 37166
rect 1822 37090 1874 37102
rect 2718 37154 2770 37166
rect 6862 37154 6914 37166
rect 3154 37102 3166 37154
rect 3218 37102 3230 37154
rect 2718 37090 2770 37102
rect 6862 37090 6914 37102
rect 7758 37154 7810 37166
rect 15262 37154 15314 37166
rect 8530 37102 8542 37154
rect 8594 37102 8606 37154
rect 11330 37102 11342 37154
rect 11394 37102 11406 37154
rect 14130 37102 14142 37154
rect 14194 37102 14206 37154
rect 7758 37090 7810 37102
rect 15262 37090 15314 37102
rect 19742 37154 19794 37166
rect 19742 37090 19794 37102
rect 35982 37154 36034 37166
rect 35982 37090 36034 37102
rect 37438 37154 37490 37166
rect 37438 37090 37490 37102
rect 13906 36990 13918 37042
rect 13970 36990 13982 37042
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 3838 36706 3890 36718
rect 3838 36642 3890 36654
rect 2494 36594 2546 36606
rect 2494 36530 2546 36542
rect 3502 36594 3554 36606
rect 4050 36542 4062 36594
rect 4114 36542 4126 36594
rect 11554 36542 11566 36594
rect 11618 36542 11630 36594
rect 14242 36542 14254 36594
rect 14306 36542 14318 36594
rect 15250 36542 15262 36594
rect 15314 36542 15326 36594
rect 16706 36542 16718 36594
rect 16770 36542 16782 36594
rect 3502 36530 3554 36542
rect 2606 36482 2658 36494
rect 2606 36418 2658 36430
rect 2942 36482 2994 36494
rect 5742 36482 5794 36494
rect 4162 36430 4174 36482
rect 4226 36430 4238 36482
rect 4834 36430 4846 36482
rect 4898 36430 4910 36482
rect 2942 36418 2994 36430
rect 5742 36418 5794 36430
rect 5854 36482 5906 36494
rect 5854 36418 5906 36430
rect 5966 36482 6018 36494
rect 12910 36482 12962 36494
rect 6962 36430 6974 36482
rect 7026 36430 7038 36482
rect 9986 36430 9998 36482
rect 10050 36430 10062 36482
rect 12226 36430 12238 36482
rect 12290 36430 12302 36482
rect 12786 36430 12798 36482
rect 12850 36430 12862 36482
rect 13794 36430 13806 36482
rect 13858 36430 13870 36482
rect 14018 36430 14030 36482
rect 14082 36430 14094 36482
rect 15138 36430 15150 36482
rect 15202 36430 15214 36482
rect 16370 36430 16382 36482
rect 16434 36430 16446 36482
rect 17266 36430 17278 36482
rect 17330 36430 17342 36482
rect 5966 36418 6018 36430
rect 12910 36418 12962 36430
rect 11006 36370 11058 36382
rect 5058 36318 5070 36370
rect 5122 36318 5134 36370
rect 8530 36318 8542 36370
rect 8594 36318 8606 36370
rect 15250 36318 15262 36370
rect 15314 36318 15326 36370
rect 11006 36306 11058 36318
rect 1710 36258 1762 36270
rect 7646 36258 7698 36270
rect 2034 36206 2046 36258
rect 2098 36206 2110 36258
rect 6402 36206 6414 36258
rect 6466 36206 6478 36258
rect 1710 36194 1762 36206
rect 7646 36194 7698 36206
rect 8094 36258 8146 36270
rect 14690 36206 14702 36258
rect 14754 36206 14766 36258
rect 17490 36206 17502 36258
rect 17554 36206 17566 36258
rect 8094 36194 8146 36206
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 6862 35922 6914 35934
rect 6862 35858 6914 35870
rect 2046 35810 2098 35822
rect 4398 35810 4450 35822
rect 7310 35810 7362 35822
rect 13694 35810 13746 35822
rect 2370 35758 2382 35810
rect 2434 35758 2446 35810
rect 4834 35758 4846 35810
rect 4898 35758 4910 35810
rect 6290 35758 6302 35810
rect 6354 35758 6366 35810
rect 10098 35758 10110 35810
rect 10162 35758 10174 35810
rect 16146 35758 16158 35810
rect 16210 35758 16222 35810
rect 2046 35746 2098 35758
rect 4398 35746 4450 35758
rect 7310 35746 7362 35758
rect 13694 35746 13746 35758
rect 12574 35698 12626 35710
rect 1810 35646 1822 35698
rect 1874 35646 1886 35698
rect 2594 35646 2606 35698
rect 2658 35646 2670 35698
rect 5282 35646 5294 35698
rect 5346 35646 5358 35698
rect 6402 35646 6414 35698
rect 6466 35646 6478 35698
rect 10994 35646 11006 35698
rect 11058 35646 11070 35698
rect 11218 35646 11230 35698
rect 11282 35646 11294 35698
rect 12574 35634 12626 35646
rect 14590 35698 14642 35710
rect 14590 35634 14642 35646
rect 17390 35698 17442 35710
rect 17390 35634 17442 35646
rect 3166 35586 3218 35598
rect 3166 35522 3218 35534
rect 3614 35586 3666 35598
rect 6066 35534 6078 35586
rect 6130 35534 6142 35586
rect 11666 35534 11678 35586
rect 11730 35534 11742 35586
rect 14018 35534 14030 35586
rect 14082 35534 14094 35586
rect 17826 35534 17838 35586
rect 17890 35534 17902 35586
rect 3614 35522 3666 35534
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 14254 35026 14306 35038
rect 4274 34974 4286 35026
rect 4338 34974 4350 35026
rect 14254 34962 14306 34974
rect 8206 34914 8258 34926
rect 3378 34862 3390 34914
rect 3442 34862 3454 34914
rect 7970 34862 7982 34914
rect 8034 34862 8046 34914
rect 8206 34850 8258 34862
rect 8318 34914 8370 34926
rect 10782 34914 10834 34926
rect 8754 34862 8766 34914
rect 8818 34862 8830 34914
rect 8318 34850 8370 34862
rect 10782 34850 10834 34862
rect 12798 34914 12850 34926
rect 16382 34914 16434 34926
rect 16034 34862 16046 34914
rect 16098 34862 16110 34914
rect 12798 34850 12850 34862
rect 16382 34850 16434 34862
rect 16942 34914 16994 34926
rect 16942 34850 16994 34862
rect 2942 34802 2994 34814
rect 2942 34738 2994 34750
rect 4734 34802 4786 34814
rect 4734 34738 4786 34750
rect 4846 34802 4898 34814
rect 4846 34738 4898 34750
rect 6190 34802 6242 34814
rect 6190 34738 6242 34750
rect 6526 34802 6578 34814
rect 10222 34802 10274 34814
rect 6850 34750 6862 34802
rect 6914 34750 6926 34802
rect 6526 34738 6578 34750
rect 10222 34738 10274 34750
rect 10894 34802 10946 34814
rect 15486 34802 15538 34814
rect 12898 34750 12910 34802
rect 12962 34750 12974 34802
rect 10894 34738 10946 34750
rect 15486 34738 15538 34750
rect 1934 34690 1986 34702
rect 1934 34626 1986 34638
rect 2270 34690 2322 34702
rect 3838 34690 3890 34702
rect 2594 34638 2606 34690
rect 2658 34638 2670 34690
rect 2270 34626 2322 34638
rect 3838 34626 3890 34638
rect 5070 34690 5122 34702
rect 5070 34626 5122 34638
rect 5630 34690 5682 34702
rect 5630 34626 5682 34638
rect 13694 34690 13746 34702
rect 13694 34626 13746 34638
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 7858 34302 7870 34354
rect 7922 34302 7934 34354
rect 6750 34242 6802 34254
rect 11790 34242 11842 34254
rect 2258 34190 2270 34242
rect 2322 34190 2334 34242
rect 4274 34190 4286 34242
rect 4338 34190 4350 34242
rect 8866 34190 8878 34242
rect 8930 34190 8942 34242
rect 6750 34178 6802 34190
rect 11790 34178 11842 34190
rect 11902 34242 11954 34254
rect 11902 34178 11954 34190
rect 12014 34242 12066 34254
rect 18062 34242 18114 34254
rect 16818 34190 16830 34242
rect 16882 34190 16894 34242
rect 12014 34178 12066 34190
rect 18062 34178 18114 34190
rect 19966 34242 20018 34254
rect 19966 34178 20018 34190
rect 5854 34130 5906 34142
rect 9550 34130 9602 34142
rect 2034 34078 2046 34130
rect 2098 34078 2110 34130
rect 2594 34078 2606 34130
rect 2658 34078 2670 34130
rect 6178 34078 6190 34130
rect 6242 34078 6254 34130
rect 8418 34078 8430 34130
rect 8482 34078 8494 34130
rect 5854 34066 5906 34078
rect 9550 34066 9602 34078
rect 9774 34130 9826 34142
rect 9774 34066 9826 34078
rect 13806 34130 13858 34142
rect 13806 34066 13858 34078
rect 14702 34130 14754 34142
rect 16494 34130 16546 34142
rect 16034 34078 16046 34130
rect 16098 34078 16110 34130
rect 14702 34066 14754 34078
rect 16494 34066 16546 34078
rect 17838 34130 17890 34142
rect 17838 34066 17890 34078
rect 18174 34130 18226 34142
rect 18174 34066 18226 34078
rect 13582 34018 13634 34030
rect 3714 33966 3726 34018
rect 3778 33966 3790 34018
rect 8754 33966 8766 34018
rect 8818 33966 8830 34018
rect 12450 33966 12462 34018
rect 12514 33966 12526 34018
rect 13582 33954 13634 33966
rect 15262 34018 15314 34030
rect 18622 34018 18674 34030
rect 15698 33966 15710 34018
rect 15762 33966 15774 34018
rect 15262 33954 15314 33966
rect 18622 33954 18674 33966
rect 14142 33906 14194 33918
rect 10098 33854 10110 33906
rect 10162 33854 10174 33906
rect 14142 33842 14194 33854
rect 19854 33906 19906 33918
rect 19854 33842 19906 33854
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 17614 33570 17666 33582
rect 17614 33506 17666 33518
rect 3490 33406 3502 33458
rect 3554 33406 3566 33458
rect 4834 33406 4846 33458
rect 4898 33406 4910 33458
rect 7074 33406 7086 33458
rect 7138 33406 7150 33458
rect 9202 33406 9214 33458
rect 9266 33406 9278 33458
rect 15586 33406 15598 33458
rect 15650 33406 15662 33458
rect 5630 33346 5682 33358
rect 2258 33294 2270 33346
rect 2322 33294 2334 33346
rect 2818 33294 2830 33346
rect 2882 33294 2894 33346
rect 4386 33294 4398 33346
rect 4450 33294 4462 33346
rect 4722 33294 4734 33346
rect 4786 33294 4798 33346
rect 5630 33282 5682 33294
rect 6862 33346 6914 33358
rect 14030 33346 14082 33358
rect 16270 33346 16322 33358
rect 6962 33294 6974 33346
rect 7026 33294 7038 33346
rect 8642 33294 8654 33346
rect 8706 33294 8718 33346
rect 10210 33294 10222 33346
rect 10274 33294 10286 33346
rect 11778 33294 11790 33346
rect 11842 33294 11854 33346
rect 13570 33294 13582 33346
rect 13634 33294 13646 33346
rect 15026 33294 15038 33346
rect 15090 33294 15102 33346
rect 16034 33294 16046 33346
rect 16098 33294 16110 33346
rect 6862 33282 6914 33294
rect 14030 33282 14082 33294
rect 16270 33282 16322 33294
rect 16494 33346 16546 33358
rect 17054 33346 17106 33358
rect 16706 33294 16718 33346
rect 16770 33294 16782 33346
rect 16494 33282 16546 33294
rect 17054 33282 17106 33294
rect 17726 33346 17778 33358
rect 19854 33346 19906 33358
rect 18050 33294 18062 33346
rect 18114 33294 18126 33346
rect 17726 33282 17778 33294
rect 19854 33282 19906 33294
rect 2494 33234 2546 33246
rect 11454 33234 11506 33246
rect 2930 33182 2942 33234
rect 2994 33182 3006 33234
rect 10322 33182 10334 33234
rect 10386 33182 10398 33234
rect 2494 33170 2546 33182
rect 11454 33170 11506 33182
rect 15262 33234 15314 33246
rect 15262 33170 15314 33182
rect 18286 33234 18338 33246
rect 18286 33170 18338 33182
rect 18398 33234 18450 33246
rect 18398 33170 18450 33182
rect 19182 33234 19234 33246
rect 19182 33170 19234 33182
rect 20078 33234 20130 33246
rect 20078 33170 20130 33182
rect 20302 33234 20354 33246
rect 20302 33170 20354 33182
rect 1822 33122 1874 33134
rect 1822 33058 1874 33070
rect 5182 33122 5234 33134
rect 7758 33122 7810 33134
rect 14702 33122 14754 33134
rect 5954 33070 5966 33122
rect 6018 33070 6030 33122
rect 12002 33070 12014 33122
rect 12066 33070 12078 33122
rect 5182 33058 5234 33070
rect 7758 33058 7810 33070
rect 14702 33058 14754 33070
rect 15486 33122 15538 33134
rect 15486 33058 15538 33070
rect 15598 33122 15650 33134
rect 15598 33058 15650 33070
rect 16382 33122 16434 33134
rect 16382 33058 16434 33070
rect 17278 33122 17330 33134
rect 17278 33058 17330 33070
rect 17502 33122 17554 33134
rect 23438 33122 23490 33134
rect 18834 33070 18846 33122
rect 18898 33070 18910 33122
rect 19506 33070 19518 33122
rect 19570 33070 19582 33122
rect 20626 33070 20638 33122
rect 20690 33070 20702 33122
rect 17502 33058 17554 33070
rect 23438 33058 23490 33070
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 12238 32786 12290 32798
rect 8306 32734 8318 32786
rect 8370 32734 8382 32786
rect 12238 32722 12290 32734
rect 12462 32786 12514 32798
rect 12462 32722 12514 32734
rect 13582 32786 13634 32798
rect 13582 32722 13634 32734
rect 19406 32786 19458 32798
rect 19406 32722 19458 32734
rect 2830 32674 2882 32686
rect 2482 32622 2494 32674
rect 2546 32622 2558 32674
rect 2830 32610 2882 32622
rect 5294 32674 5346 32686
rect 5294 32610 5346 32622
rect 7870 32674 7922 32686
rect 7870 32610 7922 32622
rect 10782 32674 10834 32686
rect 10782 32610 10834 32622
rect 12126 32674 12178 32686
rect 16830 32674 16882 32686
rect 15586 32622 15598 32674
rect 15650 32622 15662 32674
rect 12126 32610 12178 32622
rect 16830 32610 16882 32622
rect 17390 32674 17442 32686
rect 17390 32610 17442 32622
rect 21310 32674 21362 32686
rect 23090 32622 23102 32674
rect 23154 32622 23166 32674
rect 21310 32610 21362 32622
rect 3054 32562 3106 32574
rect 2258 32510 2270 32562
rect 2322 32510 2334 32562
rect 3054 32498 3106 32510
rect 4286 32562 4338 32574
rect 4286 32498 4338 32510
rect 6302 32562 6354 32574
rect 6302 32498 6354 32510
rect 6750 32562 6802 32574
rect 12798 32562 12850 32574
rect 9986 32510 9998 32562
rect 10050 32510 10062 32562
rect 6750 32498 6802 32510
rect 12798 32498 12850 32510
rect 14142 32562 14194 32574
rect 19854 32562 19906 32574
rect 21198 32562 21250 32574
rect 15362 32510 15374 32562
rect 15426 32510 15438 32562
rect 20962 32510 20974 32562
rect 21026 32510 21038 32562
rect 14142 32498 14194 32510
rect 19854 32498 19906 32510
rect 21198 32498 21250 32510
rect 23438 32562 23490 32574
rect 23438 32498 23490 32510
rect 1822 32450 1874 32462
rect 10446 32450 10498 32462
rect 18958 32450 19010 32462
rect 20526 32450 20578 32462
rect 3826 32398 3838 32450
rect 3890 32398 3902 32450
rect 17826 32398 17838 32450
rect 17890 32398 17902 32450
rect 20066 32398 20078 32450
rect 20130 32398 20142 32450
rect 1822 32386 1874 32398
rect 10446 32386 10498 32398
rect 18958 32386 19010 32398
rect 20526 32386 20578 32398
rect 22206 32450 22258 32462
rect 22206 32386 22258 32398
rect 22766 32450 22818 32462
rect 22766 32386 22818 32398
rect 23886 32450 23938 32462
rect 23886 32386 23938 32398
rect 24334 32450 24386 32462
rect 24334 32386 24386 32398
rect 3390 32338 3442 32350
rect 3390 32274 3442 32286
rect 11006 32338 11058 32350
rect 11006 32274 11058 32286
rect 11230 32338 11282 32350
rect 11230 32274 11282 32286
rect 11454 32338 11506 32350
rect 11454 32274 11506 32286
rect 11902 32338 11954 32350
rect 11902 32274 11954 32286
rect 16270 32338 16322 32350
rect 16270 32274 16322 32286
rect 16606 32338 16658 32350
rect 16606 32274 16658 32286
rect 19742 32338 19794 32350
rect 19742 32274 19794 32286
rect 20302 32338 20354 32350
rect 23774 32338 23826 32350
rect 21746 32286 21758 32338
rect 21810 32286 21822 32338
rect 20302 32274 20354 32286
rect 23774 32274 23826 32286
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 2270 32002 2322 32014
rect 2270 31938 2322 31950
rect 10110 32002 10162 32014
rect 10110 31938 10162 31950
rect 2046 31890 2098 31902
rect 2046 31826 2098 31838
rect 3502 31890 3554 31902
rect 10334 31890 10386 31902
rect 16270 31890 16322 31902
rect 4834 31838 4846 31890
rect 4898 31838 4910 31890
rect 6626 31838 6638 31890
rect 6690 31838 6702 31890
rect 11106 31838 11118 31890
rect 11170 31838 11182 31890
rect 3502 31826 3554 31838
rect 10334 31826 10386 31838
rect 16270 31826 16322 31838
rect 21310 31890 21362 31902
rect 21310 31826 21362 31838
rect 22542 31890 22594 31902
rect 22542 31826 22594 31838
rect 24110 31890 24162 31902
rect 24110 31826 24162 31838
rect 4286 31778 4338 31790
rect 5182 31778 5234 31790
rect 4386 31726 4398 31778
rect 4450 31726 4462 31778
rect 4286 31714 4338 31726
rect 5182 31714 5234 31726
rect 6190 31778 6242 31790
rect 7758 31778 7810 31790
rect 8654 31778 8706 31790
rect 6402 31726 6414 31778
rect 6466 31726 6478 31778
rect 7410 31726 7422 31778
rect 7474 31726 7486 31778
rect 7858 31726 7870 31778
rect 7922 31726 7934 31778
rect 6190 31714 6242 31726
rect 7758 31714 7810 31726
rect 8654 31714 8706 31726
rect 8878 31778 8930 31790
rect 8878 31714 8930 31726
rect 13918 31778 13970 31790
rect 15710 31778 15762 31790
rect 15362 31726 15374 31778
rect 15426 31726 15438 31778
rect 13918 31714 13970 31726
rect 15710 31714 15762 31726
rect 16606 31778 16658 31790
rect 16606 31714 16658 31726
rect 16942 31778 16994 31790
rect 16942 31714 16994 31726
rect 17502 31778 17554 31790
rect 17502 31714 17554 31726
rect 21534 31778 21586 31790
rect 21534 31714 21586 31726
rect 22318 31778 22370 31790
rect 22318 31714 22370 31726
rect 23102 31778 23154 31790
rect 23102 31714 23154 31726
rect 23886 31778 23938 31790
rect 23886 31714 23938 31726
rect 7086 31666 7138 31678
rect 7086 31602 7138 31614
rect 9438 31666 9490 31678
rect 9438 31602 9490 31614
rect 15150 31666 15202 31678
rect 15150 31602 15202 31614
rect 15598 31666 15650 31678
rect 15598 31602 15650 31614
rect 16046 31666 16098 31678
rect 16046 31602 16098 31614
rect 2942 31554 2994 31566
rect 10670 31554 10722 31566
rect 2594 31502 2606 31554
rect 2658 31502 2670 31554
rect 9762 31502 9774 31554
rect 9826 31502 9838 31554
rect 2942 31490 2994 31502
rect 10670 31490 10722 31502
rect 11678 31554 11730 31566
rect 11678 31490 11730 31502
rect 12014 31554 12066 31566
rect 17950 31554 18002 31566
rect 22654 31554 22706 31566
rect 12338 31502 12350 31554
rect 12402 31502 12414 31554
rect 14242 31502 14254 31554
rect 14306 31502 14318 31554
rect 16482 31502 16494 31554
rect 16546 31502 16558 31554
rect 21858 31502 21870 31554
rect 21922 31502 21934 31554
rect 12014 31490 12066 31502
rect 17950 31490 18002 31502
rect 22654 31490 22706 31502
rect 22878 31554 22930 31566
rect 22878 31490 22930 31502
rect 23438 31554 23490 31566
rect 23438 31490 23490 31502
rect 23662 31554 23714 31566
rect 23662 31490 23714 31502
rect 23774 31554 23826 31566
rect 23774 31490 23826 31502
rect 24222 31554 24274 31566
rect 24222 31490 24274 31502
rect 24446 31554 24498 31566
rect 24446 31490 24498 31502
rect 24894 31554 24946 31566
rect 24894 31490 24946 31502
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 7870 31218 7922 31230
rect 15598 31218 15650 31230
rect 13010 31166 13022 31218
rect 13074 31166 13086 31218
rect 20974 31218 21026 31230
rect 7870 31154 7922 31166
rect 15598 31154 15650 31166
rect 16494 31162 16546 31174
rect 2718 31106 2770 31118
rect 2034 31054 2046 31106
rect 2098 31054 2110 31106
rect 2718 31042 2770 31054
rect 3166 31106 3218 31118
rect 15150 31106 15202 31118
rect 20974 31154 21026 31166
rect 22542 31218 22594 31230
rect 22542 31154 22594 31166
rect 25454 31218 25506 31230
rect 25454 31154 25506 31166
rect 11330 31054 11342 31106
rect 11394 31054 11406 31106
rect 13234 31054 13246 31106
rect 13298 31054 13310 31106
rect 15922 31054 15934 31106
rect 15986 31054 15998 31106
rect 16494 31098 16546 31110
rect 16606 31106 16658 31118
rect 3166 31042 3218 31054
rect 15150 31042 15202 31054
rect 16606 31042 16658 31054
rect 21310 31106 21362 31118
rect 21310 31042 21362 31054
rect 21422 31106 21474 31118
rect 25230 31106 25282 31118
rect 23426 31054 23438 31106
rect 23490 31054 23502 31106
rect 23986 31054 23998 31106
rect 24050 31054 24062 31106
rect 21422 31042 21474 31054
rect 25230 31042 25282 31054
rect 1710 30994 1762 31006
rect 4286 30994 4338 31006
rect 6526 30994 6578 31006
rect 2482 30942 2494 30994
rect 2546 30942 2558 30994
rect 4722 30942 4734 30994
rect 4786 30942 4798 30994
rect 5618 30942 5630 30994
rect 5682 30942 5694 30994
rect 6066 30942 6078 30994
rect 6130 30942 6142 30994
rect 1710 30930 1762 30942
rect 4286 30930 4338 30942
rect 6526 30930 6578 30942
rect 6862 30994 6914 31006
rect 6862 30930 6914 30942
rect 10222 30994 10274 31006
rect 12910 30994 12962 31006
rect 11666 30942 11678 30994
rect 11730 30942 11742 30994
rect 12114 30942 12126 30994
rect 12178 30942 12190 30994
rect 10222 30930 10274 30942
rect 12910 30930 12962 30942
rect 13694 30994 13746 31006
rect 13694 30930 13746 30942
rect 18622 30994 18674 31006
rect 22206 30994 22258 31006
rect 21970 30942 21982 30994
rect 22034 30942 22046 30994
rect 23090 30942 23102 30994
rect 23154 30942 23166 30994
rect 18622 30930 18674 30942
rect 22206 30930 22258 30942
rect 5182 30882 5234 30894
rect 3826 30830 3838 30882
rect 3890 30830 3902 30882
rect 5182 30818 5234 30830
rect 8430 30882 8482 30894
rect 8430 30818 8482 30830
rect 9998 30882 10050 30894
rect 9998 30818 10050 30830
rect 14366 30882 14418 30894
rect 14366 30818 14418 30830
rect 14702 30882 14754 30894
rect 14702 30818 14754 30830
rect 18398 30882 18450 30894
rect 18398 30818 18450 30830
rect 20526 30882 20578 30894
rect 20526 30818 20578 30830
rect 24334 30882 24386 30894
rect 24334 30818 24386 30830
rect 25342 30882 25394 30894
rect 25342 30818 25394 30830
rect 3054 30770 3106 30782
rect 3054 30706 3106 30718
rect 10446 30770 10498 30782
rect 10446 30706 10498 30718
rect 10782 30770 10834 30782
rect 16606 30770 16658 30782
rect 14130 30718 14142 30770
rect 14194 30767 14206 30770
rect 14354 30767 14366 30770
rect 14194 30721 14366 30767
rect 14194 30718 14206 30721
rect 14354 30718 14366 30721
rect 14418 30718 14430 30770
rect 10782 30706 10834 30718
rect 16606 30706 16658 30718
rect 18958 30770 19010 30782
rect 18958 30706 19010 30718
rect 21422 30770 21474 30782
rect 21422 30706 21474 30718
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 8654 30434 8706 30446
rect 8654 30370 8706 30382
rect 8990 30434 9042 30446
rect 8990 30370 9042 30382
rect 24222 30434 24274 30446
rect 24222 30370 24274 30382
rect 3054 30322 3106 30334
rect 3054 30258 3106 30270
rect 3166 30322 3218 30334
rect 3166 30258 3218 30270
rect 6414 30322 6466 30334
rect 6414 30258 6466 30270
rect 8766 30322 8818 30334
rect 8766 30258 8818 30270
rect 9998 30322 10050 30334
rect 9998 30258 10050 30270
rect 1710 30210 1762 30222
rect 5070 30210 5122 30222
rect 9102 30210 9154 30222
rect 3602 30158 3614 30210
rect 3666 30158 3678 30210
rect 6626 30158 6638 30210
rect 6690 30158 6702 30210
rect 1710 30146 1762 30158
rect 5070 30146 5122 30158
rect 9102 30146 9154 30158
rect 9886 30210 9938 30222
rect 23998 30210 24050 30222
rect 11442 30158 11454 30210
rect 11506 30158 11518 30210
rect 14130 30158 14142 30210
rect 14194 30158 14206 30210
rect 15250 30158 15262 30210
rect 15314 30158 15326 30210
rect 15586 30158 15598 30210
rect 15650 30158 15662 30210
rect 15922 30158 15934 30210
rect 15986 30158 15998 30210
rect 18498 30158 18510 30210
rect 18562 30158 18574 30210
rect 19842 30158 19854 30210
rect 19906 30158 19918 30210
rect 9886 30146 9938 30158
rect 23998 30146 24050 30158
rect 2046 30098 2098 30110
rect 2046 30034 2098 30046
rect 4062 30098 4114 30110
rect 4062 30034 4114 30046
rect 4510 30098 4562 30110
rect 4510 30034 4562 30046
rect 7198 30098 7250 30110
rect 7198 30034 7250 30046
rect 11902 30098 11954 30110
rect 11902 30034 11954 30046
rect 12350 30098 12402 30110
rect 12350 30034 12402 30046
rect 12462 30098 12514 30110
rect 12462 30034 12514 30046
rect 12574 30098 12626 30110
rect 19406 30098 19458 30110
rect 17378 30046 17390 30098
rect 17442 30046 17454 30098
rect 12574 30034 12626 30046
rect 19406 30034 19458 30046
rect 22990 30098 23042 30110
rect 22990 30034 23042 30046
rect 2830 29986 2882 29998
rect 2830 29922 2882 29934
rect 8094 29986 8146 29998
rect 8094 29922 8146 29934
rect 9550 29986 9602 29998
rect 9550 29922 9602 29934
rect 10670 29986 10722 29998
rect 10670 29922 10722 29934
rect 13582 29986 13634 29998
rect 23102 29986 23154 29998
rect 18834 29934 18846 29986
rect 18898 29934 18910 29986
rect 13582 29922 13634 29934
rect 23102 29922 23154 29934
rect 23326 29986 23378 29998
rect 24546 29934 24558 29986
rect 24610 29934 24622 29986
rect 23326 29922 23378 29934
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 2942 29650 2994 29662
rect 2942 29586 2994 29598
rect 8766 29650 8818 29662
rect 8766 29586 8818 29598
rect 14366 29650 14418 29662
rect 14366 29586 14418 29598
rect 15038 29650 15090 29662
rect 15038 29586 15090 29598
rect 15262 29650 15314 29662
rect 15262 29586 15314 29598
rect 16494 29650 16546 29662
rect 16494 29586 16546 29598
rect 18286 29650 18338 29662
rect 18286 29586 18338 29598
rect 18510 29650 18562 29662
rect 18510 29586 18562 29598
rect 18622 29650 18674 29662
rect 18622 29586 18674 29598
rect 2046 29538 2098 29550
rect 2046 29474 2098 29486
rect 4958 29538 5010 29550
rect 4958 29474 5010 29486
rect 6974 29538 7026 29550
rect 6974 29474 7026 29486
rect 8878 29538 8930 29550
rect 23326 29538 23378 29550
rect 19058 29486 19070 29538
rect 19122 29486 19134 29538
rect 21410 29486 21422 29538
rect 21474 29486 21486 29538
rect 21858 29486 21870 29538
rect 21922 29486 21934 29538
rect 8878 29474 8930 29486
rect 23326 29474 23378 29486
rect 23438 29538 23490 29550
rect 23438 29474 23490 29486
rect 2382 29426 2434 29438
rect 8654 29426 8706 29438
rect 1810 29374 1822 29426
rect 1874 29374 1886 29426
rect 3378 29374 3390 29426
rect 3442 29374 3454 29426
rect 4386 29374 4398 29426
rect 4450 29374 4462 29426
rect 6402 29374 6414 29426
rect 6466 29374 6478 29426
rect 2382 29362 2434 29374
rect 8654 29362 8706 29374
rect 9550 29426 9602 29438
rect 9550 29362 9602 29374
rect 9998 29426 10050 29438
rect 9998 29362 10050 29374
rect 11006 29426 11058 29438
rect 11006 29362 11058 29374
rect 11902 29426 11954 29438
rect 11902 29362 11954 29374
rect 12126 29426 12178 29438
rect 12126 29362 12178 29374
rect 12350 29426 12402 29438
rect 14254 29426 14306 29438
rect 13234 29374 13246 29426
rect 13298 29374 13310 29426
rect 14018 29374 14030 29426
rect 14082 29374 14094 29426
rect 12350 29362 12402 29374
rect 14254 29362 14306 29374
rect 14478 29426 14530 29438
rect 14478 29362 14530 29374
rect 14590 29426 14642 29438
rect 14590 29362 14642 29374
rect 15150 29426 15202 29438
rect 19406 29426 19458 29438
rect 15586 29374 15598 29426
rect 15650 29374 15662 29426
rect 18050 29374 18062 29426
rect 18114 29374 18126 29426
rect 15150 29362 15202 29374
rect 19406 29362 19458 29374
rect 21198 29426 21250 29438
rect 21198 29362 21250 29374
rect 23662 29426 23714 29438
rect 23662 29362 23714 29374
rect 3838 29314 3890 29326
rect 10334 29314 10386 29326
rect 7746 29262 7758 29314
rect 7810 29262 7822 29314
rect 3838 29250 3890 29262
rect 10334 29250 10386 29262
rect 10782 29314 10834 29326
rect 10782 29250 10834 29262
rect 11230 29314 11282 29326
rect 11230 29250 11282 29262
rect 11678 29314 11730 29326
rect 11678 29250 11730 29262
rect 12014 29314 12066 29326
rect 16046 29314 16098 29326
rect 20974 29314 21026 29326
rect 13570 29262 13582 29314
rect 13634 29262 13646 29314
rect 15586 29262 15598 29314
rect 15650 29311 15662 29314
rect 15650 29265 15871 29311
rect 15650 29262 15662 29265
rect 12014 29250 12066 29262
rect 15825 29199 15871 29265
rect 16370 29262 16382 29314
rect 16434 29262 16446 29314
rect 18498 29262 18510 29314
rect 18562 29262 18574 29314
rect 16046 29250 16098 29262
rect 16385 29199 16431 29262
rect 20974 29250 21026 29262
rect 15825 29153 16431 29199
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 23214 28866 23266 28878
rect 9874 28814 9886 28866
rect 9938 28814 9950 28866
rect 23214 28802 23266 28814
rect 23662 28866 23714 28878
rect 23662 28802 23714 28814
rect 24782 28866 24834 28878
rect 24782 28802 24834 28814
rect 5070 28754 5122 28766
rect 3602 28702 3614 28754
rect 3666 28702 3678 28754
rect 5070 28690 5122 28702
rect 7646 28754 7698 28766
rect 7646 28690 7698 28702
rect 8094 28754 8146 28766
rect 21310 28754 21362 28766
rect 8978 28702 8990 28754
rect 9042 28702 9054 28754
rect 11890 28702 11902 28754
rect 11954 28702 11966 28754
rect 8094 28690 8146 28702
rect 21310 28690 21362 28702
rect 21758 28754 21810 28766
rect 21758 28690 21810 28702
rect 22990 28754 23042 28766
rect 22990 28690 23042 28702
rect 1710 28642 1762 28654
rect 1710 28578 1762 28590
rect 2830 28642 2882 28654
rect 13694 28642 13746 28654
rect 4162 28590 4174 28642
rect 4226 28590 4238 28642
rect 5618 28590 5630 28642
rect 5682 28590 5694 28642
rect 7186 28590 7198 28642
rect 7250 28590 7262 28642
rect 8866 28590 8878 28642
rect 8930 28590 8942 28642
rect 10434 28590 10446 28642
rect 10498 28590 10510 28642
rect 11442 28590 11454 28642
rect 11506 28590 11518 28642
rect 2830 28578 2882 28590
rect 13694 28578 13746 28590
rect 14590 28642 14642 28654
rect 14590 28578 14642 28590
rect 15262 28642 15314 28654
rect 15262 28578 15314 28590
rect 16606 28642 16658 28654
rect 16606 28578 16658 28590
rect 17502 28642 17554 28654
rect 17502 28578 17554 28590
rect 18622 28642 18674 28654
rect 19406 28642 19458 28654
rect 19058 28590 19070 28642
rect 19122 28590 19134 28642
rect 18622 28578 18674 28590
rect 19406 28578 19458 28590
rect 21534 28642 21586 28654
rect 21534 28578 21586 28590
rect 21982 28642 22034 28654
rect 21982 28578 22034 28590
rect 22430 28642 22482 28654
rect 22430 28578 22482 28590
rect 23886 28642 23938 28654
rect 23886 28578 23938 28590
rect 24110 28642 24162 28654
rect 24110 28578 24162 28590
rect 24894 28642 24946 28654
rect 24894 28578 24946 28590
rect 25342 28642 25394 28654
rect 25342 28578 25394 28590
rect 25678 28642 25730 28654
rect 25678 28578 25730 28590
rect 26238 28642 26290 28654
rect 26238 28578 26290 28590
rect 15710 28530 15762 28542
rect 5730 28478 5742 28530
rect 5794 28478 5806 28530
rect 6178 28478 6190 28530
rect 6242 28478 6254 28530
rect 15710 28466 15762 28478
rect 16046 28530 16098 28542
rect 16046 28466 16098 28478
rect 17166 28530 17218 28542
rect 17166 28466 17218 28478
rect 19294 28530 19346 28542
rect 19294 28466 19346 28478
rect 20190 28530 20242 28542
rect 20190 28466 20242 28478
rect 20302 28530 20354 28542
rect 20302 28466 20354 28478
rect 24334 28530 24386 28542
rect 24334 28466 24386 28478
rect 24670 28530 24722 28542
rect 24670 28466 24722 28478
rect 2046 28418 2098 28430
rect 13358 28418 13410 28430
rect 6626 28366 6638 28418
rect 6690 28366 6702 28418
rect 2046 28354 2098 28366
rect 13358 28354 13410 28366
rect 13582 28418 13634 28430
rect 13582 28354 13634 28366
rect 14030 28418 14082 28430
rect 17278 28418 17330 28430
rect 14914 28366 14926 28418
rect 14978 28366 14990 28418
rect 14030 28354 14082 28366
rect 17278 28354 17330 28366
rect 17838 28418 17890 28430
rect 20526 28418 20578 28430
rect 18274 28366 18286 28418
rect 18338 28366 18350 28418
rect 19842 28366 19854 28418
rect 19906 28366 19918 28418
rect 17838 28354 17890 28366
rect 20526 28354 20578 28366
rect 25118 28418 25170 28430
rect 25118 28354 25170 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 11230 28082 11282 28094
rect 8866 28030 8878 28082
rect 8930 28030 8942 28082
rect 11230 28018 11282 28030
rect 15486 28082 15538 28094
rect 15486 28018 15538 28030
rect 16270 28082 16322 28094
rect 16270 28018 16322 28030
rect 18062 28082 18114 28094
rect 18062 28018 18114 28030
rect 18622 28082 18674 28094
rect 18622 28018 18674 28030
rect 20750 28082 20802 28094
rect 20750 28018 20802 28030
rect 3614 27970 3666 27982
rect 3614 27906 3666 27918
rect 5070 27970 5122 27982
rect 5070 27906 5122 27918
rect 6526 27970 6578 27982
rect 6526 27906 6578 27918
rect 8318 27970 8370 27982
rect 8318 27906 8370 27918
rect 12238 27970 12290 27982
rect 12238 27906 12290 27918
rect 13694 27970 13746 27982
rect 15822 27970 15874 27982
rect 14914 27918 14926 27970
rect 14978 27918 14990 27970
rect 13694 27906 13746 27918
rect 15822 27906 15874 27918
rect 23774 27970 23826 27982
rect 25566 27970 25618 27982
rect 23986 27918 23998 27970
rect 24050 27918 24062 27970
rect 23774 27906 23826 27918
rect 25566 27906 25618 27918
rect 26014 27970 26066 27982
rect 26014 27906 26066 27918
rect 7646 27858 7698 27870
rect 2930 27806 2942 27858
rect 2994 27806 3006 27858
rect 3378 27806 3390 27858
rect 3442 27806 3454 27858
rect 3938 27806 3950 27858
rect 4002 27806 4014 27858
rect 7646 27794 7698 27806
rect 8542 27858 8594 27870
rect 11118 27858 11170 27870
rect 12462 27858 12514 27870
rect 16046 27858 16098 27870
rect 9762 27806 9774 27858
rect 9826 27806 9838 27858
rect 11330 27806 11342 27858
rect 11394 27806 11406 27858
rect 13458 27806 13470 27858
rect 13522 27806 13534 27858
rect 14802 27806 14814 27858
rect 14866 27806 14878 27858
rect 8542 27794 8594 27806
rect 11118 27794 11170 27806
rect 12462 27794 12514 27806
rect 16046 27794 16098 27806
rect 16382 27858 16434 27870
rect 16382 27794 16434 27806
rect 18398 27858 18450 27870
rect 18398 27794 18450 27806
rect 18846 27858 18898 27870
rect 18846 27794 18898 27806
rect 19070 27858 19122 27870
rect 23326 27858 23378 27870
rect 19842 27806 19854 27858
rect 19906 27806 19918 27858
rect 19070 27794 19122 27806
rect 23326 27794 23378 27806
rect 24110 27858 24162 27870
rect 24110 27794 24162 27806
rect 25230 27858 25282 27870
rect 25230 27794 25282 27806
rect 25790 27858 25842 27870
rect 25790 27794 25842 27806
rect 26126 27858 26178 27870
rect 26126 27794 26178 27806
rect 20302 27746 20354 27758
rect 2258 27694 2270 27746
rect 2322 27694 2334 27746
rect 7186 27694 7198 27746
rect 7250 27694 7262 27746
rect 10658 27694 10670 27746
rect 10722 27694 10734 27746
rect 14578 27694 14590 27746
rect 14642 27694 14654 27746
rect 16258 27694 16270 27746
rect 16322 27694 16334 27746
rect 17602 27694 17614 27746
rect 17666 27694 17678 27746
rect 20302 27682 20354 27694
rect 22542 27746 22594 27758
rect 22542 27682 22594 27694
rect 22990 27746 23042 27758
rect 22990 27682 23042 27694
rect 26574 27746 26626 27758
rect 26574 27682 26626 27694
rect 12798 27634 12850 27646
rect 12798 27570 12850 27582
rect 18958 27634 19010 27646
rect 18958 27570 19010 27582
rect 23102 27634 23154 27646
rect 23102 27570 23154 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 19742 27298 19794 27310
rect 11666 27246 11678 27298
rect 11730 27246 11742 27298
rect 19742 27234 19794 27246
rect 21422 27298 21474 27310
rect 21422 27234 21474 27246
rect 22318 27298 22370 27310
rect 26002 27246 26014 27298
rect 26066 27246 26078 27298
rect 22318 27234 22370 27246
rect 20302 27186 20354 27198
rect 4946 27134 4958 27186
rect 5010 27134 5022 27186
rect 9202 27134 9214 27186
rect 9266 27134 9278 27186
rect 12338 27134 12350 27186
rect 12402 27134 12414 27186
rect 13794 27134 13806 27186
rect 13858 27134 13870 27186
rect 20302 27122 20354 27134
rect 23102 27186 23154 27198
rect 23102 27122 23154 27134
rect 7310 27074 7362 27086
rect 3154 27022 3166 27074
rect 3218 27022 3230 27074
rect 5058 27022 5070 27074
rect 5122 27022 5134 27074
rect 6514 27022 6526 27074
rect 6578 27022 6590 27074
rect 7310 27010 7362 27022
rect 7870 27074 7922 27086
rect 14254 27074 14306 27086
rect 9762 27022 9774 27074
rect 9826 27022 9838 27074
rect 10434 27022 10446 27074
rect 10498 27022 10510 27074
rect 11778 27022 11790 27074
rect 11842 27022 11854 27074
rect 7870 27010 7922 27022
rect 14254 27010 14306 27022
rect 14814 27074 14866 27086
rect 22206 27074 22258 27086
rect 15138 27022 15150 27074
rect 15202 27022 15214 27074
rect 16594 27022 16606 27074
rect 16658 27022 16670 27074
rect 17154 27022 17166 27074
rect 17218 27022 17230 27074
rect 18498 27022 18510 27074
rect 18562 27022 18574 27074
rect 23538 27022 23550 27074
rect 23602 27022 23614 27074
rect 24770 27022 24782 27074
rect 24834 27022 24846 27074
rect 26226 27022 26238 27074
rect 26290 27022 26302 27074
rect 14814 27010 14866 27022
rect 22206 27010 22258 27022
rect 5518 26962 5570 26974
rect 2594 26910 2606 26962
rect 2658 26910 2670 26962
rect 3378 26910 3390 26962
rect 3442 26910 3454 26962
rect 5518 26898 5570 26910
rect 7758 26962 7810 26974
rect 7758 26898 7810 26910
rect 19630 26962 19682 26974
rect 19630 26898 19682 26910
rect 22318 26962 22370 26974
rect 26338 26910 26350 26962
rect 26402 26910 26414 26962
rect 22318 26898 22370 26910
rect 7534 26850 7586 26862
rect 19294 26850 19346 26862
rect 16482 26798 16494 26850
rect 16546 26798 16558 26850
rect 18722 26798 18734 26850
rect 18786 26798 18798 26850
rect 7534 26786 7586 26798
rect 19294 26786 19346 26798
rect 19742 26850 19794 26862
rect 19742 26786 19794 26798
rect 21534 26850 21586 26862
rect 21534 26786 21586 26798
rect 21646 26850 21698 26862
rect 21646 26786 21698 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 8430 26514 8482 26526
rect 17390 26514 17442 26526
rect 16706 26462 16718 26514
rect 16770 26462 16782 26514
rect 8430 26450 8482 26462
rect 17390 26450 17442 26462
rect 21646 26514 21698 26526
rect 21646 26450 21698 26462
rect 22318 26514 22370 26526
rect 22318 26450 22370 26462
rect 22878 26514 22930 26526
rect 22878 26450 22930 26462
rect 23774 26514 23826 26526
rect 23774 26450 23826 26462
rect 23998 26514 24050 26526
rect 23998 26450 24050 26462
rect 24334 26514 24386 26526
rect 26674 26462 26686 26514
rect 26738 26462 26750 26514
rect 24334 26450 24386 26462
rect 8766 26402 8818 26414
rect 5282 26350 5294 26402
rect 5346 26350 5358 26402
rect 6514 26350 6526 26402
rect 6578 26350 6590 26402
rect 8766 26338 8818 26350
rect 8878 26402 8930 26414
rect 8878 26338 8930 26350
rect 9998 26402 10050 26414
rect 19294 26402 19346 26414
rect 15362 26350 15374 26402
rect 15426 26350 15438 26402
rect 9998 26338 10050 26350
rect 19294 26338 19346 26350
rect 21422 26402 21474 26414
rect 21422 26338 21474 26350
rect 22654 26402 22706 26414
rect 28478 26402 28530 26414
rect 24658 26350 24670 26402
rect 24722 26350 24734 26402
rect 25218 26350 25230 26402
rect 25282 26350 25294 26402
rect 26786 26350 26798 26402
rect 26850 26350 26862 26402
rect 27570 26350 27582 26402
rect 27634 26350 27646 26402
rect 28130 26350 28142 26402
rect 28194 26350 28206 26402
rect 22654 26338 22706 26350
rect 28478 26338 28530 26350
rect 2606 26290 2658 26302
rect 7870 26290 7922 26302
rect 3154 26238 3166 26290
rect 3218 26238 3230 26290
rect 5954 26238 5966 26290
rect 6018 26238 6030 26290
rect 2606 26226 2658 26238
rect 7870 26226 7922 26238
rect 9102 26290 9154 26302
rect 19182 26290 19234 26302
rect 11554 26238 11566 26290
rect 11618 26238 11630 26290
rect 13010 26238 13022 26290
rect 13074 26238 13086 26290
rect 13234 26238 13246 26290
rect 13298 26238 13310 26290
rect 13570 26238 13582 26290
rect 13634 26238 13646 26290
rect 14242 26238 14254 26290
rect 14306 26238 14318 26290
rect 16482 26238 16494 26290
rect 16546 26238 16558 26290
rect 18386 26238 18398 26290
rect 18450 26238 18462 26290
rect 9102 26226 9154 26238
rect 19182 26226 19234 26238
rect 19518 26290 19570 26302
rect 19518 26226 19570 26238
rect 20638 26290 20690 26302
rect 20638 26226 20690 26238
rect 21086 26290 21138 26302
rect 21086 26226 21138 26238
rect 21310 26290 21362 26302
rect 21310 26226 21362 26238
rect 23214 26290 23266 26302
rect 23214 26226 23266 26238
rect 23326 26290 23378 26302
rect 25778 26238 25790 26290
rect 25842 26238 25854 26290
rect 26226 26238 26238 26290
rect 26290 26238 26302 26290
rect 27234 26238 27246 26290
rect 27298 26238 27310 26290
rect 23326 26226 23378 26238
rect 17950 26178 18002 26190
rect 19966 26178 20018 26190
rect 2146 26126 2158 26178
rect 2210 26126 2222 26178
rect 4050 26126 4062 26178
rect 4114 26126 4126 26178
rect 8082 26126 8094 26178
rect 8146 26126 8158 26178
rect 10882 26126 10894 26178
rect 10946 26126 10958 26178
rect 18722 26126 18734 26178
rect 18786 26126 18798 26178
rect 17950 26114 18002 26126
rect 19966 26114 20018 26126
rect 20190 26178 20242 26190
rect 20190 26114 20242 26126
rect 23886 26178 23938 26190
rect 23886 26114 23938 26126
rect 20414 26066 20466 26078
rect 20414 26002 20466 26014
rect 22542 26066 22594 26078
rect 22542 26002 22594 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 17378 25678 17390 25730
rect 17442 25678 17454 25730
rect 14478 25618 14530 25630
rect 4946 25566 4958 25618
rect 5010 25566 5022 25618
rect 5842 25566 5854 25618
rect 5906 25566 5918 25618
rect 9202 25566 9214 25618
rect 9266 25566 9278 25618
rect 12898 25566 12910 25618
rect 12962 25566 12974 25618
rect 13906 25566 13918 25618
rect 13970 25566 13982 25618
rect 14478 25554 14530 25566
rect 19630 25618 19682 25630
rect 19630 25554 19682 25566
rect 7646 25506 7698 25518
rect 17838 25506 17890 25518
rect 1810 25454 1822 25506
rect 1874 25454 1886 25506
rect 3378 25454 3390 25506
rect 3442 25454 3454 25506
rect 5058 25454 5070 25506
rect 5122 25454 5134 25506
rect 5954 25454 5966 25506
rect 6018 25454 6030 25506
rect 6178 25454 6190 25506
rect 6242 25454 6254 25506
rect 9538 25454 9550 25506
rect 9602 25454 9614 25506
rect 10994 25454 11006 25506
rect 11058 25454 11070 25506
rect 11778 25454 11790 25506
rect 11842 25454 11854 25506
rect 12786 25454 12798 25506
rect 12850 25454 12862 25506
rect 14802 25454 14814 25506
rect 14866 25454 14878 25506
rect 15922 25454 15934 25506
rect 15986 25454 15998 25506
rect 17266 25454 17278 25506
rect 17330 25454 17342 25506
rect 7646 25442 7698 25454
rect 17838 25442 17890 25454
rect 19406 25506 19458 25518
rect 20514 25454 20526 25506
rect 20578 25454 20590 25506
rect 24882 25454 24894 25506
rect 24946 25454 24958 25506
rect 25330 25454 25342 25506
rect 25394 25454 25406 25506
rect 19406 25442 19458 25454
rect 7310 25394 7362 25406
rect 4498 25342 4510 25394
rect 4562 25342 4574 25394
rect 7310 25330 7362 25342
rect 17726 25394 17778 25406
rect 19518 25394 19570 25406
rect 18050 25342 18062 25394
rect 18114 25342 18126 25394
rect 18610 25342 18622 25394
rect 18674 25342 18686 25394
rect 17726 25330 17778 25342
rect 19518 25330 19570 25342
rect 19742 25394 19794 25406
rect 19742 25330 19794 25342
rect 19966 25394 20018 25406
rect 19966 25330 20018 25342
rect 23774 25394 23826 25406
rect 23774 25330 23826 25342
rect 25790 25394 25842 25406
rect 25790 25330 25842 25342
rect 27246 25394 27298 25406
rect 27246 25330 27298 25342
rect 2046 25282 2098 25294
rect 7534 25282 7586 25294
rect 6514 25230 6526 25282
rect 6578 25230 6590 25282
rect 2046 25218 2098 25230
rect 7534 25218 7586 25230
rect 7758 25282 7810 25294
rect 7758 25218 7810 25230
rect 13470 25282 13522 25294
rect 27358 25282 27410 25294
rect 20738 25230 20750 25282
rect 20802 25230 20814 25282
rect 26786 25230 26798 25282
rect 26850 25230 26862 25282
rect 13470 25218 13522 25230
rect 27358 25218 27410 25230
rect 27582 25282 27634 25294
rect 27582 25218 27634 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 4062 24946 4114 24958
rect 4062 24882 4114 24894
rect 8878 24946 8930 24958
rect 8878 24882 8930 24894
rect 15262 24946 15314 24958
rect 17502 24946 17554 24958
rect 15362 24894 15374 24946
rect 15426 24894 15438 24946
rect 15262 24882 15314 24894
rect 17502 24882 17554 24894
rect 20078 24946 20130 24958
rect 20078 24882 20130 24894
rect 21646 24946 21698 24958
rect 21646 24882 21698 24894
rect 22094 24946 22146 24958
rect 22094 24882 22146 24894
rect 22766 24946 22818 24958
rect 22766 24882 22818 24894
rect 2046 24834 2098 24846
rect 2046 24770 2098 24782
rect 2382 24834 2434 24846
rect 2382 24770 2434 24782
rect 2718 24834 2770 24846
rect 11790 24834 11842 24846
rect 18958 24834 19010 24846
rect 3602 24782 3614 24834
rect 3666 24782 3678 24834
rect 5730 24782 5742 24834
rect 5794 24782 5806 24834
rect 6402 24782 6414 24834
rect 6466 24782 6478 24834
rect 9874 24782 9886 24834
rect 9938 24782 9950 24834
rect 14354 24782 14366 24834
rect 14418 24782 14430 24834
rect 16034 24782 16046 24834
rect 16098 24782 16110 24834
rect 18610 24782 18622 24834
rect 18674 24782 18686 24834
rect 2718 24770 2770 24782
rect 11790 24770 11842 24782
rect 18958 24770 19010 24782
rect 19182 24834 19234 24846
rect 23998 24834 24050 24846
rect 20850 24782 20862 24834
rect 20914 24782 20926 24834
rect 26114 24782 26126 24834
rect 26178 24782 26190 24834
rect 27010 24782 27022 24834
rect 27074 24782 27086 24834
rect 19182 24770 19234 24782
rect 23998 24770 24050 24782
rect 1710 24722 1762 24734
rect 4174 24722 4226 24734
rect 3378 24670 3390 24722
rect 3442 24670 3454 24722
rect 1710 24658 1762 24670
rect 4174 24658 4226 24670
rect 4398 24722 4450 24734
rect 17390 24722 17442 24734
rect 5954 24670 5966 24722
rect 6018 24670 6030 24722
rect 6514 24670 6526 24722
rect 6578 24670 6590 24722
rect 9538 24670 9550 24722
rect 9602 24670 9614 24722
rect 10658 24670 10670 24722
rect 10722 24670 10734 24722
rect 12674 24670 12686 24722
rect 12738 24670 12750 24722
rect 15586 24670 15598 24722
rect 15650 24670 15662 24722
rect 15922 24670 15934 24722
rect 15986 24670 15998 24722
rect 4398 24658 4450 24670
rect 17390 24658 17442 24670
rect 17614 24722 17666 24734
rect 17614 24658 17666 24670
rect 18062 24722 18114 24734
rect 18062 24658 18114 24670
rect 18286 24722 18338 24734
rect 18286 24658 18338 24670
rect 19406 24722 19458 24734
rect 19966 24722 20018 24734
rect 19618 24670 19630 24722
rect 19682 24670 19694 24722
rect 19406 24658 19458 24670
rect 19966 24658 20018 24670
rect 20190 24722 20242 24734
rect 23774 24722 23826 24734
rect 20514 24670 20526 24722
rect 20578 24670 20590 24722
rect 21074 24670 21086 24722
rect 21138 24670 21150 24722
rect 20190 24658 20242 24670
rect 23774 24658 23826 24670
rect 24110 24722 24162 24734
rect 28366 24722 28418 24734
rect 24322 24670 24334 24722
rect 24386 24670 24398 24722
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 24110 24658 24162 24670
rect 28366 24658 28418 24670
rect 8766 24610 8818 24622
rect 23326 24610 23378 24622
rect 8082 24558 8094 24610
rect 8146 24558 8158 24610
rect 10210 24558 10222 24610
rect 10274 24558 10286 24610
rect 14018 24558 14030 24610
rect 14082 24558 14094 24610
rect 19506 24558 19518 24610
rect 19570 24558 19582 24610
rect 25330 24558 25342 24610
rect 25394 24558 25406 24610
rect 8766 24546 8818 24558
rect 23326 24546 23378 24558
rect 4062 24498 4114 24510
rect 4062 24434 4114 24446
rect 8654 24498 8706 24510
rect 8654 24434 8706 24446
rect 24782 24498 24834 24510
rect 24782 24434 24834 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 21422 24162 21474 24174
rect 11778 24110 11790 24162
rect 11842 24110 11854 24162
rect 19394 24110 19406 24162
rect 19458 24159 19470 24162
rect 19458 24113 19903 24159
rect 19458 24110 19470 24113
rect 2494 24050 2546 24062
rect 2494 23986 2546 23998
rect 2942 24050 2994 24062
rect 2942 23986 2994 23998
rect 4734 24050 4786 24062
rect 4734 23986 4786 23998
rect 10782 24050 10834 24062
rect 19857 24050 19903 24113
rect 21422 24098 21474 24110
rect 28142 24050 28194 24062
rect 19842 23998 19854 24050
rect 19906 23998 19918 24050
rect 10782 23986 10834 23998
rect 28142 23986 28194 23998
rect 3950 23938 4002 23950
rect 1922 23886 1934 23938
rect 1986 23886 1998 23938
rect 3950 23874 4002 23886
rect 4286 23938 4338 23950
rect 7646 23938 7698 23950
rect 14142 23938 14194 23950
rect 5618 23886 5630 23938
rect 5682 23886 5694 23938
rect 6626 23886 6638 23938
rect 6690 23886 6702 23938
rect 8418 23886 8430 23938
rect 8482 23886 8494 23938
rect 10098 23886 10110 23938
rect 10162 23886 10174 23938
rect 11666 23886 11678 23938
rect 11730 23886 11742 23938
rect 12114 23886 12126 23938
rect 12178 23886 12190 23938
rect 12786 23886 12798 23938
rect 12850 23886 12862 23938
rect 4286 23874 4338 23886
rect 7646 23874 7698 23886
rect 14142 23874 14194 23886
rect 14702 23938 14754 23950
rect 17726 23938 17778 23950
rect 19742 23938 19794 23950
rect 15362 23886 15374 23938
rect 15426 23886 15438 23938
rect 17266 23886 17278 23938
rect 17330 23886 17342 23938
rect 18946 23886 18958 23938
rect 19010 23886 19022 23938
rect 14702 23874 14754 23886
rect 17726 23874 17778 23886
rect 19742 23874 19794 23886
rect 19854 23938 19906 23950
rect 19854 23874 19906 23886
rect 20302 23938 20354 23950
rect 20302 23874 20354 23886
rect 20526 23938 20578 23950
rect 20526 23874 20578 23886
rect 21310 23938 21362 23950
rect 23998 23938 24050 23950
rect 23650 23886 23662 23938
rect 23714 23886 23726 23938
rect 26898 23886 26910 23938
rect 26962 23886 26974 23938
rect 21310 23874 21362 23886
rect 23998 23874 24050 23886
rect 4174 23826 4226 23838
rect 4174 23762 4226 23774
rect 4622 23826 4674 23838
rect 4622 23762 4674 23774
rect 5070 23826 5122 23838
rect 7310 23826 7362 23838
rect 5842 23774 5854 23826
rect 5906 23774 5918 23826
rect 5070 23762 5122 23774
rect 7310 23762 7362 23774
rect 7422 23826 7474 23838
rect 24558 23826 24610 23838
rect 8194 23774 8206 23826
rect 8258 23774 8270 23826
rect 10322 23774 10334 23826
rect 10386 23774 10398 23826
rect 12898 23774 12910 23826
rect 12962 23774 12974 23826
rect 15810 23774 15822 23826
rect 15874 23774 15886 23826
rect 21858 23774 21870 23826
rect 21922 23774 21934 23826
rect 27234 23774 27246 23826
rect 27298 23774 27310 23826
rect 27794 23774 27806 23826
rect 27858 23774 27870 23826
rect 7422 23762 7474 23774
rect 24558 23762 24610 23774
rect 1710 23714 1762 23726
rect 1710 23650 1762 23662
rect 4846 23714 4898 23726
rect 14926 23714 14978 23726
rect 6626 23662 6638 23714
rect 6690 23662 6702 23714
rect 4846 23650 4898 23662
rect 14926 23650 14978 23662
rect 20414 23714 20466 23726
rect 20414 23650 20466 23662
rect 21422 23714 21474 23726
rect 21422 23650 21474 23662
rect 22654 23714 22706 23726
rect 22654 23650 22706 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 2270 23378 2322 23390
rect 2270 23314 2322 23326
rect 6862 23378 6914 23390
rect 25566 23378 25618 23390
rect 16706 23326 16718 23378
rect 16770 23326 16782 23378
rect 23650 23326 23662 23378
rect 23714 23326 23726 23378
rect 6862 23314 6914 23326
rect 25566 23314 25618 23326
rect 17390 23266 17442 23278
rect 5506 23214 5518 23266
rect 5570 23214 5582 23266
rect 8306 23214 8318 23266
rect 8370 23214 8382 23266
rect 15026 23214 15038 23266
rect 15090 23214 15102 23266
rect 16146 23214 16158 23266
rect 16210 23214 16222 23266
rect 17390 23202 17442 23214
rect 18622 23266 18674 23278
rect 18622 23202 18674 23214
rect 18734 23266 18786 23278
rect 26910 23266 26962 23278
rect 22418 23214 22430 23266
rect 22482 23214 22494 23266
rect 23762 23214 23774 23266
rect 23826 23214 23838 23266
rect 24322 23214 24334 23266
rect 24386 23214 24398 23266
rect 18734 23202 18786 23214
rect 26910 23202 26962 23214
rect 1934 23154 1986 23166
rect 1934 23090 1986 23102
rect 3838 23154 3890 23166
rect 17614 23154 17666 23166
rect 5282 23102 5294 23154
rect 5346 23102 5358 23154
rect 7746 23102 7758 23154
rect 7810 23102 7822 23154
rect 8082 23102 8094 23154
rect 8146 23102 8158 23154
rect 9090 23102 9102 23154
rect 9154 23102 9166 23154
rect 10210 23102 10222 23154
rect 10274 23102 10286 23154
rect 11330 23102 11342 23154
rect 11394 23102 11406 23154
rect 12450 23102 12462 23154
rect 12514 23102 12526 23154
rect 13234 23102 13246 23154
rect 13298 23102 13310 23154
rect 13906 23102 13918 23154
rect 13970 23102 13982 23154
rect 16482 23102 16494 23154
rect 16546 23102 16558 23154
rect 3838 23090 3890 23102
rect 17614 23090 17666 23102
rect 17838 23154 17890 23166
rect 18958 23154 19010 23166
rect 26462 23154 26514 23166
rect 18050 23102 18062 23154
rect 18114 23102 18126 23154
rect 19506 23102 19518 23154
rect 19570 23102 19582 23154
rect 20962 23102 20974 23154
rect 21026 23102 21038 23154
rect 22306 23102 22318 23154
rect 22370 23102 22382 23154
rect 24546 23102 24558 23154
rect 24610 23102 24622 23154
rect 17838 23090 17890 23102
rect 18958 23090 19010 23102
rect 26462 23090 26514 23102
rect 27358 23154 27410 23166
rect 27358 23090 27410 23102
rect 27582 23154 27634 23166
rect 27582 23090 27634 23102
rect 27806 23154 27858 23166
rect 28366 23154 28418 23166
rect 28130 23102 28142 23154
rect 28194 23102 28206 23154
rect 27806 23090 27858 23102
rect 28366 23090 28418 23102
rect 28478 23154 28530 23166
rect 28478 23090 28530 23102
rect 2718 23042 2770 23054
rect 2718 22978 2770 22990
rect 7422 23042 7474 23054
rect 7422 22978 7474 22990
rect 10110 23042 10162 23054
rect 17726 23042 17778 23054
rect 26686 23042 26738 23054
rect 11106 22990 11118 23042
rect 11170 22990 11182 23042
rect 22754 22990 22766 23042
rect 22818 22990 22830 23042
rect 10110 22978 10162 22990
rect 17726 22978 17778 22990
rect 26686 22978 26738 22990
rect 6078 22930 6130 22942
rect 1810 22878 1822 22930
rect 1874 22927 1886 22930
rect 2706 22927 2718 22930
rect 1874 22881 2718 22927
rect 1874 22878 1886 22881
rect 2706 22878 2718 22881
rect 2770 22878 2782 22930
rect 6078 22866 6130 22878
rect 26014 22930 26066 22942
rect 26014 22866 26066 22878
rect 26238 22930 26290 22942
rect 28914 22878 28926 22930
rect 28978 22878 28990 22930
rect 26238 22866 26290 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 5070 22594 5122 22606
rect 5070 22530 5122 22542
rect 5966 22594 6018 22606
rect 5966 22530 6018 22542
rect 6638 22594 6690 22606
rect 8754 22542 8766 22594
rect 8818 22542 8830 22594
rect 24546 22542 24558 22594
rect 24610 22591 24622 22594
rect 25106 22591 25118 22594
rect 24610 22545 25118 22591
rect 24610 22542 24622 22545
rect 25106 22542 25118 22545
rect 25170 22542 25182 22594
rect 6638 22530 6690 22542
rect 7982 22482 8034 22494
rect 18510 22482 18562 22494
rect 4162 22430 4174 22482
rect 4226 22430 4238 22482
rect 10434 22430 10446 22482
rect 10498 22430 10510 22482
rect 13570 22430 13582 22482
rect 13634 22430 13646 22482
rect 7982 22418 8034 22430
rect 18510 22418 18562 22430
rect 18734 22482 18786 22494
rect 18734 22418 18786 22430
rect 20638 22482 20690 22494
rect 20638 22418 20690 22430
rect 24222 22482 24274 22494
rect 24222 22418 24274 22430
rect 2942 22370 2994 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 2706 22318 2718 22370
rect 2770 22318 2782 22370
rect 2942 22306 2994 22318
rect 3166 22370 3218 22382
rect 4286 22370 4338 22382
rect 9774 22370 9826 22382
rect 12238 22370 12290 22382
rect 3378 22318 3390 22370
rect 3442 22318 3454 22370
rect 8530 22318 8542 22370
rect 8594 22318 8606 22370
rect 10210 22318 10222 22370
rect 10274 22318 10286 22370
rect 3166 22306 3218 22318
rect 4286 22306 4338 22318
rect 9774 22306 9826 22318
rect 12238 22306 12290 22318
rect 12574 22370 12626 22382
rect 18846 22370 18898 22382
rect 13794 22318 13806 22370
rect 13858 22318 13870 22370
rect 14914 22318 14926 22370
rect 14978 22318 14990 22370
rect 16146 22318 16158 22370
rect 16210 22318 16222 22370
rect 16930 22318 16942 22370
rect 16994 22318 17006 22370
rect 17154 22318 17166 22370
rect 17218 22318 17230 22370
rect 17490 22318 17502 22370
rect 17554 22318 17566 22370
rect 12574 22306 12626 22318
rect 18846 22306 18898 22318
rect 19182 22370 19234 22382
rect 19182 22306 19234 22318
rect 19294 22370 19346 22382
rect 19294 22306 19346 22318
rect 19630 22370 19682 22382
rect 23550 22370 23602 22382
rect 25342 22370 25394 22382
rect 27694 22370 27746 22382
rect 19842 22318 19854 22370
rect 19906 22318 19918 22370
rect 22642 22318 22654 22370
rect 22706 22318 22718 22370
rect 23874 22318 23886 22370
rect 23938 22318 23950 22370
rect 25890 22318 25902 22370
rect 25954 22318 25966 22370
rect 19630 22306 19682 22318
rect 23550 22306 23602 22318
rect 25342 22306 25394 22318
rect 27694 22306 27746 22318
rect 3726 22258 3778 22270
rect 3726 22194 3778 22206
rect 5742 22258 5794 22270
rect 5742 22194 5794 22206
rect 6414 22258 6466 22270
rect 6414 22194 6466 22206
rect 12462 22258 12514 22270
rect 13570 22206 13582 22258
rect 13634 22206 13646 22258
rect 15810 22218 15822 22270
rect 15874 22218 15886 22270
rect 20750 22258 20802 22270
rect 26462 22258 26514 22270
rect 17714 22206 17726 22258
rect 17778 22206 17790 22258
rect 21858 22206 21870 22258
rect 21922 22206 21934 22258
rect 22418 22206 22430 22258
rect 22482 22206 22494 22258
rect 12462 22194 12514 22206
rect 20750 22194 20802 22206
rect 26462 22194 26514 22206
rect 2046 22146 2098 22158
rect 2046 22082 2098 22094
rect 3054 22146 3106 22158
rect 3054 22082 3106 22094
rect 3950 22146 4002 22158
rect 3950 22082 4002 22094
rect 4174 22146 4226 22158
rect 4174 22082 4226 22094
rect 4846 22146 4898 22158
rect 4846 22082 4898 22094
rect 4958 22146 5010 22158
rect 4958 22082 5010 22094
rect 5854 22146 5906 22158
rect 5854 22082 5906 22094
rect 6526 22146 6578 22158
rect 6526 22082 6578 22094
rect 7422 22146 7474 22158
rect 18174 22146 18226 22158
rect 14802 22094 14814 22146
rect 14866 22094 14878 22146
rect 7422 22082 7474 22094
rect 18174 22082 18226 22094
rect 20302 22146 20354 22158
rect 20302 22082 20354 22094
rect 20526 22146 20578 22158
rect 24110 22146 24162 22158
rect 22194 22094 22206 22146
rect 22258 22094 22270 22146
rect 20526 22082 20578 22094
rect 24110 22082 24162 22094
rect 24558 22146 24610 22158
rect 24558 22082 24610 22094
rect 25006 22146 25058 22158
rect 25006 22082 25058 22094
rect 25454 22146 25506 22158
rect 25454 22082 25506 22094
rect 25678 22146 25730 22158
rect 25678 22082 25730 22094
rect 28254 22146 28306 22158
rect 28254 22082 28306 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 2942 21810 2994 21822
rect 2370 21758 2382 21810
rect 2434 21758 2446 21810
rect 2942 21746 2994 21758
rect 3166 21810 3218 21822
rect 9998 21810 10050 21822
rect 3826 21758 3838 21810
rect 3890 21758 3902 21810
rect 3166 21746 3218 21758
rect 9998 21746 10050 21758
rect 10110 21810 10162 21822
rect 10110 21746 10162 21758
rect 11678 21810 11730 21822
rect 11678 21746 11730 21758
rect 12686 21810 12738 21822
rect 21758 21810 21810 21822
rect 21298 21758 21310 21810
rect 21362 21758 21374 21810
rect 12686 21746 12738 21758
rect 21758 21746 21810 21758
rect 26686 21810 26738 21822
rect 26686 21746 26738 21758
rect 2046 21698 2098 21710
rect 9662 21698 9714 21710
rect 4386 21646 4398 21698
rect 4450 21646 4462 21698
rect 5506 21646 5518 21698
rect 5570 21646 5582 21698
rect 2046 21634 2098 21646
rect 9662 21634 9714 21646
rect 11566 21698 11618 21710
rect 11566 21634 11618 21646
rect 14030 21698 14082 21710
rect 22878 21698 22930 21710
rect 25566 21698 25618 21710
rect 17490 21646 17502 21698
rect 17554 21646 17566 21698
rect 21410 21646 21422 21698
rect 21474 21646 21486 21698
rect 24210 21646 24222 21698
rect 24274 21646 24286 21698
rect 27458 21646 27470 21698
rect 27522 21646 27534 21698
rect 28690 21646 28702 21698
rect 28754 21646 28766 21698
rect 14030 21634 14082 21646
rect 22878 21634 22930 21646
rect 25566 21634 25618 21646
rect 9886 21586 9938 21598
rect 2706 21534 2718 21586
rect 2770 21534 2782 21586
rect 3378 21534 3390 21586
rect 3442 21534 3454 21586
rect 3714 21534 3726 21586
rect 3778 21534 3790 21586
rect 6290 21534 6302 21586
rect 6354 21534 6366 21586
rect 7298 21534 7310 21586
rect 7362 21534 7374 21586
rect 8642 21534 8654 21586
rect 8706 21534 8718 21586
rect 9886 21522 9938 21534
rect 10446 21586 10498 21598
rect 10446 21522 10498 21534
rect 11006 21586 11058 21598
rect 11006 21522 11058 21534
rect 13022 21586 13074 21598
rect 13022 21522 13074 21534
rect 13246 21586 13298 21598
rect 22430 21586 22482 21598
rect 15698 21534 15710 21586
rect 15762 21534 15774 21586
rect 17378 21534 17390 21586
rect 17442 21534 17454 21586
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 20850 21534 20862 21586
rect 20914 21534 20926 21586
rect 13246 21522 13298 21534
rect 22430 21522 22482 21534
rect 22654 21586 22706 21598
rect 22654 21522 22706 21534
rect 23998 21586 24050 21598
rect 26238 21586 26290 21598
rect 24322 21534 24334 21586
rect 24386 21534 24398 21586
rect 28130 21534 28142 21586
rect 28194 21534 28206 21586
rect 28578 21534 28590 21586
rect 28642 21534 28654 21586
rect 23998 21522 24050 21534
rect 26238 21522 26290 21534
rect 12126 21474 12178 21486
rect 16830 21474 16882 21486
rect 3266 21422 3278 21474
rect 3330 21422 3342 21474
rect 15362 21422 15374 21474
rect 15426 21422 15438 21474
rect 12126 21410 12178 21422
rect 16830 21410 16882 21422
rect 23774 21474 23826 21486
rect 28802 21422 28814 21474
rect 28866 21422 28878 21474
rect 23774 21410 23826 21422
rect 11678 21362 11730 21374
rect 22206 21362 22258 21374
rect 13570 21310 13582 21362
rect 13634 21310 13646 21362
rect 11678 21298 11730 21310
rect 22206 21298 22258 21310
rect 24782 21362 24834 21374
rect 24782 21298 24834 21310
rect 25790 21362 25842 21374
rect 25790 21298 25842 21310
rect 26014 21362 26066 21374
rect 26014 21298 26066 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 8318 21026 8370 21038
rect 19406 21026 19458 21038
rect 18498 20974 18510 21026
rect 18562 21023 18574 21026
rect 18834 21023 18846 21026
rect 18562 20977 18846 21023
rect 18562 20974 18574 20977
rect 18834 20974 18846 20977
rect 18898 20974 18910 21026
rect 8318 20962 8370 20974
rect 19406 20962 19458 20974
rect 20302 21026 20354 21038
rect 22318 21026 22370 21038
rect 20626 20974 20638 21026
rect 20690 20974 20702 21026
rect 20302 20962 20354 20974
rect 22318 20962 22370 20974
rect 4286 20914 4338 20926
rect 4286 20850 4338 20862
rect 7198 20914 7250 20926
rect 7198 20850 7250 20862
rect 12238 20914 12290 20926
rect 12238 20850 12290 20862
rect 12686 20914 12738 20926
rect 12686 20850 12738 20862
rect 18062 20914 18114 20926
rect 18062 20850 18114 20862
rect 18510 20914 18562 20926
rect 18510 20850 18562 20862
rect 21310 20914 21362 20926
rect 27458 20862 27470 20914
rect 27522 20862 27534 20914
rect 21310 20850 21362 20862
rect 2942 20802 2994 20814
rect 2942 20738 2994 20750
rect 3054 20802 3106 20814
rect 3054 20738 3106 20750
rect 3166 20802 3218 20814
rect 3726 20802 3778 20814
rect 6190 20802 6242 20814
rect 6862 20802 6914 20814
rect 3378 20750 3390 20802
rect 3442 20750 3454 20802
rect 5842 20750 5854 20802
rect 5906 20750 5918 20802
rect 6626 20750 6638 20802
rect 6690 20750 6702 20802
rect 3166 20738 3218 20750
rect 3726 20738 3778 20750
rect 6190 20738 6242 20750
rect 6862 20738 6914 20750
rect 7646 20802 7698 20814
rect 10446 20802 10498 20814
rect 8194 20750 8206 20802
rect 8258 20750 8270 20802
rect 9090 20750 9102 20802
rect 9154 20750 9166 20802
rect 9538 20750 9550 20802
rect 9602 20750 9614 20802
rect 7646 20738 7698 20750
rect 10446 20738 10498 20750
rect 11454 20802 11506 20814
rect 16158 20802 16210 20814
rect 19294 20802 19346 20814
rect 13794 20750 13806 20802
rect 13858 20750 13870 20802
rect 15138 20750 15150 20802
rect 15202 20750 15214 20802
rect 16930 20750 16942 20802
rect 16994 20750 17006 20802
rect 11454 20738 11506 20750
rect 16158 20738 16210 20750
rect 19294 20738 19346 20750
rect 20078 20802 20130 20814
rect 20078 20738 20130 20750
rect 21646 20802 21698 20814
rect 21646 20738 21698 20750
rect 22094 20802 22146 20814
rect 22094 20738 22146 20750
rect 22542 20802 22594 20814
rect 24770 20750 24782 20802
rect 24834 20750 24846 20802
rect 26786 20750 26798 20802
rect 26850 20750 26862 20802
rect 22542 20738 22594 20750
rect 1710 20690 1762 20702
rect 1710 20626 1762 20638
rect 2718 20690 2770 20702
rect 2718 20626 2770 20638
rect 5182 20690 5234 20702
rect 10222 20690 10274 20702
rect 22766 20690 22818 20702
rect 8978 20638 8990 20690
rect 9042 20638 9054 20690
rect 14354 20638 14366 20690
rect 14418 20638 14430 20690
rect 15922 20638 15934 20690
rect 15986 20638 15998 20690
rect 21410 20638 21422 20690
rect 21474 20638 21486 20690
rect 5182 20626 5234 20638
rect 10222 20626 10274 20638
rect 22766 20626 22818 20638
rect 22878 20690 22930 20702
rect 27358 20690 27410 20702
rect 24882 20638 24894 20690
rect 24946 20638 24958 20690
rect 22878 20626 22930 20638
rect 27358 20626 27410 20638
rect 2046 20578 2098 20590
rect 2046 20514 2098 20526
rect 6078 20578 6130 20590
rect 6078 20514 6130 20526
rect 7198 20578 7250 20590
rect 7198 20514 7250 20526
rect 9774 20578 9826 20590
rect 11566 20578 11618 20590
rect 10770 20526 10782 20578
rect 10834 20526 10846 20578
rect 9774 20514 9826 20526
rect 11566 20514 11618 20526
rect 11790 20578 11842 20590
rect 11790 20514 11842 20526
rect 18958 20578 19010 20590
rect 18958 20514 19010 20526
rect 19406 20578 19458 20590
rect 19406 20514 19458 20526
rect 23326 20578 23378 20590
rect 23326 20514 23378 20526
rect 24446 20578 24498 20590
rect 24446 20514 24498 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 2718 20242 2770 20254
rect 2718 20178 2770 20190
rect 3166 20242 3218 20254
rect 3166 20178 3218 20190
rect 3502 20242 3554 20254
rect 3502 20178 3554 20190
rect 8878 20242 8930 20254
rect 8878 20178 8930 20190
rect 10558 20242 10610 20254
rect 10558 20178 10610 20190
rect 12798 20242 12850 20254
rect 12798 20178 12850 20190
rect 16606 20242 16658 20254
rect 16606 20178 16658 20190
rect 17614 20242 17666 20254
rect 17614 20178 17666 20190
rect 20302 20242 20354 20254
rect 20302 20178 20354 20190
rect 1710 20130 1762 20142
rect 1710 20066 1762 20078
rect 2046 20130 2098 20142
rect 2046 20066 2098 20078
rect 5406 20130 5458 20142
rect 8766 20130 8818 20142
rect 7746 20078 7758 20130
rect 7810 20078 7822 20130
rect 5406 20066 5458 20078
rect 8766 20066 8818 20078
rect 10782 20130 10834 20142
rect 10782 20066 10834 20078
rect 11678 20130 11730 20142
rect 12462 20130 12514 20142
rect 16382 20130 16434 20142
rect 11890 20078 11902 20130
rect 11954 20078 11966 20130
rect 14354 20078 14366 20130
rect 14418 20078 14430 20130
rect 11678 20066 11730 20078
rect 12462 20066 12514 20078
rect 16382 20066 16434 20078
rect 21534 20130 21586 20142
rect 21534 20066 21586 20078
rect 21982 20130 22034 20142
rect 24782 20130 24834 20142
rect 23874 20078 23886 20130
rect 23938 20078 23950 20130
rect 24322 20078 24334 20130
rect 24386 20078 24398 20130
rect 26674 20078 26686 20130
rect 26738 20078 26750 20130
rect 27906 20078 27918 20130
rect 27970 20078 27982 20130
rect 21982 20066 22034 20078
rect 24782 20066 24834 20078
rect 2382 20018 2434 20030
rect 2382 19954 2434 19966
rect 4958 20018 5010 20030
rect 4958 19954 5010 19966
rect 5294 20018 5346 20030
rect 5294 19954 5346 19966
rect 5630 20018 5682 20030
rect 5630 19954 5682 19966
rect 7422 20018 7474 20030
rect 7422 19954 7474 19966
rect 7982 20018 8034 20030
rect 7982 19954 8034 19966
rect 8990 20018 9042 20030
rect 8990 19954 9042 19966
rect 10334 20018 10386 20030
rect 10334 19954 10386 19966
rect 10894 20018 10946 20030
rect 10894 19954 10946 19966
rect 11454 20018 11506 20030
rect 14590 20018 14642 20030
rect 12002 19966 12014 20018
rect 12066 19966 12078 20018
rect 13346 19966 13358 20018
rect 13410 19966 13422 20018
rect 13906 19966 13918 20018
rect 13970 19966 13982 20018
rect 11454 19954 11506 19966
rect 14590 19954 14642 19966
rect 14702 20018 14754 20030
rect 14702 19954 14754 19966
rect 14926 20018 14978 20030
rect 16270 20018 16322 20030
rect 17726 20018 17778 20030
rect 21310 20018 21362 20030
rect 15138 19966 15150 20018
rect 15202 19966 15214 20018
rect 16818 19966 16830 20018
rect 16882 19966 16894 20018
rect 18162 19966 18174 20018
rect 18226 19966 18238 20018
rect 18386 19966 18398 20018
rect 18450 19966 18462 20018
rect 14926 19954 14978 19966
rect 16270 19954 16322 19966
rect 17726 19954 17778 19966
rect 21310 19954 21362 19966
rect 21758 20018 21810 20030
rect 23538 19966 23550 20018
rect 23602 19966 23614 20018
rect 26114 19966 26126 20018
rect 26178 19966 26190 20018
rect 27682 19966 27694 20018
rect 27746 19966 27758 20018
rect 21758 19954 21810 19966
rect 4062 19906 4114 19918
rect 4062 19842 4114 19854
rect 4398 19906 4450 19918
rect 4398 19842 4450 19854
rect 6078 19906 6130 19918
rect 6078 19842 6130 19854
rect 6414 19906 6466 19918
rect 6414 19842 6466 19854
rect 6974 19906 7026 19918
rect 6974 19842 7026 19854
rect 8206 19906 8258 19918
rect 15710 19906 15762 19918
rect 20190 19906 20242 19918
rect 9874 19854 9886 19906
rect 9938 19854 9950 19906
rect 16706 19854 16718 19906
rect 16770 19854 16782 19906
rect 18722 19854 18734 19906
rect 18786 19854 18798 19906
rect 8206 19842 8258 19854
rect 15710 19842 15762 19854
rect 20190 19842 20242 19854
rect 21086 19906 21138 19918
rect 21086 19842 21138 19854
rect 22094 19906 22146 19918
rect 22094 19842 22146 19854
rect 22430 19906 22482 19918
rect 29474 19854 29486 19906
rect 29538 19854 29550 19906
rect 22430 19842 22482 19854
rect 7198 19794 7250 19806
rect 6066 19742 6078 19794
rect 6130 19791 6142 19794
rect 6514 19791 6526 19794
rect 6130 19745 6526 19791
rect 6130 19742 6142 19745
rect 6514 19742 6526 19745
rect 6578 19742 6590 19794
rect 7198 19730 7250 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 24110 19458 24162 19470
rect 15474 19406 15486 19458
rect 15538 19455 15550 19458
rect 15698 19455 15710 19458
rect 15538 19409 15710 19455
rect 15538 19406 15550 19409
rect 15698 19406 15710 19409
rect 15762 19406 15774 19458
rect 24110 19394 24162 19406
rect 25678 19458 25730 19470
rect 25678 19394 25730 19406
rect 8878 19346 8930 19358
rect 8878 19282 8930 19294
rect 12350 19346 12402 19358
rect 15374 19346 15426 19358
rect 20190 19346 20242 19358
rect 13570 19294 13582 19346
rect 13634 19294 13646 19346
rect 19394 19294 19406 19346
rect 19458 19294 19470 19346
rect 12350 19282 12402 19294
rect 15374 19282 15426 19294
rect 20190 19282 20242 19294
rect 22430 19346 22482 19358
rect 22430 19282 22482 19294
rect 23214 19346 23266 19358
rect 23214 19282 23266 19294
rect 11342 19234 11394 19246
rect 3042 19182 3054 19234
rect 3106 19182 3118 19234
rect 3490 19182 3502 19234
rect 3554 19182 3566 19234
rect 3938 19182 3950 19234
rect 4002 19182 4014 19234
rect 9538 19182 9550 19234
rect 9602 19182 9614 19234
rect 10994 19182 11006 19234
rect 11058 19182 11070 19234
rect 11342 19170 11394 19182
rect 11902 19234 11954 19246
rect 11902 19170 11954 19182
rect 12910 19234 12962 19246
rect 20078 19234 20130 19246
rect 24670 19234 24722 19246
rect 14018 19182 14030 19234
rect 14082 19182 14094 19234
rect 14802 19182 14814 19234
rect 14866 19182 14878 19234
rect 16370 19182 16382 19234
rect 16434 19182 16446 19234
rect 17826 19182 17838 19234
rect 17890 19182 17902 19234
rect 18498 19182 18510 19234
rect 18562 19182 18574 19234
rect 20626 19182 20638 19234
rect 20690 19182 20702 19234
rect 21410 19182 21422 19234
rect 21474 19182 21486 19234
rect 12910 19170 12962 19182
rect 20078 19170 20130 19182
rect 24670 19170 24722 19182
rect 24894 19234 24946 19246
rect 25218 19182 25230 19234
rect 25282 19182 25294 19234
rect 24894 19170 24946 19182
rect 1710 19122 1762 19134
rect 5742 19122 5794 19134
rect 14702 19122 14754 19134
rect 23998 19122 24050 19134
rect 2482 19070 2494 19122
rect 2546 19070 2558 19122
rect 4386 19070 4398 19122
rect 4450 19070 4462 19122
rect 10770 19070 10782 19122
rect 10834 19070 10846 19122
rect 13906 19070 13918 19122
rect 13970 19070 13982 19122
rect 19170 19070 19182 19122
rect 19234 19070 19246 19122
rect 21522 19070 21534 19122
rect 21586 19070 21598 19122
rect 21970 19070 21982 19122
rect 22034 19070 22046 19122
rect 1710 19058 1762 19070
rect 5742 19058 5794 19070
rect 14702 19058 14754 19070
rect 23998 19058 24050 19070
rect 25006 19122 25058 19134
rect 25006 19058 25058 19070
rect 2046 19010 2098 19022
rect 4846 19010 4898 19022
rect 4162 18958 4174 19010
rect 4226 18958 4238 19010
rect 2046 18946 2098 18958
rect 4846 18946 4898 18958
rect 9326 19010 9378 19022
rect 9326 18946 9378 18958
rect 9774 19010 9826 19022
rect 20302 19010 20354 19022
rect 10434 18958 10446 19010
rect 10498 18958 10510 19010
rect 9774 18946 9826 18958
rect 20302 18946 20354 18958
rect 24110 19010 24162 19022
rect 24110 18946 24162 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 2046 18674 2098 18686
rect 2046 18610 2098 18622
rect 3278 18674 3330 18686
rect 3278 18610 3330 18622
rect 10558 18674 10610 18686
rect 10558 18610 10610 18622
rect 15598 18674 15650 18686
rect 15598 18610 15650 18622
rect 16942 18674 16994 18686
rect 16942 18610 16994 18622
rect 18286 18674 18338 18686
rect 18286 18610 18338 18622
rect 19854 18674 19906 18686
rect 19854 18610 19906 18622
rect 20414 18674 20466 18686
rect 20414 18610 20466 18622
rect 20862 18674 20914 18686
rect 20862 18610 20914 18622
rect 22318 18674 22370 18686
rect 22318 18610 22370 18622
rect 23774 18674 23826 18686
rect 23774 18610 23826 18622
rect 2942 18562 2994 18574
rect 2942 18498 2994 18510
rect 3166 18562 3218 18574
rect 3166 18498 3218 18510
rect 4510 18562 4562 18574
rect 4510 18498 4562 18510
rect 5070 18562 5122 18574
rect 5070 18498 5122 18510
rect 7534 18562 7586 18574
rect 18174 18562 18226 18574
rect 11554 18510 11566 18562
rect 11618 18510 11630 18562
rect 14690 18510 14702 18562
rect 14754 18510 14766 18562
rect 7534 18498 7586 18510
rect 18174 18498 18226 18510
rect 20638 18562 20690 18574
rect 20638 18498 20690 18510
rect 22094 18562 22146 18574
rect 22094 18498 22146 18510
rect 1710 18450 1762 18462
rect 3838 18450 3890 18462
rect 7422 18450 7474 18462
rect 2706 18398 2718 18450
rect 2770 18398 2782 18450
rect 5842 18398 5854 18450
rect 5906 18398 5918 18450
rect 1710 18386 1762 18398
rect 3838 18386 3890 18398
rect 7422 18386 7474 18398
rect 8990 18450 9042 18462
rect 8990 18386 9042 18398
rect 9550 18450 9602 18462
rect 9550 18386 9602 18398
rect 10110 18450 10162 18462
rect 17950 18450 18002 18462
rect 10994 18398 11006 18450
rect 11058 18398 11070 18450
rect 12338 18398 12350 18450
rect 12402 18398 12414 18450
rect 14130 18398 14142 18450
rect 14194 18398 14206 18450
rect 10110 18386 10162 18398
rect 17950 18386 18002 18398
rect 19182 18450 19234 18462
rect 19182 18386 19234 18398
rect 19406 18450 19458 18462
rect 19406 18386 19458 18398
rect 19966 18450 20018 18462
rect 19966 18386 20018 18398
rect 20078 18450 20130 18462
rect 20078 18386 20130 18398
rect 21646 18450 21698 18462
rect 21646 18386 21698 18398
rect 21982 18450 22034 18462
rect 21982 18386 22034 18398
rect 22766 18450 22818 18462
rect 22766 18386 22818 18398
rect 23550 18450 23602 18462
rect 23550 18386 23602 18398
rect 23774 18450 23826 18462
rect 23774 18386 23826 18398
rect 24110 18450 24162 18462
rect 24110 18386 24162 18398
rect 3054 18338 3106 18350
rect 3054 18274 3106 18286
rect 5406 18338 5458 18350
rect 5406 18274 5458 18286
rect 15822 18338 15874 18350
rect 15822 18274 15874 18286
rect 20526 18338 20578 18350
rect 20526 18274 20578 18286
rect 22542 18338 22594 18350
rect 22542 18274 22594 18286
rect 7534 18226 7586 18238
rect 7534 18162 7586 18174
rect 16046 18226 16098 18238
rect 16046 18162 16098 18174
rect 16270 18226 16322 18238
rect 16270 18162 16322 18174
rect 16494 18226 16546 18238
rect 16494 18162 16546 18174
rect 18286 18226 18338 18238
rect 23090 18174 23102 18226
rect 23154 18174 23166 18226
rect 18286 18162 18338 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 18958 17890 19010 17902
rect 10546 17838 10558 17890
rect 10610 17887 10622 17890
rect 11218 17887 11230 17890
rect 10610 17841 11230 17887
rect 10610 17838 10622 17841
rect 11218 17838 11230 17841
rect 11282 17838 11294 17890
rect 18958 17826 19010 17838
rect 4622 17778 4674 17790
rect 13582 17778 13634 17790
rect 2258 17726 2270 17778
rect 2322 17726 2334 17778
rect 9874 17726 9886 17778
rect 9938 17726 9950 17778
rect 4622 17714 4674 17726
rect 13582 17714 13634 17726
rect 15710 17778 15762 17790
rect 17390 17778 17442 17790
rect 16706 17726 16718 17778
rect 16770 17726 16782 17778
rect 15710 17714 15762 17726
rect 17390 17714 17442 17726
rect 18622 17778 18674 17790
rect 18622 17714 18674 17726
rect 20638 17778 20690 17790
rect 23202 17726 23214 17778
rect 23266 17726 23278 17778
rect 20638 17714 20690 17726
rect 1822 17666 1874 17678
rect 1822 17602 1874 17614
rect 1934 17666 1986 17678
rect 11230 17666 11282 17678
rect 13470 17666 13522 17678
rect 14926 17666 14978 17678
rect 2370 17614 2382 17666
rect 2434 17614 2446 17666
rect 3266 17614 3278 17666
rect 3330 17614 3342 17666
rect 3714 17614 3726 17666
rect 3778 17614 3790 17666
rect 6850 17614 6862 17666
rect 6914 17614 6926 17666
rect 8754 17614 8766 17666
rect 8818 17614 8830 17666
rect 12002 17614 12014 17666
rect 12066 17614 12078 17666
rect 12338 17614 12350 17666
rect 12402 17614 12414 17666
rect 14018 17614 14030 17666
rect 14082 17614 14094 17666
rect 1934 17602 1986 17614
rect 11230 17602 11282 17614
rect 13470 17602 13522 17614
rect 14926 17602 14978 17614
rect 15374 17666 15426 17678
rect 15374 17602 15426 17614
rect 15598 17666 15650 17678
rect 16382 17666 16434 17678
rect 16146 17614 16158 17666
rect 16210 17614 16222 17666
rect 15598 17602 15650 17614
rect 16382 17602 16434 17614
rect 16606 17666 16658 17678
rect 16606 17602 16658 17614
rect 18846 17666 18898 17678
rect 21646 17666 21698 17678
rect 19394 17614 19406 17666
rect 19458 17614 19470 17666
rect 18846 17602 18898 17614
rect 21646 17602 21698 17614
rect 22206 17666 22258 17678
rect 22754 17614 22766 17666
rect 22818 17614 22830 17666
rect 24434 17614 24446 17666
rect 24498 17614 24510 17666
rect 25666 17614 25678 17666
rect 25730 17614 25742 17666
rect 22206 17602 22258 17614
rect 15150 17554 15202 17566
rect 2818 17502 2830 17554
rect 2882 17502 2894 17554
rect 8306 17502 8318 17554
rect 8370 17502 8382 17554
rect 9426 17502 9438 17554
rect 9490 17502 9502 17554
rect 12786 17502 12798 17554
rect 12850 17502 12862 17554
rect 15150 17490 15202 17502
rect 16718 17554 16770 17566
rect 19618 17502 19630 17554
rect 19682 17502 19694 17554
rect 20066 17502 20078 17554
rect 20130 17502 20142 17554
rect 22866 17502 22878 17554
rect 22930 17502 22942 17554
rect 16718 17490 16770 17502
rect 2158 17442 2210 17454
rect 10670 17442 10722 17454
rect 13694 17442 13746 17454
rect 3826 17390 3838 17442
rect 3890 17390 3902 17442
rect 4050 17390 4062 17442
rect 4114 17390 4126 17442
rect 11554 17390 11566 17442
rect 11618 17390 11630 17442
rect 12562 17390 12574 17442
rect 12626 17390 12638 17442
rect 2158 17378 2210 17390
rect 10670 17378 10722 17390
rect 13694 17378 13746 17390
rect 14590 17442 14642 17454
rect 14590 17378 14642 17390
rect 18062 17442 18114 17454
rect 18062 17378 18114 17390
rect 18958 17442 19010 17454
rect 18958 17378 19010 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 1934 17106 1986 17118
rect 4734 17106 4786 17118
rect 3826 17054 3838 17106
rect 3890 17054 3902 17106
rect 4050 17054 4062 17106
rect 4114 17054 4126 17106
rect 1934 17042 1986 17054
rect 4734 17042 4786 17054
rect 7198 17106 7250 17118
rect 7198 17042 7250 17054
rect 7310 17106 7362 17118
rect 7310 17042 7362 17054
rect 8654 17106 8706 17118
rect 10334 17106 10386 17118
rect 8978 17054 8990 17106
rect 9042 17054 9054 17106
rect 8654 17042 8706 17054
rect 10334 17042 10386 17054
rect 11566 17106 11618 17118
rect 11566 17042 11618 17054
rect 11678 17106 11730 17118
rect 11678 17042 11730 17054
rect 15374 17106 15426 17118
rect 15374 17042 15426 17054
rect 15598 17106 15650 17118
rect 15598 17042 15650 17054
rect 17502 17106 17554 17118
rect 17502 17042 17554 17054
rect 17614 17106 17666 17118
rect 17614 17042 17666 17054
rect 17726 17106 17778 17118
rect 19406 17106 19458 17118
rect 18834 17054 18846 17106
rect 18898 17054 18910 17106
rect 17726 17042 17778 17054
rect 19406 17042 19458 17054
rect 19630 17106 19682 17118
rect 19630 17042 19682 17054
rect 21198 17106 21250 17118
rect 21198 17042 21250 17054
rect 8094 16994 8146 17006
rect 2818 16942 2830 16994
rect 2882 16942 2894 16994
rect 7858 16942 7870 16994
rect 7922 16942 7934 16994
rect 8094 16930 8146 16942
rect 10558 16994 10610 17006
rect 10558 16930 10610 16942
rect 10670 16994 10722 17006
rect 10670 16930 10722 16942
rect 11230 16994 11282 17006
rect 11230 16930 11282 16942
rect 15822 16994 15874 17006
rect 15822 16930 15874 16942
rect 16382 16994 16434 17006
rect 16382 16930 16434 16942
rect 16830 16994 16882 17006
rect 16830 16930 16882 16942
rect 18510 16994 18562 17006
rect 18510 16930 18562 16942
rect 20526 16994 20578 17006
rect 21970 16942 21982 16994
rect 22034 16942 22046 16994
rect 22978 16942 22990 16994
rect 23042 16942 23054 16994
rect 20526 16930 20578 16942
rect 1822 16882 1874 16894
rect 1822 16818 1874 16830
rect 2158 16882 2210 16894
rect 2158 16818 2210 16830
rect 2270 16882 2322 16894
rect 4958 16882 5010 16894
rect 3154 16830 3166 16882
rect 3218 16830 3230 16882
rect 3602 16830 3614 16882
rect 3666 16830 3678 16882
rect 4498 16830 4510 16882
rect 4562 16830 4574 16882
rect 2270 16818 2322 16830
rect 4958 16818 5010 16830
rect 5070 16882 5122 16894
rect 8318 16882 8370 16894
rect 11790 16882 11842 16894
rect 7746 16830 7758 16882
rect 7810 16830 7822 16882
rect 9650 16830 9662 16882
rect 9714 16830 9726 16882
rect 5070 16818 5122 16830
rect 8318 16818 8370 16830
rect 11790 16818 11842 16830
rect 12238 16882 12290 16894
rect 12238 16818 12290 16830
rect 12462 16882 12514 16894
rect 12462 16818 12514 16830
rect 13022 16882 13074 16894
rect 13918 16882 13970 16894
rect 13458 16830 13470 16882
rect 13522 16830 13534 16882
rect 13022 16818 13074 16830
rect 13918 16818 13970 16830
rect 14254 16882 14306 16894
rect 14254 16818 14306 16830
rect 14590 16882 14642 16894
rect 14590 16818 14642 16830
rect 14702 16882 14754 16894
rect 14702 16818 14754 16830
rect 14926 16882 14978 16894
rect 16158 16882 16210 16894
rect 15138 16830 15150 16882
rect 15202 16830 15214 16882
rect 14926 16818 14978 16830
rect 16158 16818 16210 16830
rect 16606 16882 16658 16894
rect 16606 16818 16658 16830
rect 17838 16882 17890 16894
rect 17838 16818 17890 16830
rect 17950 16882 18002 16894
rect 20414 16882 20466 16894
rect 24558 16882 24610 16894
rect 19170 16830 19182 16882
rect 19234 16830 19246 16882
rect 19842 16830 19854 16882
rect 19906 16830 19918 16882
rect 20738 16830 20750 16882
rect 20802 16830 20814 16882
rect 22418 16830 22430 16882
rect 22482 16830 22494 16882
rect 17950 16818 18002 16830
rect 20414 16818 20466 16830
rect 24558 16818 24610 16830
rect 2046 16770 2098 16782
rect 2046 16706 2098 16718
rect 4846 16770 4898 16782
rect 19518 16770 19570 16782
rect 9986 16718 9998 16770
rect 10050 16718 10062 16770
rect 15250 16718 15262 16770
rect 15314 16718 15326 16770
rect 4846 16706 4898 16718
rect 19518 16706 19570 16718
rect 20190 16770 20242 16782
rect 24770 16718 24782 16770
rect 24834 16718 24846 16770
rect 20190 16706 20242 16718
rect 16270 16658 16322 16670
rect 16270 16594 16322 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 22430 16322 22482 16334
rect 14018 16270 14030 16322
rect 14082 16270 14094 16322
rect 22430 16258 22482 16270
rect 11006 16210 11058 16222
rect 4610 16158 4622 16210
rect 4674 16158 4686 16210
rect 11006 16146 11058 16158
rect 13470 16210 13522 16222
rect 13470 16146 13522 16158
rect 13694 16210 13746 16222
rect 19406 16210 19458 16222
rect 15250 16158 15262 16210
rect 15314 16158 15326 16210
rect 18610 16158 18622 16210
rect 18674 16158 18686 16210
rect 13694 16146 13746 16158
rect 19406 16146 19458 16158
rect 20414 16210 20466 16222
rect 20414 16146 20466 16158
rect 21646 16210 21698 16222
rect 24322 16158 24334 16210
rect 24386 16158 24398 16210
rect 21646 16146 21698 16158
rect 1710 16098 1762 16110
rect 5070 16098 5122 16110
rect 7870 16098 7922 16110
rect 10446 16098 10498 16110
rect 11790 16098 11842 16110
rect 3266 16046 3278 16098
rect 3330 16046 3342 16098
rect 3602 16046 3614 16098
rect 3666 16046 3678 16098
rect 5842 16046 5854 16098
rect 5906 16046 5918 16098
rect 9538 16046 9550 16098
rect 9602 16046 9614 16098
rect 11330 16046 11342 16098
rect 11394 16046 11406 16098
rect 1710 16034 1762 16046
rect 5070 16034 5122 16046
rect 7870 16034 7922 16046
rect 10446 16034 10498 16046
rect 11790 16034 11842 16046
rect 12238 16098 12290 16110
rect 12238 16034 12290 16046
rect 12462 16098 12514 16110
rect 12462 16034 12514 16046
rect 14926 16098 14978 16110
rect 15934 16098 15986 16110
rect 17502 16098 17554 16110
rect 15698 16046 15710 16098
rect 15762 16046 15774 16098
rect 16370 16046 16382 16098
rect 16434 16046 16446 16098
rect 17042 16046 17054 16098
rect 17106 16046 17118 16098
rect 14926 16034 14978 16046
rect 15934 16034 15986 16046
rect 17502 16034 17554 16046
rect 17614 16098 17666 16110
rect 20526 16098 20578 16110
rect 21534 16098 21586 16110
rect 18050 16046 18062 16098
rect 18114 16046 18126 16098
rect 19058 16046 19070 16098
rect 19122 16046 19134 16098
rect 19730 16046 19742 16098
rect 19794 16046 19806 16098
rect 20738 16046 20750 16098
rect 20802 16046 20814 16098
rect 21298 16046 21310 16098
rect 21362 16046 21374 16098
rect 17614 16034 17666 16046
rect 20526 16034 20578 16046
rect 21534 16034 21586 16046
rect 21758 16098 21810 16110
rect 21758 16034 21810 16046
rect 21870 16098 21922 16110
rect 21870 16034 21922 16046
rect 22542 16098 22594 16110
rect 23090 16046 23102 16098
rect 23154 16046 23166 16098
rect 24658 16046 24670 16098
rect 24722 16046 24734 16098
rect 26002 16046 26014 16098
rect 26066 16046 26078 16098
rect 22542 16034 22594 16046
rect 2046 15986 2098 15998
rect 8206 15986 8258 15998
rect 9886 15986 9938 15998
rect 2818 15934 2830 15986
rect 2882 15934 2894 15986
rect 5618 15934 5630 15986
rect 5682 15934 5694 15986
rect 8978 15934 8990 15986
rect 9042 15934 9054 15986
rect 9202 15934 9214 15986
rect 9266 15934 9278 15986
rect 2046 15922 2098 15934
rect 8206 15922 8258 15934
rect 9886 15922 9938 15934
rect 9998 15986 10050 15998
rect 9998 15922 10050 15934
rect 10222 15986 10274 15998
rect 10222 15922 10274 15934
rect 14702 15986 14754 15998
rect 14702 15922 14754 15934
rect 16158 15986 16210 15998
rect 18274 15934 18286 15986
rect 18338 15934 18350 15986
rect 23202 15934 23214 15986
rect 23266 15934 23278 15986
rect 16158 15922 16210 15934
rect 7982 15874 8034 15886
rect 11678 15874 11730 15886
rect 3826 15822 3838 15874
rect 3890 15822 3902 15874
rect 4050 15822 4062 15874
rect 4114 15822 4126 15874
rect 8530 15822 8542 15874
rect 8594 15822 8606 15874
rect 7982 15810 8034 15822
rect 11678 15810 11730 15822
rect 11902 15874 11954 15886
rect 15150 15874 15202 15886
rect 12786 15822 12798 15874
rect 12850 15822 12862 15874
rect 11902 15810 11954 15822
rect 15150 15810 15202 15822
rect 15262 15874 15314 15886
rect 15262 15810 15314 15822
rect 16046 15874 16098 15886
rect 16046 15810 16098 15822
rect 17278 15874 17330 15886
rect 17278 15810 17330 15822
rect 17390 15874 17442 15886
rect 17390 15810 17442 15822
rect 19294 15874 19346 15886
rect 19294 15810 19346 15822
rect 19518 15874 19570 15886
rect 19518 15810 19570 15822
rect 20190 15874 20242 15886
rect 20190 15810 20242 15822
rect 20302 15874 20354 15886
rect 20302 15810 20354 15822
rect 22430 15874 22482 15886
rect 22430 15810 22482 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 2046 15538 2098 15550
rect 2046 15474 2098 15486
rect 2718 15538 2770 15550
rect 2718 15474 2770 15486
rect 3278 15538 3330 15550
rect 8990 15538 9042 15550
rect 13918 15538 13970 15550
rect 8642 15486 8654 15538
rect 8706 15486 8718 15538
rect 10882 15486 10894 15538
rect 10946 15486 10958 15538
rect 13234 15486 13246 15538
rect 13298 15486 13310 15538
rect 3278 15474 3330 15486
rect 8990 15474 9042 15486
rect 13918 15474 13970 15486
rect 16046 15538 16098 15550
rect 16046 15474 16098 15486
rect 16382 15538 16434 15550
rect 16382 15474 16434 15486
rect 18734 15538 18786 15550
rect 18734 15474 18786 15486
rect 19406 15538 19458 15550
rect 22094 15538 22146 15550
rect 21410 15486 21422 15538
rect 21474 15486 21486 15538
rect 19406 15474 19458 15486
rect 22094 15474 22146 15486
rect 22766 15538 22818 15550
rect 22766 15474 22818 15486
rect 1710 15426 1762 15438
rect 1710 15362 1762 15374
rect 3502 15426 3554 15438
rect 11230 15426 11282 15438
rect 4274 15374 4286 15426
rect 4338 15374 4350 15426
rect 6178 15374 6190 15426
rect 6242 15374 6254 15426
rect 6962 15374 6974 15426
rect 7026 15374 7038 15426
rect 3502 15362 3554 15374
rect 11230 15362 11282 15374
rect 12910 15426 12962 15438
rect 12910 15362 12962 15374
rect 14814 15426 14866 15438
rect 23214 15426 23266 15438
rect 17378 15374 17390 15426
rect 17442 15374 17454 15426
rect 19730 15374 19742 15426
rect 19794 15374 19806 15426
rect 21634 15374 21646 15426
rect 21698 15374 21710 15426
rect 14814 15362 14866 15374
rect 23214 15362 23266 15374
rect 2382 15314 2434 15326
rect 2382 15250 2434 15262
rect 3166 15314 3218 15326
rect 9550 15314 9602 15326
rect 12574 15314 12626 15326
rect 14478 15314 14530 15326
rect 3938 15262 3950 15314
rect 4002 15262 4014 15314
rect 6066 15262 6078 15314
rect 6130 15262 6142 15314
rect 7186 15262 7198 15314
rect 7250 15262 7262 15314
rect 9986 15262 9998 15314
rect 10050 15262 10062 15314
rect 10658 15262 10670 15314
rect 10722 15262 10734 15314
rect 13458 15262 13470 15314
rect 13522 15262 13534 15314
rect 3166 15250 3218 15262
rect 9550 15250 9602 15262
rect 12574 15250 12626 15262
rect 14478 15250 14530 15262
rect 15374 15314 15426 15326
rect 15374 15250 15426 15262
rect 15934 15314 15986 15326
rect 15934 15250 15986 15262
rect 16158 15314 16210 15326
rect 16158 15250 16210 15262
rect 16270 15314 16322 15326
rect 17490 15262 17502 15314
rect 17554 15262 17566 15314
rect 18162 15262 18174 15314
rect 18226 15262 18238 15314
rect 18610 15262 18622 15314
rect 18674 15262 18686 15314
rect 20290 15262 20302 15314
rect 20354 15262 20366 15314
rect 20514 15262 20526 15314
rect 20578 15262 20590 15314
rect 21186 15262 21198 15314
rect 21250 15262 21262 15314
rect 16270 15250 16322 15262
rect 11666 15150 11678 15202
rect 11730 15150 11742 15202
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 3838 14754 3890 14766
rect 21982 14754 22034 14766
rect 2258 14702 2270 14754
rect 2322 14751 2334 14754
rect 2706 14751 2718 14754
rect 2322 14705 2718 14751
rect 2322 14702 2334 14705
rect 2706 14702 2718 14705
rect 2770 14702 2782 14754
rect 10770 14702 10782 14754
rect 10834 14751 10846 14754
rect 11666 14751 11678 14754
rect 10834 14705 11678 14751
rect 10834 14702 10846 14705
rect 11666 14702 11678 14705
rect 11730 14702 11742 14754
rect 3838 14690 3890 14702
rect 21982 14690 22034 14702
rect 2494 14642 2546 14654
rect 2494 14578 2546 14590
rect 2942 14642 2994 14654
rect 2942 14578 2994 14590
rect 9326 14642 9378 14654
rect 9326 14578 9378 14590
rect 10222 14642 10274 14654
rect 10222 14578 10274 14590
rect 10782 14642 10834 14654
rect 10782 14578 10834 14590
rect 11230 14642 11282 14654
rect 11230 14578 11282 14590
rect 11678 14642 11730 14654
rect 11678 14578 11730 14590
rect 13022 14642 13074 14654
rect 16158 14642 16210 14654
rect 14690 14590 14702 14642
rect 14754 14590 14766 14642
rect 13022 14578 13074 14590
rect 16158 14578 16210 14590
rect 16494 14642 16546 14654
rect 20862 14642 20914 14654
rect 18162 14590 18174 14642
rect 18226 14590 18238 14642
rect 18610 14590 18622 14642
rect 18674 14590 18686 14642
rect 16494 14578 16546 14590
rect 20862 14578 20914 14590
rect 21422 14642 21474 14654
rect 21422 14578 21474 14590
rect 22542 14642 22594 14654
rect 22542 14578 22594 14590
rect 3726 14530 3778 14542
rect 14030 14530 14082 14542
rect 19518 14530 19570 14542
rect 13570 14478 13582 14530
rect 13634 14478 13646 14530
rect 15362 14478 15374 14530
rect 15426 14478 15438 14530
rect 16930 14478 16942 14530
rect 16994 14478 17006 14530
rect 17602 14478 17614 14530
rect 17666 14478 17678 14530
rect 18946 14478 18958 14530
rect 19010 14478 19022 14530
rect 3726 14466 3778 14478
rect 14030 14466 14082 14478
rect 19518 14466 19570 14478
rect 22094 14530 22146 14542
rect 22094 14466 22146 14478
rect 1710 14418 1762 14430
rect 1710 14354 1762 14366
rect 2046 14418 2098 14430
rect 21982 14418 22034 14430
rect 17490 14366 17502 14418
rect 17554 14366 17566 14418
rect 2046 14354 2098 14366
rect 21982 14354 22034 14366
rect 3390 14306 3442 14318
rect 3390 14242 3442 14254
rect 3838 14306 3890 14318
rect 3838 14242 3890 14254
rect 9886 14306 9938 14318
rect 9886 14242 9938 14254
rect 12238 14306 12290 14318
rect 12238 14242 12290 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 2046 13970 2098 13982
rect 2046 13906 2098 13918
rect 2494 13970 2546 13982
rect 2494 13906 2546 13918
rect 10334 13970 10386 13982
rect 10334 13906 10386 13918
rect 11006 13970 11058 13982
rect 15150 13970 15202 13982
rect 14018 13918 14030 13970
rect 14082 13918 14094 13970
rect 14802 13918 14814 13970
rect 14866 13918 14878 13970
rect 11006 13906 11058 13918
rect 15150 13906 15202 13918
rect 15710 13970 15762 13982
rect 15710 13906 15762 13918
rect 16270 13970 16322 13982
rect 16270 13906 16322 13918
rect 18062 13970 18114 13982
rect 18062 13906 18114 13918
rect 18510 13970 18562 13982
rect 18510 13906 18562 13918
rect 18958 13970 19010 13982
rect 18958 13906 19010 13918
rect 12798 13858 12850 13870
rect 12798 13794 12850 13806
rect 13246 13858 13298 13870
rect 13246 13794 13298 13806
rect 13694 13858 13746 13870
rect 13694 13794 13746 13806
rect 1710 13746 1762 13758
rect 1710 13682 1762 13694
rect 2942 13634 2994 13646
rect 2942 13570 2994 13582
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 2034 12798 2046 12850
rect 2098 12798 2110 12850
rect 1710 12738 1762 12750
rect 1710 12674 1762 12686
rect 2494 12738 2546 12750
rect 2494 12674 2546 12686
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 2046 12402 2098 12414
rect 2046 12338 2098 12350
rect 1710 12178 1762 12190
rect 1710 12114 1762 12126
rect 2494 12066 2546 12078
rect 2494 12002 2546 12014
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1710 11282 1762 11294
rect 1710 11218 1762 11230
rect 2046 11282 2098 11294
rect 2046 11218 2098 11230
rect 2494 11170 2546 11182
rect 2494 11106 2546 11118
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1922 9774 1934 9826
rect 1986 9774 1998 9826
rect 1710 9714 1762 9726
rect 1710 9650 1762 9662
rect 2494 9714 2546 9726
rect 2494 9650 2546 9662
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 2034 9214 2046 9266
rect 2098 9214 2110 9266
rect 1710 9042 1762 9054
rect 1710 8978 1762 8990
rect 2494 8930 2546 8942
rect 2494 8866 2546 8878
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1710 8146 1762 8158
rect 1710 8082 1762 8094
rect 2046 8146 2098 8158
rect 2046 8082 2098 8094
rect 2494 8034 2546 8046
rect 2494 7970 2546 7982
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 2046 7698 2098 7710
rect 2046 7634 2098 7646
rect 1710 7474 1762 7486
rect 1710 7410 1762 7422
rect 2494 7362 2546 7374
rect 2494 7298 2546 7310
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1710 6578 1762 6590
rect 1710 6514 1762 6526
rect 2046 6578 2098 6590
rect 2046 6514 2098 6526
rect 2494 6466 2546 6478
rect 2494 6402 2546 6414
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 2034 6078 2046 6130
rect 2098 6078 2110 6130
rect 1710 5906 1762 5918
rect 1710 5842 1762 5854
rect 2494 5794 2546 5806
rect 2494 5730 2546 5742
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 2494 5122 2546 5134
rect 2494 5058 2546 5070
rect 1710 5010 1762 5022
rect 1710 4946 1762 4958
rect 2046 5010 2098 5022
rect 2046 4946 2098 4958
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 1710 3442 1762 3454
rect 1710 3378 1762 3390
rect 2046 3442 2098 3454
rect 2046 3378 2098 3390
rect 2494 3442 2546 3454
rect 2494 3378 2546 3390
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 3614 38558 3666 38610
rect 6750 38558 6802 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 6862 38222 6914 38274
rect 7086 38222 7138 38274
rect 8094 38222 8146 38274
rect 17166 38222 17218 38274
rect 25566 38222 25618 38274
rect 30046 38222 30098 38274
rect 33854 38222 33906 38274
rect 37326 38222 37378 38274
rect 7758 38110 7810 38162
rect 8878 38110 8930 38162
rect 9886 38110 9938 38162
rect 11006 38110 11058 38162
rect 11790 38110 11842 38162
rect 1822 37998 1874 38050
rect 3390 37998 3442 38050
rect 4286 37998 4338 38050
rect 5966 37998 6018 38050
rect 7310 37998 7362 38050
rect 9438 37998 9490 38050
rect 12350 37998 12402 38050
rect 13134 37998 13186 38050
rect 14254 37998 14306 38050
rect 15038 37998 15090 38050
rect 19518 37998 19570 38050
rect 19966 37998 20018 38050
rect 24558 37998 24610 38050
rect 29038 37998 29090 38050
rect 32846 37998 32898 38050
rect 36430 37998 36482 38050
rect 2382 37886 2434 37938
rect 3614 37886 3666 37938
rect 4958 37886 5010 37938
rect 6526 37886 6578 37938
rect 6750 37886 6802 37938
rect 8206 37886 8258 37938
rect 13358 37886 13410 37938
rect 13470 37886 13522 37938
rect 21310 37886 21362 37938
rect 2046 37774 2098 37826
rect 2718 37774 2770 37826
rect 3950 37774 4002 37826
rect 4622 37774 4674 37826
rect 6190 37774 6242 37826
rect 10446 37774 10498 37826
rect 13918 37774 13970 37826
rect 14590 37774 14642 37826
rect 20974 37774 21026 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 3614 37438 3666 37490
rect 14702 37438 14754 37490
rect 23662 37438 23714 37490
rect 27246 37438 27298 37490
rect 6750 37326 6802 37378
rect 10222 37326 10274 37378
rect 11118 37326 11170 37378
rect 25902 37326 25954 37378
rect 39454 37326 39506 37378
rect 2270 37214 2322 37266
rect 4286 37214 4338 37266
rect 5406 37214 5458 37266
rect 5966 37214 6018 37266
rect 6414 37214 6466 37266
rect 7310 37214 7362 37266
rect 8206 37214 8258 37266
rect 10782 37214 10834 37266
rect 12686 37214 12738 37266
rect 13470 37214 13522 37266
rect 13694 37214 13746 37266
rect 21646 37214 21698 37266
rect 23326 37214 23378 37266
rect 25678 37214 25730 37266
rect 26238 37214 26290 37266
rect 37662 37214 37714 37266
rect 1822 37102 1874 37154
rect 2718 37102 2770 37154
rect 3166 37102 3218 37154
rect 6862 37102 6914 37154
rect 7758 37102 7810 37154
rect 8542 37102 8594 37154
rect 11342 37102 11394 37154
rect 14142 37102 14194 37154
rect 15262 37102 15314 37154
rect 19742 37102 19794 37154
rect 35982 37102 36034 37154
rect 37438 37102 37490 37154
rect 13918 36990 13970 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 3838 36654 3890 36706
rect 2494 36542 2546 36594
rect 3502 36542 3554 36594
rect 4062 36542 4114 36594
rect 11566 36542 11618 36594
rect 14254 36542 14306 36594
rect 15262 36542 15314 36594
rect 16718 36542 16770 36594
rect 2606 36430 2658 36482
rect 2942 36430 2994 36482
rect 4174 36430 4226 36482
rect 4846 36430 4898 36482
rect 5742 36430 5794 36482
rect 5854 36430 5906 36482
rect 5966 36430 6018 36482
rect 6974 36430 7026 36482
rect 9998 36430 10050 36482
rect 12238 36430 12290 36482
rect 12798 36430 12850 36482
rect 12910 36430 12962 36482
rect 13806 36430 13858 36482
rect 14030 36430 14082 36482
rect 15150 36430 15202 36482
rect 16382 36430 16434 36482
rect 17278 36430 17330 36482
rect 5070 36318 5122 36370
rect 8542 36318 8594 36370
rect 11006 36318 11058 36370
rect 15262 36318 15314 36370
rect 1710 36206 1762 36258
rect 2046 36206 2098 36258
rect 6414 36206 6466 36258
rect 7646 36206 7698 36258
rect 8094 36206 8146 36258
rect 14702 36206 14754 36258
rect 17502 36206 17554 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 6862 35870 6914 35922
rect 2046 35758 2098 35810
rect 2382 35758 2434 35810
rect 4398 35758 4450 35810
rect 4846 35758 4898 35810
rect 6302 35758 6354 35810
rect 7310 35758 7362 35810
rect 10110 35758 10162 35810
rect 13694 35758 13746 35810
rect 16158 35758 16210 35810
rect 1822 35646 1874 35698
rect 2606 35646 2658 35698
rect 5294 35646 5346 35698
rect 6414 35646 6466 35698
rect 11006 35646 11058 35698
rect 11230 35646 11282 35698
rect 12574 35646 12626 35698
rect 14590 35646 14642 35698
rect 17390 35646 17442 35698
rect 3166 35534 3218 35586
rect 3614 35534 3666 35586
rect 6078 35534 6130 35586
rect 11678 35534 11730 35586
rect 14030 35534 14082 35586
rect 17838 35534 17890 35586
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 4286 34974 4338 35026
rect 14254 34974 14306 35026
rect 3390 34862 3442 34914
rect 7982 34862 8034 34914
rect 8206 34862 8258 34914
rect 8318 34862 8370 34914
rect 8766 34862 8818 34914
rect 10782 34862 10834 34914
rect 12798 34862 12850 34914
rect 16046 34862 16098 34914
rect 16382 34862 16434 34914
rect 16942 34862 16994 34914
rect 2942 34750 2994 34802
rect 4734 34750 4786 34802
rect 4846 34750 4898 34802
rect 6190 34750 6242 34802
rect 6526 34750 6578 34802
rect 6862 34750 6914 34802
rect 10222 34750 10274 34802
rect 10894 34750 10946 34802
rect 12910 34750 12962 34802
rect 15486 34750 15538 34802
rect 1934 34638 1986 34690
rect 2270 34638 2322 34690
rect 2606 34638 2658 34690
rect 3838 34638 3890 34690
rect 5070 34638 5122 34690
rect 5630 34638 5682 34690
rect 13694 34638 13746 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 7870 34302 7922 34354
rect 2270 34190 2322 34242
rect 4286 34190 4338 34242
rect 6750 34190 6802 34242
rect 8878 34190 8930 34242
rect 11790 34190 11842 34242
rect 11902 34190 11954 34242
rect 12014 34190 12066 34242
rect 16830 34190 16882 34242
rect 18062 34190 18114 34242
rect 19966 34190 20018 34242
rect 2046 34078 2098 34130
rect 2606 34078 2658 34130
rect 5854 34078 5906 34130
rect 6190 34078 6242 34130
rect 8430 34078 8482 34130
rect 9550 34078 9602 34130
rect 9774 34078 9826 34130
rect 13806 34078 13858 34130
rect 14702 34078 14754 34130
rect 16046 34078 16098 34130
rect 16494 34078 16546 34130
rect 17838 34078 17890 34130
rect 18174 34078 18226 34130
rect 3726 33966 3778 34018
rect 8766 33966 8818 34018
rect 12462 33966 12514 34018
rect 13582 33966 13634 34018
rect 15262 33966 15314 34018
rect 15710 33966 15762 34018
rect 18622 33966 18674 34018
rect 10110 33854 10162 33906
rect 14142 33854 14194 33906
rect 19854 33854 19906 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 17614 33518 17666 33570
rect 3502 33406 3554 33458
rect 4846 33406 4898 33458
rect 7086 33406 7138 33458
rect 9214 33406 9266 33458
rect 15598 33406 15650 33458
rect 2270 33294 2322 33346
rect 2830 33294 2882 33346
rect 4398 33294 4450 33346
rect 4734 33294 4786 33346
rect 5630 33294 5682 33346
rect 6862 33294 6914 33346
rect 6974 33294 7026 33346
rect 8654 33294 8706 33346
rect 10222 33294 10274 33346
rect 11790 33294 11842 33346
rect 13582 33294 13634 33346
rect 14030 33294 14082 33346
rect 15038 33294 15090 33346
rect 16046 33294 16098 33346
rect 16270 33294 16322 33346
rect 16494 33294 16546 33346
rect 16718 33294 16770 33346
rect 17054 33294 17106 33346
rect 17726 33294 17778 33346
rect 18062 33294 18114 33346
rect 19854 33294 19906 33346
rect 2494 33182 2546 33234
rect 2942 33182 2994 33234
rect 10334 33182 10386 33234
rect 11454 33182 11506 33234
rect 15262 33182 15314 33234
rect 18286 33182 18338 33234
rect 18398 33182 18450 33234
rect 19182 33182 19234 33234
rect 20078 33182 20130 33234
rect 20302 33182 20354 33234
rect 1822 33070 1874 33122
rect 5182 33070 5234 33122
rect 5966 33070 6018 33122
rect 7758 33070 7810 33122
rect 12014 33070 12066 33122
rect 14702 33070 14754 33122
rect 15486 33070 15538 33122
rect 15598 33070 15650 33122
rect 16382 33070 16434 33122
rect 17278 33070 17330 33122
rect 17502 33070 17554 33122
rect 18846 33070 18898 33122
rect 19518 33070 19570 33122
rect 20638 33070 20690 33122
rect 23438 33070 23490 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 8318 32734 8370 32786
rect 12238 32734 12290 32786
rect 12462 32734 12514 32786
rect 13582 32734 13634 32786
rect 19406 32734 19458 32786
rect 2494 32622 2546 32674
rect 2830 32622 2882 32674
rect 5294 32622 5346 32674
rect 7870 32622 7922 32674
rect 10782 32622 10834 32674
rect 12126 32622 12178 32674
rect 15598 32622 15650 32674
rect 16830 32622 16882 32674
rect 17390 32622 17442 32674
rect 21310 32622 21362 32674
rect 23102 32622 23154 32674
rect 2270 32510 2322 32562
rect 3054 32510 3106 32562
rect 4286 32510 4338 32562
rect 6302 32510 6354 32562
rect 6750 32510 6802 32562
rect 9998 32510 10050 32562
rect 12798 32510 12850 32562
rect 14142 32510 14194 32562
rect 15374 32510 15426 32562
rect 19854 32510 19906 32562
rect 20974 32510 21026 32562
rect 21198 32510 21250 32562
rect 23438 32510 23490 32562
rect 1822 32398 1874 32450
rect 3838 32398 3890 32450
rect 10446 32398 10498 32450
rect 17838 32398 17890 32450
rect 18958 32398 19010 32450
rect 20078 32398 20130 32450
rect 20526 32398 20578 32450
rect 22206 32398 22258 32450
rect 22766 32398 22818 32450
rect 23886 32398 23938 32450
rect 24334 32398 24386 32450
rect 3390 32286 3442 32338
rect 11006 32286 11058 32338
rect 11230 32286 11282 32338
rect 11454 32286 11506 32338
rect 11902 32286 11954 32338
rect 16270 32286 16322 32338
rect 16606 32286 16658 32338
rect 19742 32286 19794 32338
rect 20302 32286 20354 32338
rect 21758 32286 21810 32338
rect 23774 32286 23826 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 2270 31950 2322 32002
rect 10110 31950 10162 32002
rect 2046 31838 2098 31890
rect 3502 31838 3554 31890
rect 4846 31838 4898 31890
rect 6638 31838 6690 31890
rect 10334 31838 10386 31890
rect 11118 31838 11170 31890
rect 16270 31838 16322 31890
rect 21310 31838 21362 31890
rect 22542 31838 22594 31890
rect 24110 31838 24162 31890
rect 4286 31726 4338 31778
rect 4398 31726 4450 31778
rect 5182 31726 5234 31778
rect 6190 31726 6242 31778
rect 6414 31726 6466 31778
rect 7422 31726 7474 31778
rect 7758 31726 7810 31778
rect 7870 31726 7922 31778
rect 8654 31726 8706 31778
rect 8878 31726 8930 31778
rect 13918 31726 13970 31778
rect 15374 31726 15426 31778
rect 15710 31726 15762 31778
rect 16606 31726 16658 31778
rect 16942 31726 16994 31778
rect 17502 31726 17554 31778
rect 21534 31726 21586 31778
rect 22318 31726 22370 31778
rect 23102 31726 23154 31778
rect 23886 31726 23938 31778
rect 7086 31614 7138 31666
rect 9438 31614 9490 31666
rect 15150 31614 15202 31666
rect 15598 31614 15650 31666
rect 16046 31614 16098 31666
rect 2606 31502 2658 31554
rect 2942 31502 2994 31554
rect 9774 31502 9826 31554
rect 10670 31502 10722 31554
rect 11678 31502 11730 31554
rect 12014 31502 12066 31554
rect 12350 31502 12402 31554
rect 14254 31502 14306 31554
rect 16494 31502 16546 31554
rect 17950 31502 18002 31554
rect 21870 31502 21922 31554
rect 22654 31502 22706 31554
rect 22878 31502 22930 31554
rect 23438 31502 23490 31554
rect 23662 31502 23714 31554
rect 23774 31502 23826 31554
rect 24222 31502 24274 31554
rect 24446 31502 24498 31554
rect 24894 31502 24946 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 7870 31166 7922 31218
rect 13022 31166 13074 31218
rect 15598 31166 15650 31218
rect 2046 31054 2098 31106
rect 2718 31054 2770 31106
rect 16494 31110 16546 31162
rect 20974 31166 21026 31218
rect 22542 31166 22594 31218
rect 25454 31166 25506 31218
rect 3166 31054 3218 31106
rect 11342 31054 11394 31106
rect 13246 31054 13298 31106
rect 15150 31054 15202 31106
rect 15934 31054 15986 31106
rect 16606 31054 16658 31106
rect 21310 31054 21362 31106
rect 21422 31054 21474 31106
rect 23438 31054 23490 31106
rect 23998 31054 24050 31106
rect 25230 31054 25282 31106
rect 1710 30942 1762 30994
rect 2494 30942 2546 30994
rect 4286 30942 4338 30994
rect 4734 30942 4786 30994
rect 5630 30942 5682 30994
rect 6078 30942 6130 30994
rect 6526 30942 6578 30994
rect 6862 30942 6914 30994
rect 10222 30942 10274 30994
rect 11678 30942 11730 30994
rect 12126 30942 12178 30994
rect 12910 30942 12962 30994
rect 13694 30942 13746 30994
rect 18622 30942 18674 30994
rect 21982 30942 22034 30994
rect 22206 30942 22258 30994
rect 23102 30942 23154 30994
rect 3838 30830 3890 30882
rect 5182 30830 5234 30882
rect 8430 30830 8482 30882
rect 9998 30830 10050 30882
rect 14366 30830 14418 30882
rect 14702 30830 14754 30882
rect 18398 30830 18450 30882
rect 20526 30830 20578 30882
rect 24334 30830 24386 30882
rect 25342 30830 25394 30882
rect 3054 30718 3106 30770
rect 10446 30718 10498 30770
rect 10782 30718 10834 30770
rect 14142 30718 14194 30770
rect 14366 30718 14418 30770
rect 16606 30718 16658 30770
rect 18958 30718 19010 30770
rect 21422 30718 21474 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 8654 30382 8706 30434
rect 8990 30382 9042 30434
rect 24222 30382 24274 30434
rect 3054 30270 3106 30322
rect 3166 30270 3218 30322
rect 6414 30270 6466 30322
rect 8766 30270 8818 30322
rect 9998 30270 10050 30322
rect 1710 30158 1762 30210
rect 3614 30158 3666 30210
rect 5070 30158 5122 30210
rect 6638 30158 6690 30210
rect 9102 30158 9154 30210
rect 9886 30158 9938 30210
rect 11454 30158 11506 30210
rect 14142 30158 14194 30210
rect 15262 30158 15314 30210
rect 15598 30158 15650 30210
rect 15934 30158 15986 30210
rect 18510 30158 18562 30210
rect 19854 30158 19906 30210
rect 23998 30158 24050 30210
rect 2046 30046 2098 30098
rect 4062 30046 4114 30098
rect 4510 30046 4562 30098
rect 7198 30046 7250 30098
rect 11902 30046 11954 30098
rect 12350 30046 12402 30098
rect 12462 30046 12514 30098
rect 12574 30046 12626 30098
rect 17390 30046 17442 30098
rect 19406 30046 19458 30098
rect 22990 30046 23042 30098
rect 2830 29934 2882 29986
rect 8094 29934 8146 29986
rect 9550 29934 9602 29986
rect 10670 29934 10722 29986
rect 13582 29934 13634 29986
rect 18846 29934 18898 29986
rect 23102 29934 23154 29986
rect 23326 29934 23378 29986
rect 24558 29934 24610 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 2942 29598 2994 29650
rect 8766 29598 8818 29650
rect 14366 29598 14418 29650
rect 15038 29598 15090 29650
rect 15262 29598 15314 29650
rect 16494 29598 16546 29650
rect 18286 29598 18338 29650
rect 18510 29598 18562 29650
rect 18622 29598 18674 29650
rect 2046 29486 2098 29538
rect 4958 29486 5010 29538
rect 6974 29486 7026 29538
rect 8878 29486 8930 29538
rect 19070 29486 19122 29538
rect 21422 29486 21474 29538
rect 21870 29486 21922 29538
rect 23326 29486 23378 29538
rect 23438 29486 23490 29538
rect 1822 29374 1874 29426
rect 2382 29374 2434 29426
rect 3390 29374 3442 29426
rect 4398 29374 4450 29426
rect 6414 29374 6466 29426
rect 8654 29374 8706 29426
rect 9550 29374 9602 29426
rect 9998 29374 10050 29426
rect 11006 29374 11058 29426
rect 11902 29374 11954 29426
rect 12126 29374 12178 29426
rect 12350 29374 12402 29426
rect 13246 29374 13298 29426
rect 14030 29374 14082 29426
rect 14254 29374 14306 29426
rect 14478 29374 14530 29426
rect 14590 29374 14642 29426
rect 15150 29374 15202 29426
rect 15598 29374 15650 29426
rect 18062 29374 18114 29426
rect 19406 29374 19458 29426
rect 21198 29374 21250 29426
rect 23662 29374 23714 29426
rect 3838 29262 3890 29314
rect 7758 29262 7810 29314
rect 10334 29262 10386 29314
rect 10782 29262 10834 29314
rect 11230 29262 11282 29314
rect 11678 29262 11730 29314
rect 12014 29262 12066 29314
rect 13582 29262 13634 29314
rect 15598 29262 15650 29314
rect 16046 29262 16098 29314
rect 16382 29262 16434 29314
rect 18510 29262 18562 29314
rect 20974 29262 21026 29314
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 9886 28814 9938 28866
rect 23214 28814 23266 28866
rect 23662 28814 23714 28866
rect 24782 28814 24834 28866
rect 3614 28702 3666 28754
rect 5070 28702 5122 28754
rect 7646 28702 7698 28754
rect 8094 28702 8146 28754
rect 8990 28702 9042 28754
rect 11902 28702 11954 28754
rect 21310 28702 21362 28754
rect 21758 28702 21810 28754
rect 22990 28702 23042 28754
rect 1710 28590 1762 28642
rect 2830 28590 2882 28642
rect 4174 28590 4226 28642
rect 5630 28590 5682 28642
rect 7198 28590 7250 28642
rect 8878 28590 8930 28642
rect 10446 28590 10498 28642
rect 11454 28590 11506 28642
rect 13694 28590 13746 28642
rect 14590 28590 14642 28642
rect 15262 28590 15314 28642
rect 16606 28590 16658 28642
rect 17502 28590 17554 28642
rect 18622 28590 18674 28642
rect 19070 28590 19122 28642
rect 19406 28590 19458 28642
rect 21534 28590 21586 28642
rect 21982 28590 22034 28642
rect 22430 28590 22482 28642
rect 23886 28590 23938 28642
rect 24110 28590 24162 28642
rect 24894 28590 24946 28642
rect 25342 28590 25394 28642
rect 25678 28590 25730 28642
rect 26238 28590 26290 28642
rect 5742 28478 5794 28530
rect 6190 28478 6242 28530
rect 15710 28478 15762 28530
rect 16046 28478 16098 28530
rect 17166 28478 17218 28530
rect 19294 28478 19346 28530
rect 20190 28478 20242 28530
rect 20302 28478 20354 28530
rect 24334 28478 24386 28530
rect 24670 28478 24722 28530
rect 2046 28366 2098 28418
rect 6638 28366 6690 28418
rect 13358 28366 13410 28418
rect 13582 28366 13634 28418
rect 14030 28366 14082 28418
rect 14926 28366 14978 28418
rect 17278 28366 17330 28418
rect 17838 28366 17890 28418
rect 18286 28366 18338 28418
rect 19854 28366 19906 28418
rect 20526 28366 20578 28418
rect 25118 28366 25170 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 8878 28030 8930 28082
rect 11230 28030 11282 28082
rect 15486 28030 15538 28082
rect 16270 28030 16322 28082
rect 18062 28030 18114 28082
rect 18622 28030 18674 28082
rect 20750 28030 20802 28082
rect 3614 27918 3666 27970
rect 5070 27918 5122 27970
rect 6526 27918 6578 27970
rect 8318 27918 8370 27970
rect 12238 27918 12290 27970
rect 13694 27918 13746 27970
rect 14926 27918 14978 27970
rect 15822 27918 15874 27970
rect 23774 27918 23826 27970
rect 23998 27918 24050 27970
rect 25566 27918 25618 27970
rect 26014 27918 26066 27970
rect 2942 27806 2994 27858
rect 3390 27806 3442 27858
rect 3950 27806 4002 27858
rect 7646 27806 7698 27858
rect 8542 27806 8594 27858
rect 9774 27806 9826 27858
rect 11118 27806 11170 27858
rect 11342 27806 11394 27858
rect 12462 27806 12514 27858
rect 13470 27806 13522 27858
rect 14814 27806 14866 27858
rect 16046 27806 16098 27858
rect 16382 27806 16434 27858
rect 18398 27806 18450 27858
rect 18846 27806 18898 27858
rect 19070 27806 19122 27858
rect 19854 27806 19906 27858
rect 23326 27806 23378 27858
rect 24110 27806 24162 27858
rect 25230 27806 25282 27858
rect 25790 27806 25842 27858
rect 26126 27806 26178 27858
rect 2270 27694 2322 27746
rect 7198 27694 7250 27746
rect 10670 27694 10722 27746
rect 14590 27694 14642 27746
rect 16270 27694 16322 27746
rect 17614 27694 17666 27746
rect 20302 27694 20354 27746
rect 22542 27694 22594 27746
rect 22990 27694 23042 27746
rect 26574 27694 26626 27746
rect 12798 27582 12850 27634
rect 18958 27582 19010 27634
rect 23102 27582 23154 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 11678 27246 11730 27298
rect 19742 27246 19794 27298
rect 21422 27246 21474 27298
rect 22318 27246 22370 27298
rect 26014 27246 26066 27298
rect 4958 27134 5010 27186
rect 9214 27134 9266 27186
rect 12350 27134 12402 27186
rect 13806 27134 13858 27186
rect 20302 27134 20354 27186
rect 23102 27134 23154 27186
rect 3166 27022 3218 27074
rect 5070 27022 5122 27074
rect 6526 27022 6578 27074
rect 7310 27022 7362 27074
rect 7870 27022 7922 27074
rect 9774 27022 9826 27074
rect 10446 27022 10498 27074
rect 11790 27022 11842 27074
rect 14254 27022 14306 27074
rect 14814 27022 14866 27074
rect 15150 27022 15202 27074
rect 16606 27022 16658 27074
rect 17166 27022 17218 27074
rect 18510 27022 18562 27074
rect 22206 27022 22258 27074
rect 23550 27022 23602 27074
rect 24782 27022 24834 27074
rect 26238 27022 26290 27074
rect 2606 26910 2658 26962
rect 3390 26910 3442 26962
rect 5518 26910 5570 26962
rect 7758 26910 7810 26962
rect 19630 26910 19682 26962
rect 22318 26910 22370 26962
rect 26350 26910 26402 26962
rect 7534 26798 7586 26850
rect 16494 26798 16546 26850
rect 18734 26798 18786 26850
rect 19294 26798 19346 26850
rect 19742 26798 19794 26850
rect 21534 26798 21586 26850
rect 21646 26798 21698 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 8430 26462 8482 26514
rect 16718 26462 16770 26514
rect 17390 26462 17442 26514
rect 21646 26462 21698 26514
rect 22318 26462 22370 26514
rect 22878 26462 22930 26514
rect 23774 26462 23826 26514
rect 23998 26462 24050 26514
rect 24334 26462 24386 26514
rect 26686 26462 26738 26514
rect 5294 26350 5346 26402
rect 6526 26350 6578 26402
rect 8766 26350 8818 26402
rect 8878 26350 8930 26402
rect 9998 26350 10050 26402
rect 15374 26350 15426 26402
rect 19294 26350 19346 26402
rect 21422 26350 21474 26402
rect 22654 26350 22706 26402
rect 24670 26350 24722 26402
rect 25230 26350 25282 26402
rect 26798 26350 26850 26402
rect 27582 26350 27634 26402
rect 28142 26350 28194 26402
rect 28478 26350 28530 26402
rect 2606 26238 2658 26290
rect 3166 26238 3218 26290
rect 5966 26238 6018 26290
rect 7870 26238 7922 26290
rect 9102 26238 9154 26290
rect 11566 26238 11618 26290
rect 13022 26238 13074 26290
rect 13246 26238 13298 26290
rect 13582 26238 13634 26290
rect 14254 26238 14306 26290
rect 16494 26238 16546 26290
rect 18398 26238 18450 26290
rect 19182 26238 19234 26290
rect 19518 26238 19570 26290
rect 20638 26238 20690 26290
rect 21086 26238 21138 26290
rect 21310 26238 21362 26290
rect 23214 26238 23266 26290
rect 23326 26238 23378 26290
rect 25790 26238 25842 26290
rect 26238 26238 26290 26290
rect 27246 26238 27298 26290
rect 2158 26126 2210 26178
rect 4062 26126 4114 26178
rect 8094 26126 8146 26178
rect 10894 26126 10946 26178
rect 17950 26126 18002 26178
rect 18734 26126 18786 26178
rect 19966 26126 20018 26178
rect 20190 26126 20242 26178
rect 23886 26126 23938 26178
rect 20414 26014 20466 26066
rect 22542 26014 22594 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 17390 25678 17442 25730
rect 4958 25566 5010 25618
rect 5854 25566 5906 25618
rect 9214 25566 9266 25618
rect 12910 25566 12962 25618
rect 13918 25566 13970 25618
rect 14478 25566 14530 25618
rect 19630 25566 19682 25618
rect 1822 25454 1874 25506
rect 3390 25454 3442 25506
rect 5070 25454 5122 25506
rect 5966 25454 6018 25506
rect 6190 25454 6242 25506
rect 7646 25454 7698 25506
rect 9550 25454 9602 25506
rect 11006 25454 11058 25506
rect 11790 25454 11842 25506
rect 12798 25454 12850 25506
rect 14814 25454 14866 25506
rect 15934 25454 15986 25506
rect 17278 25454 17330 25506
rect 17838 25454 17890 25506
rect 19406 25454 19458 25506
rect 20526 25454 20578 25506
rect 24894 25454 24946 25506
rect 25342 25454 25394 25506
rect 4510 25342 4562 25394
rect 7310 25342 7362 25394
rect 17726 25342 17778 25394
rect 18062 25342 18114 25394
rect 18622 25342 18674 25394
rect 19518 25342 19570 25394
rect 19742 25342 19794 25394
rect 19966 25342 20018 25394
rect 23774 25342 23826 25394
rect 25790 25342 25842 25394
rect 27246 25342 27298 25394
rect 2046 25230 2098 25282
rect 6526 25230 6578 25282
rect 7534 25230 7586 25282
rect 7758 25230 7810 25282
rect 13470 25230 13522 25282
rect 20750 25230 20802 25282
rect 26798 25230 26850 25282
rect 27358 25230 27410 25282
rect 27582 25230 27634 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 4062 24894 4114 24946
rect 8878 24894 8930 24946
rect 15262 24894 15314 24946
rect 15374 24894 15426 24946
rect 17502 24894 17554 24946
rect 20078 24894 20130 24946
rect 21646 24894 21698 24946
rect 22094 24894 22146 24946
rect 22766 24894 22818 24946
rect 2046 24782 2098 24834
rect 2382 24782 2434 24834
rect 2718 24782 2770 24834
rect 3614 24782 3666 24834
rect 5742 24782 5794 24834
rect 6414 24782 6466 24834
rect 9886 24782 9938 24834
rect 11790 24782 11842 24834
rect 14366 24782 14418 24834
rect 16046 24782 16098 24834
rect 18622 24782 18674 24834
rect 18958 24782 19010 24834
rect 19182 24782 19234 24834
rect 20862 24782 20914 24834
rect 23998 24782 24050 24834
rect 26126 24782 26178 24834
rect 27022 24782 27074 24834
rect 1710 24670 1762 24722
rect 3390 24670 3442 24722
rect 4174 24670 4226 24722
rect 4398 24670 4450 24722
rect 5966 24670 6018 24722
rect 6526 24670 6578 24722
rect 9550 24670 9602 24722
rect 10670 24670 10722 24722
rect 12686 24670 12738 24722
rect 15598 24670 15650 24722
rect 15934 24670 15986 24722
rect 17390 24670 17442 24722
rect 17614 24670 17666 24722
rect 18062 24670 18114 24722
rect 18286 24670 18338 24722
rect 19406 24670 19458 24722
rect 19630 24670 19682 24722
rect 19966 24670 20018 24722
rect 20190 24670 20242 24722
rect 20526 24670 20578 24722
rect 21086 24670 21138 24722
rect 23774 24670 23826 24722
rect 24110 24670 24162 24722
rect 24334 24670 24386 24722
rect 25230 24670 25282 24722
rect 28366 24670 28418 24722
rect 8094 24558 8146 24610
rect 8766 24558 8818 24610
rect 10222 24558 10274 24610
rect 14030 24558 14082 24610
rect 19518 24558 19570 24610
rect 23326 24558 23378 24610
rect 25342 24558 25394 24610
rect 4062 24446 4114 24498
rect 8654 24446 8706 24498
rect 24782 24446 24834 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 11790 24110 11842 24162
rect 19406 24110 19458 24162
rect 2494 23998 2546 24050
rect 2942 23998 2994 24050
rect 4734 23998 4786 24050
rect 21422 24110 21474 24162
rect 10782 23998 10834 24050
rect 19854 23998 19906 24050
rect 28142 23998 28194 24050
rect 1934 23886 1986 23938
rect 3950 23886 4002 23938
rect 4286 23886 4338 23938
rect 5630 23886 5682 23938
rect 6638 23886 6690 23938
rect 7646 23886 7698 23938
rect 8430 23886 8482 23938
rect 10110 23886 10162 23938
rect 11678 23886 11730 23938
rect 12126 23886 12178 23938
rect 12798 23886 12850 23938
rect 14142 23886 14194 23938
rect 14702 23886 14754 23938
rect 15374 23886 15426 23938
rect 17278 23886 17330 23938
rect 17726 23886 17778 23938
rect 18958 23886 19010 23938
rect 19742 23886 19794 23938
rect 19854 23886 19906 23938
rect 20302 23886 20354 23938
rect 20526 23886 20578 23938
rect 21310 23886 21362 23938
rect 23662 23886 23714 23938
rect 23998 23886 24050 23938
rect 26910 23886 26962 23938
rect 4174 23774 4226 23826
rect 4622 23774 4674 23826
rect 5070 23774 5122 23826
rect 5854 23774 5906 23826
rect 7310 23774 7362 23826
rect 7422 23774 7474 23826
rect 8206 23774 8258 23826
rect 10334 23774 10386 23826
rect 12910 23774 12962 23826
rect 15822 23774 15874 23826
rect 21870 23774 21922 23826
rect 24558 23774 24610 23826
rect 27246 23774 27298 23826
rect 27806 23774 27858 23826
rect 1710 23662 1762 23714
rect 4846 23662 4898 23714
rect 6638 23662 6690 23714
rect 14926 23662 14978 23714
rect 20414 23662 20466 23714
rect 21422 23662 21474 23714
rect 22654 23662 22706 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 2270 23326 2322 23378
rect 6862 23326 6914 23378
rect 16718 23326 16770 23378
rect 23662 23326 23714 23378
rect 25566 23326 25618 23378
rect 5518 23214 5570 23266
rect 8318 23214 8370 23266
rect 15038 23214 15090 23266
rect 16158 23214 16210 23266
rect 17390 23214 17442 23266
rect 18622 23214 18674 23266
rect 18734 23214 18786 23266
rect 22430 23214 22482 23266
rect 23774 23214 23826 23266
rect 24334 23214 24386 23266
rect 26910 23214 26962 23266
rect 1934 23102 1986 23154
rect 3838 23102 3890 23154
rect 5294 23102 5346 23154
rect 7758 23102 7810 23154
rect 8094 23102 8146 23154
rect 9102 23102 9154 23154
rect 10222 23102 10274 23154
rect 11342 23102 11394 23154
rect 12462 23102 12514 23154
rect 13246 23102 13298 23154
rect 13918 23102 13970 23154
rect 16494 23102 16546 23154
rect 17614 23102 17666 23154
rect 17838 23102 17890 23154
rect 18062 23102 18114 23154
rect 18958 23102 19010 23154
rect 19518 23102 19570 23154
rect 20974 23102 21026 23154
rect 22318 23102 22370 23154
rect 24558 23102 24610 23154
rect 26462 23102 26514 23154
rect 27358 23102 27410 23154
rect 27582 23102 27634 23154
rect 27806 23102 27858 23154
rect 28142 23102 28194 23154
rect 28366 23102 28418 23154
rect 28478 23102 28530 23154
rect 2718 22990 2770 23042
rect 7422 22990 7474 23042
rect 10110 22990 10162 23042
rect 11118 22990 11170 23042
rect 17726 22990 17778 23042
rect 22766 22990 22818 23042
rect 26686 22990 26738 23042
rect 1822 22878 1874 22930
rect 2718 22878 2770 22930
rect 6078 22878 6130 22930
rect 26014 22878 26066 22930
rect 26238 22878 26290 22930
rect 28926 22878 28978 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 5070 22542 5122 22594
rect 5966 22542 6018 22594
rect 6638 22542 6690 22594
rect 8766 22542 8818 22594
rect 24558 22542 24610 22594
rect 25118 22542 25170 22594
rect 4174 22430 4226 22482
rect 7982 22430 8034 22482
rect 10446 22430 10498 22482
rect 13582 22430 13634 22482
rect 18510 22430 18562 22482
rect 18734 22430 18786 22482
rect 20638 22430 20690 22482
rect 24222 22430 24274 22482
rect 1822 22318 1874 22370
rect 2718 22318 2770 22370
rect 2942 22318 2994 22370
rect 3166 22318 3218 22370
rect 3390 22318 3442 22370
rect 4286 22318 4338 22370
rect 8542 22318 8594 22370
rect 9774 22318 9826 22370
rect 10222 22318 10274 22370
rect 12238 22318 12290 22370
rect 12574 22318 12626 22370
rect 13806 22318 13858 22370
rect 14926 22318 14978 22370
rect 16158 22318 16210 22370
rect 16942 22318 16994 22370
rect 17166 22318 17218 22370
rect 17502 22318 17554 22370
rect 18846 22318 18898 22370
rect 19182 22318 19234 22370
rect 19294 22318 19346 22370
rect 19630 22318 19682 22370
rect 19854 22318 19906 22370
rect 22654 22318 22706 22370
rect 23550 22318 23602 22370
rect 23886 22318 23938 22370
rect 25342 22318 25394 22370
rect 25902 22318 25954 22370
rect 27694 22318 27746 22370
rect 3726 22206 3778 22258
rect 5742 22206 5794 22258
rect 6414 22206 6466 22258
rect 12462 22206 12514 22258
rect 13582 22206 13634 22258
rect 15822 22218 15874 22270
rect 17726 22206 17778 22258
rect 20750 22206 20802 22258
rect 21870 22206 21922 22258
rect 22430 22206 22482 22258
rect 26462 22206 26514 22258
rect 2046 22094 2098 22146
rect 3054 22094 3106 22146
rect 3950 22094 4002 22146
rect 4174 22094 4226 22146
rect 4846 22094 4898 22146
rect 4958 22094 5010 22146
rect 5854 22094 5906 22146
rect 6526 22094 6578 22146
rect 7422 22094 7474 22146
rect 14814 22094 14866 22146
rect 18174 22094 18226 22146
rect 20302 22094 20354 22146
rect 20526 22094 20578 22146
rect 22206 22094 22258 22146
rect 24110 22094 24162 22146
rect 24558 22094 24610 22146
rect 25006 22094 25058 22146
rect 25454 22094 25506 22146
rect 25678 22094 25730 22146
rect 28254 22094 28306 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 2382 21758 2434 21810
rect 2942 21758 2994 21810
rect 3166 21758 3218 21810
rect 3838 21758 3890 21810
rect 9998 21758 10050 21810
rect 10110 21758 10162 21810
rect 11678 21758 11730 21810
rect 12686 21758 12738 21810
rect 21310 21758 21362 21810
rect 21758 21758 21810 21810
rect 26686 21758 26738 21810
rect 2046 21646 2098 21698
rect 4398 21646 4450 21698
rect 5518 21646 5570 21698
rect 9662 21646 9714 21698
rect 11566 21646 11618 21698
rect 14030 21646 14082 21698
rect 17502 21646 17554 21698
rect 21422 21646 21474 21698
rect 22878 21646 22930 21698
rect 24222 21646 24274 21698
rect 25566 21646 25618 21698
rect 27470 21646 27522 21698
rect 28702 21646 28754 21698
rect 2718 21534 2770 21586
rect 3390 21534 3442 21586
rect 3726 21534 3778 21586
rect 6302 21534 6354 21586
rect 7310 21534 7362 21586
rect 8654 21534 8706 21586
rect 9886 21534 9938 21586
rect 10446 21534 10498 21586
rect 11006 21534 11058 21586
rect 13022 21534 13074 21586
rect 13246 21534 13298 21586
rect 15710 21534 15762 21586
rect 17390 21534 17442 21586
rect 19406 21534 19458 21586
rect 20862 21534 20914 21586
rect 22430 21534 22482 21586
rect 22654 21534 22706 21586
rect 23998 21534 24050 21586
rect 24334 21534 24386 21586
rect 26238 21534 26290 21586
rect 28142 21534 28194 21586
rect 28590 21534 28642 21586
rect 3278 21422 3330 21474
rect 12126 21422 12178 21474
rect 15374 21422 15426 21474
rect 16830 21422 16882 21474
rect 23774 21422 23826 21474
rect 28814 21422 28866 21474
rect 11678 21310 11730 21362
rect 13582 21310 13634 21362
rect 22206 21310 22258 21362
rect 24782 21310 24834 21362
rect 25790 21310 25842 21362
rect 26014 21310 26066 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 8318 20974 8370 21026
rect 18510 20974 18562 21026
rect 18846 20974 18898 21026
rect 19406 20974 19458 21026
rect 20302 20974 20354 21026
rect 20638 20974 20690 21026
rect 22318 20974 22370 21026
rect 4286 20862 4338 20914
rect 7198 20862 7250 20914
rect 12238 20862 12290 20914
rect 12686 20862 12738 20914
rect 18062 20862 18114 20914
rect 18510 20862 18562 20914
rect 21310 20862 21362 20914
rect 27470 20862 27522 20914
rect 2942 20750 2994 20802
rect 3054 20750 3106 20802
rect 3166 20750 3218 20802
rect 3390 20750 3442 20802
rect 3726 20750 3778 20802
rect 5854 20750 5906 20802
rect 6190 20750 6242 20802
rect 6638 20750 6690 20802
rect 6862 20750 6914 20802
rect 7646 20750 7698 20802
rect 8206 20750 8258 20802
rect 9102 20750 9154 20802
rect 9550 20750 9602 20802
rect 10446 20750 10498 20802
rect 11454 20750 11506 20802
rect 13806 20750 13858 20802
rect 15150 20750 15202 20802
rect 16158 20750 16210 20802
rect 16942 20750 16994 20802
rect 19294 20750 19346 20802
rect 20078 20750 20130 20802
rect 21646 20750 21698 20802
rect 22094 20750 22146 20802
rect 22542 20750 22594 20802
rect 24782 20750 24834 20802
rect 26798 20750 26850 20802
rect 1710 20638 1762 20690
rect 2718 20638 2770 20690
rect 5182 20638 5234 20690
rect 8990 20638 9042 20690
rect 10222 20638 10274 20690
rect 14366 20638 14418 20690
rect 15934 20638 15986 20690
rect 21422 20638 21474 20690
rect 22766 20638 22818 20690
rect 22878 20638 22930 20690
rect 24894 20638 24946 20690
rect 27358 20638 27410 20690
rect 2046 20526 2098 20578
rect 6078 20526 6130 20578
rect 7198 20526 7250 20578
rect 9774 20526 9826 20578
rect 10782 20526 10834 20578
rect 11566 20526 11618 20578
rect 11790 20526 11842 20578
rect 18958 20526 19010 20578
rect 19406 20526 19458 20578
rect 23326 20526 23378 20578
rect 24446 20526 24498 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 2718 20190 2770 20242
rect 3166 20190 3218 20242
rect 3502 20190 3554 20242
rect 8878 20190 8930 20242
rect 10558 20190 10610 20242
rect 12798 20190 12850 20242
rect 16606 20190 16658 20242
rect 17614 20190 17666 20242
rect 20302 20190 20354 20242
rect 1710 20078 1762 20130
rect 2046 20078 2098 20130
rect 5406 20078 5458 20130
rect 7758 20078 7810 20130
rect 8766 20078 8818 20130
rect 10782 20078 10834 20130
rect 11678 20078 11730 20130
rect 11902 20078 11954 20130
rect 12462 20078 12514 20130
rect 14366 20078 14418 20130
rect 16382 20078 16434 20130
rect 21534 20078 21586 20130
rect 21982 20078 22034 20130
rect 23886 20078 23938 20130
rect 24334 20078 24386 20130
rect 24782 20078 24834 20130
rect 26686 20078 26738 20130
rect 27918 20078 27970 20130
rect 2382 19966 2434 20018
rect 4958 19966 5010 20018
rect 5294 19966 5346 20018
rect 5630 19966 5682 20018
rect 7422 19966 7474 20018
rect 7982 19966 8034 20018
rect 8990 19966 9042 20018
rect 10334 19966 10386 20018
rect 10894 19966 10946 20018
rect 11454 19966 11506 20018
rect 12014 19966 12066 20018
rect 13358 19966 13410 20018
rect 13918 19966 13970 20018
rect 14590 19966 14642 20018
rect 14702 19966 14754 20018
rect 14926 19966 14978 20018
rect 15150 19966 15202 20018
rect 16270 19966 16322 20018
rect 16830 19966 16882 20018
rect 17726 19966 17778 20018
rect 18174 19966 18226 20018
rect 18398 19966 18450 20018
rect 21310 19966 21362 20018
rect 21758 19966 21810 20018
rect 23550 19966 23602 20018
rect 26126 19966 26178 20018
rect 27694 19966 27746 20018
rect 4062 19854 4114 19906
rect 4398 19854 4450 19906
rect 6078 19854 6130 19906
rect 6414 19854 6466 19906
rect 6974 19854 7026 19906
rect 8206 19854 8258 19906
rect 9886 19854 9938 19906
rect 15710 19854 15762 19906
rect 16718 19854 16770 19906
rect 18734 19854 18786 19906
rect 20190 19854 20242 19906
rect 21086 19854 21138 19906
rect 22094 19854 22146 19906
rect 22430 19854 22482 19906
rect 29486 19854 29538 19906
rect 6078 19742 6130 19794
rect 6526 19742 6578 19794
rect 7198 19742 7250 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 15486 19406 15538 19458
rect 15710 19406 15762 19458
rect 24110 19406 24162 19458
rect 25678 19406 25730 19458
rect 8878 19294 8930 19346
rect 12350 19294 12402 19346
rect 13582 19294 13634 19346
rect 15374 19294 15426 19346
rect 19406 19294 19458 19346
rect 20190 19294 20242 19346
rect 22430 19294 22482 19346
rect 23214 19294 23266 19346
rect 3054 19182 3106 19234
rect 3502 19182 3554 19234
rect 3950 19182 4002 19234
rect 9550 19182 9602 19234
rect 11006 19182 11058 19234
rect 11342 19182 11394 19234
rect 11902 19182 11954 19234
rect 12910 19182 12962 19234
rect 14030 19182 14082 19234
rect 14814 19182 14866 19234
rect 16382 19182 16434 19234
rect 17838 19182 17890 19234
rect 18510 19182 18562 19234
rect 20078 19182 20130 19234
rect 20638 19182 20690 19234
rect 21422 19182 21474 19234
rect 24670 19182 24722 19234
rect 24894 19182 24946 19234
rect 25230 19182 25282 19234
rect 1710 19070 1762 19122
rect 2494 19070 2546 19122
rect 4398 19070 4450 19122
rect 5742 19070 5794 19122
rect 10782 19070 10834 19122
rect 13918 19070 13970 19122
rect 14702 19070 14754 19122
rect 19182 19070 19234 19122
rect 21534 19070 21586 19122
rect 21982 19070 22034 19122
rect 23998 19070 24050 19122
rect 25006 19070 25058 19122
rect 2046 18958 2098 19010
rect 4174 18958 4226 19010
rect 4846 18958 4898 19010
rect 9326 18958 9378 19010
rect 9774 18958 9826 19010
rect 10446 18958 10498 19010
rect 20302 18958 20354 19010
rect 24110 18958 24162 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 2046 18622 2098 18674
rect 3278 18622 3330 18674
rect 10558 18622 10610 18674
rect 15598 18622 15650 18674
rect 16942 18622 16994 18674
rect 18286 18622 18338 18674
rect 19854 18622 19906 18674
rect 20414 18622 20466 18674
rect 20862 18622 20914 18674
rect 22318 18622 22370 18674
rect 23774 18622 23826 18674
rect 2942 18510 2994 18562
rect 3166 18510 3218 18562
rect 4510 18510 4562 18562
rect 5070 18510 5122 18562
rect 7534 18510 7586 18562
rect 11566 18510 11618 18562
rect 14702 18510 14754 18562
rect 18174 18510 18226 18562
rect 20638 18510 20690 18562
rect 22094 18510 22146 18562
rect 1710 18398 1762 18450
rect 2718 18398 2770 18450
rect 3838 18398 3890 18450
rect 5854 18398 5906 18450
rect 7422 18398 7474 18450
rect 8990 18398 9042 18450
rect 9550 18398 9602 18450
rect 10110 18398 10162 18450
rect 11006 18398 11058 18450
rect 12350 18398 12402 18450
rect 14142 18398 14194 18450
rect 17950 18398 18002 18450
rect 19182 18398 19234 18450
rect 19406 18398 19458 18450
rect 19966 18398 20018 18450
rect 20078 18398 20130 18450
rect 21646 18398 21698 18450
rect 21982 18398 22034 18450
rect 22766 18398 22818 18450
rect 23550 18398 23602 18450
rect 23774 18398 23826 18450
rect 24110 18398 24162 18450
rect 3054 18286 3106 18338
rect 5406 18286 5458 18338
rect 15822 18286 15874 18338
rect 20526 18286 20578 18338
rect 22542 18286 22594 18338
rect 7534 18174 7586 18226
rect 16046 18174 16098 18226
rect 16270 18174 16322 18226
rect 16494 18174 16546 18226
rect 18286 18174 18338 18226
rect 23102 18174 23154 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 10558 17838 10610 17890
rect 11230 17838 11282 17890
rect 18958 17838 19010 17890
rect 2270 17726 2322 17778
rect 4622 17726 4674 17778
rect 9886 17726 9938 17778
rect 13582 17726 13634 17778
rect 15710 17726 15762 17778
rect 16718 17726 16770 17778
rect 17390 17726 17442 17778
rect 18622 17726 18674 17778
rect 20638 17726 20690 17778
rect 23214 17726 23266 17778
rect 1822 17614 1874 17666
rect 1934 17614 1986 17666
rect 2382 17614 2434 17666
rect 3278 17614 3330 17666
rect 3726 17614 3778 17666
rect 6862 17614 6914 17666
rect 8766 17614 8818 17666
rect 11230 17614 11282 17666
rect 12014 17614 12066 17666
rect 12350 17614 12402 17666
rect 13470 17614 13522 17666
rect 14030 17614 14082 17666
rect 14926 17614 14978 17666
rect 15374 17614 15426 17666
rect 15598 17614 15650 17666
rect 16158 17614 16210 17666
rect 16382 17614 16434 17666
rect 16606 17614 16658 17666
rect 18846 17614 18898 17666
rect 19406 17614 19458 17666
rect 21646 17614 21698 17666
rect 22206 17614 22258 17666
rect 22766 17614 22818 17666
rect 24446 17614 24498 17666
rect 25678 17614 25730 17666
rect 2830 17502 2882 17554
rect 8318 17502 8370 17554
rect 9438 17502 9490 17554
rect 12798 17502 12850 17554
rect 15150 17502 15202 17554
rect 16718 17502 16770 17554
rect 19630 17502 19682 17554
rect 20078 17502 20130 17554
rect 22878 17502 22930 17554
rect 2158 17390 2210 17442
rect 3838 17390 3890 17442
rect 4062 17390 4114 17442
rect 10670 17390 10722 17442
rect 11566 17390 11618 17442
rect 12574 17390 12626 17442
rect 13694 17390 13746 17442
rect 14590 17390 14642 17442
rect 18062 17390 18114 17442
rect 18958 17390 19010 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 1934 17054 1986 17106
rect 3838 17054 3890 17106
rect 4062 17054 4114 17106
rect 4734 17054 4786 17106
rect 7198 17054 7250 17106
rect 7310 17054 7362 17106
rect 8654 17054 8706 17106
rect 8990 17054 9042 17106
rect 10334 17054 10386 17106
rect 11566 17054 11618 17106
rect 11678 17054 11730 17106
rect 15374 17054 15426 17106
rect 15598 17054 15650 17106
rect 17502 17054 17554 17106
rect 17614 17054 17666 17106
rect 17726 17054 17778 17106
rect 18846 17054 18898 17106
rect 19406 17054 19458 17106
rect 19630 17054 19682 17106
rect 21198 17054 21250 17106
rect 2830 16942 2882 16994
rect 7870 16942 7922 16994
rect 8094 16942 8146 16994
rect 10558 16942 10610 16994
rect 10670 16942 10722 16994
rect 11230 16942 11282 16994
rect 15822 16942 15874 16994
rect 16382 16942 16434 16994
rect 16830 16942 16882 16994
rect 18510 16942 18562 16994
rect 20526 16942 20578 16994
rect 21982 16942 22034 16994
rect 22990 16942 23042 16994
rect 1822 16830 1874 16882
rect 2158 16830 2210 16882
rect 2270 16830 2322 16882
rect 3166 16830 3218 16882
rect 3614 16830 3666 16882
rect 4510 16830 4562 16882
rect 4958 16830 5010 16882
rect 5070 16830 5122 16882
rect 7758 16830 7810 16882
rect 8318 16830 8370 16882
rect 9662 16830 9714 16882
rect 11790 16830 11842 16882
rect 12238 16830 12290 16882
rect 12462 16830 12514 16882
rect 13022 16830 13074 16882
rect 13470 16830 13522 16882
rect 13918 16830 13970 16882
rect 14254 16830 14306 16882
rect 14590 16830 14642 16882
rect 14702 16830 14754 16882
rect 14926 16830 14978 16882
rect 15150 16830 15202 16882
rect 16158 16830 16210 16882
rect 16606 16830 16658 16882
rect 17838 16830 17890 16882
rect 17950 16830 18002 16882
rect 19182 16830 19234 16882
rect 19854 16830 19906 16882
rect 20414 16830 20466 16882
rect 20750 16830 20802 16882
rect 22430 16830 22482 16882
rect 24558 16830 24610 16882
rect 2046 16718 2098 16770
rect 4846 16718 4898 16770
rect 9998 16718 10050 16770
rect 15262 16718 15314 16770
rect 19518 16718 19570 16770
rect 20190 16718 20242 16770
rect 24782 16718 24834 16770
rect 16270 16606 16322 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 14030 16270 14082 16322
rect 22430 16270 22482 16322
rect 4622 16158 4674 16210
rect 11006 16158 11058 16210
rect 13470 16158 13522 16210
rect 13694 16158 13746 16210
rect 15262 16158 15314 16210
rect 18622 16158 18674 16210
rect 19406 16158 19458 16210
rect 20414 16158 20466 16210
rect 21646 16158 21698 16210
rect 24334 16158 24386 16210
rect 1710 16046 1762 16098
rect 3278 16046 3330 16098
rect 3614 16046 3666 16098
rect 5070 16046 5122 16098
rect 5854 16046 5906 16098
rect 7870 16046 7922 16098
rect 9550 16046 9602 16098
rect 10446 16046 10498 16098
rect 11342 16046 11394 16098
rect 11790 16046 11842 16098
rect 12238 16046 12290 16098
rect 12462 16046 12514 16098
rect 14926 16046 14978 16098
rect 15710 16046 15762 16098
rect 15934 16046 15986 16098
rect 16382 16046 16434 16098
rect 17054 16046 17106 16098
rect 17502 16046 17554 16098
rect 17614 16046 17666 16098
rect 18062 16046 18114 16098
rect 19070 16046 19122 16098
rect 19742 16046 19794 16098
rect 20526 16046 20578 16098
rect 20750 16046 20802 16098
rect 21310 16046 21362 16098
rect 21534 16046 21586 16098
rect 21758 16046 21810 16098
rect 21870 16046 21922 16098
rect 22542 16046 22594 16098
rect 23102 16046 23154 16098
rect 24670 16046 24722 16098
rect 26014 16046 26066 16098
rect 2046 15934 2098 15986
rect 2830 15934 2882 15986
rect 5630 15934 5682 15986
rect 8206 15934 8258 15986
rect 8990 15934 9042 15986
rect 9214 15934 9266 15986
rect 9886 15934 9938 15986
rect 9998 15934 10050 15986
rect 10222 15934 10274 15986
rect 14702 15934 14754 15986
rect 16158 15934 16210 15986
rect 18286 15934 18338 15986
rect 23214 15934 23266 15986
rect 3838 15822 3890 15874
rect 4062 15822 4114 15874
rect 7982 15822 8034 15874
rect 8542 15822 8594 15874
rect 11678 15822 11730 15874
rect 11902 15822 11954 15874
rect 12798 15822 12850 15874
rect 15150 15822 15202 15874
rect 15262 15822 15314 15874
rect 16046 15822 16098 15874
rect 17278 15822 17330 15874
rect 17390 15822 17442 15874
rect 19294 15822 19346 15874
rect 19518 15822 19570 15874
rect 20190 15822 20242 15874
rect 20302 15822 20354 15874
rect 22430 15822 22482 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 2046 15486 2098 15538
rect 2718 15486 2770 15538
rect 3278 15486 3330 15538
rect 8654 15486 8706 15538
rect 8990 15486 9042 15538
rect 10894 15486 10946 15538
rect 13246 15486 13298 15538
rect 13918 15486 13970 15538
rect 16046 15486 16098 15538
rect 16382 15486 16434 15538
rect 18734 15486 18786 15538
rect 19406 15486 19458 15538
rect 21422 15486 21474 15538
rect 22094 15486 22146 15538
rect 22766 15486 22818 15538
rect 1710 15374 1762 15426
rect 3502 15374 3554 15426
rect 4286 15374 4338 15426
rect 6190 15374 6242 15426
rect 6974 15374 7026 15426
rect 11230 15374 11282 15426
rect 12910 15374 12962 15426
rect 14814 15374 14866 15426
rect 17390 15374 17442 15426
rect 19742 15374 19794 15426
rect 21646 15374 21698 15426
rect 23214 15374 23266 15426
rect 2382 15262 2434 15314
rect 3166 15262 3218 15314
rect 3950 15262 4002 15314
rect 6078 15262 6130 15314
rect 7198 15262 7250 15314
rect 9550 15262 9602 15314
rect 9998 15262 10050 15314
rect 10670 15262 10722 15314
rect 12574 15262 12626 15314
rect 13470 15262 13522 15314
rect 14478 15262 14530 15314
rect 15374 15262 15426 15314
rect 15934 15262 15986 15314
rect 16158 15262 16210 15314
rect 16270 15262 16322 15314
rect 17502 15262 17554 15314
rect 18174 15262 18226 15314
rect 18622 15262 18674 15314
rect 20302 15262 20354 15314
rect 20526 15262 20578 15314
rect 21198 15262 21250 15314
rect 11678 15150 11730 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 2270 14702 2322 14754
rect 2718 14702 2770 14754
rect 3838 14702 3890 14754
rect 10782 14702 10834 14754
rect 11678 14702 11730 14754
rect 21982 14702 22034 14754
rect 2494 14590 2546 14642
rect 2942 14590 2994 14642
rect 9326 14590 9378 14642
rect 10222 14590 10274 14642
rect 10782 14590 10834 14642
rect 11230 14590 11282 14642
rect 11678 14590 11730 14642
rect 13022 14590 13074 14642
rect 14702 14590 14754 14642
rect 16158 14590 16210 14642
rect 16494 14590 16546 14642
rect 18174 14590 18226 14642
rect 18622 14590 18674 14642
rect 20862 14590 20914 14642
rect 21422 14590 21474 14642
rect 22542 14590 22594 14642
rect 3726 14478 3778 14530
rect 13582 14478 13634 14530
rect 14030 14478 14082 14530
rect 15374 14478 15426 14530
rect 16942 14478 16994 14530
rect 17614 14478 17666 14530
rect 18958 14478 19010 14530
rect 19518 14478 19570 14530
rect 22094 14478 22146 14530
rect 1710 14366 1762 14418
rect 2046 14366 2098 14418
rect 17502 14366 17554 14418
rect 21982 14366 22034 14418
rect 3390 14254 3442 14306
rect 3838 14254 3890 14306
rect 9886 14254 9938 14306
rect 12238 14254 12290 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 2046 13918 2098 13970
rect 2494 13918 2546 13970
rect 10334 13918 10386 13970
rect 11006 13918 11058 13970
rect 14030 13918 14082 13970
rect 14814 13918 14866 13970
rect 15150 13918 15202 13970
rect 15710 13918 15762 13970
rect 16270 13918 16322 13970
rect 18062 13918 18114 13970
rect 18510 13918 18562 13970
rect 18958 13918 19010 13970
rect 12798 13806 12850 13858
rect 13246 13806 13298 13858
rect 13694 13806 13746 13858
rect 1710 13694 1762 13746
rect 2942 13582 2994 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 2046 12798 2098 12850
rect 1710 12686 1762 12738
rect 2494 12686 2546 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 2046 12350 2098 12402
rect 1710 12126 1762 12178
rect 2494 12014 2546 12066
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 1710 11230 1762 11282
rect 2046 11230 2098 11282
rect 2494 11118 2546 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 1934 9774 1986 9826
rect 1710 9662 1762 9714
rect 2494 9662 2546 9714
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 2046 9214 2098 9266
rect 1710 8990 1762 9042
rect 2494 8878 2546 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 1710 8094 1762 8146
rect 2046 8094 2098 8146
rect 2494 7982 2546 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 2046 7646 2098 7698
rect 1710 7422 1762 7474
rect 2494 7310 2546 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 1710 6526 1762 6578
rect 2046 6526 2098 6578
rect 2494 6414 2546 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 2046 6078 2098 6130
rect 1710 5854 1762 5906
rect 2494 5742 2546 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 2494 5070 2546 5122
rect 1710 4958 1762 5010
rect 2046 4958 2098 5010
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 1710 3390 1762 3442
rect 2046 3390 2098 3442
rect 2494 3390 2546 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 2464 41200 2576 42000
rect 5824 41200 5936 42000
rect 9184 41200 9296 42000
rect 12544 41200 12656 42000
rect 15904 41200 16016 42000
rect 19264 41200 19376 42000
rect 22624 41200 22736 42000
rect 25984 41200 26096 42000
rect 29344 41200 29456 42000
rect 29708 41244 30100 41300
rect 5852 38668 5908 41200
rect 9212 38948 9268 41200
rect 8876 38892 9492 38948
rect 3612 38610 3668 38622
rect 5852 38612 6020 38668
rect 3612 38558 3614 38610
rect 3666 38558 3668 38610
rect 1820 38052 1876 38062
rect 1820 38050 1988 38052
rect 1820 37998 1822 38050
rect 1874 37998 1988 38050
rect 1820 37996 1988 37998
rect 1820 37986 1876 37996
rect 1820 37154 1876 37166
rect 1820 37102 1822 37154
rect 1874 37102 1876 37154
rect 1708 36258 1764 36270
rect 1708 36206 1710 36258
rect 1762 36206 1764 36258
rect 1708 36148 1764 36206
rect 1596 36092 1764 36148
rect 1148 36036 1204 36046
rect 1148 13860 1204 35980
rect 1596 35924 1652 36092
rect 1820 36036 1876 37102
rect 1932 36708 1988 37996
rect 3388 38050 3444 38062
rect 3388 37998 3390 38050
rect 3442 37998 3444 38050
rect 2380 37940 2436 37950
rect 2044 37826 2100 37838
rect 2044 37774 2046 37826
rect 2098 37774 2100 37826
rect 2044 36932 2100 37774
rect 2268 37828 2324 37838
rect 2268 37268 2324 37772
rect 2380 37492 2436 37884
rect 2380 37426 2436 37436
rect 2716 37826 2772 37838
rect 2716 37774 2718 37826
rect 2770 37774 2772 37826
rect 2716 37380 2772 37774
rect 2716 37314 2772 37324
rect 3388 37380 3444 37998
rect 3612 37938 3668 38558
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4284 38164 4340 38174
rect 4284 38050 4340 38108
rect 4284 37998 4286 38050
rect 4338 37998 4340 38050
rect 4284 37986 4340 37998
rect 5964 38052 6020 38612
rect 5964 37958 6020 37996
rect 6748 38610 6804 38622
rect 6748 38558 6750 38610
rect 6802 38558 6804 38610
rect 3612 37886 3614 37938
rect 3666 37886 3668 37938
rect 3612 37874 3668 37886
rect 4956 37938 5012 37950
rect 4956 37886 4958 37938
rect 5010 37886 5012 37938
rect 3948 37828 4004 37838
rect 4620 37828 4676 37838
rect 3948 37734 4004 37772
rect 4396 37826 4676 37828
rect 4396 37774 4622 37826
rect 4674 37774 4676 37826
rect 4396 37772 4676 37774
rect 4396 37604 4452 37772
rect 4620 37762 4676 37772
rect 3612 37548 4452 37604
rect 3612 37490 3668 37548
rect 3612 37438 3614 37490
rect 3666 37438 3668 37490
rect 3612 37426 3668 37438
rect 3388 37314 3444 37324
rect 3164 37268 3220 37278
rect 2268 37266 2548 37268
rect 2268 37214 2270 37266
rect 2322 37214 2548 37266
rect 2268 37212 2548 37214
rect 2268 37202 2324 37212
rect 2044 36866 2100 36876
rect 1932 36652 2212 36708
rect 2044 36260 2100 36270
rect 1596 33908 1652 35868
rect 1596 33842 1652 33852
rect 1708 35980 1876 36036
rect 1932 36258 2100 36260
rect 1932 36206 2046 36258
rect 2098 36206 2100 36258
rect 1932 36204 2100 36206
rect 1708 33348 1764 35980
rect 1820 35812 1876 35822
rect 1820 35698 1876 35756
rect 1820 35646 1822 35698
rect 1874 35646 1876 35698
rect 1820 35634 1876 35646
rect 1932 34916 1988 36204
rect 2044 36194 2100 36204
rect 2156 36148 2212 36652
rect 2492 36594 2548 37212
rect 2716 37156 2772 37166
rect 2716 37062 2772 37100
rect 3164 37154 3220 37212
rect 3164 37102 3166 37154
rect 3218 37102 3220 37154
rect 3164 37090 3220 37102
rect 2492 36542 2494 36594
rect 2546 36542 2548 36594
rect 2492 36530 2548 36542
rect 2940 36932 2996 36942
rect 2604 36484 2660 36494
rect 2604 36390 2660 36428
rect 2940 36482 2996 36876
rect 3836 36932 3892 36942
rect 3500 36708 3556 36718
rect 3500 36594 3556 36652
rect 3836 36706 3892 36876
rect 3836 36654 3838 36706
rect 3890 36654 3892 36706
rect 3836 36642 3892 36654
rect 3500 36542 3502 36594
rect 3554 36542 3556 36594
rect 3500 36530 3556 36542
rect 4060 36596 4116 36606
rect 4060 36502 4116 36540
rect 2940 36430 2942 36482
rect 2994 36430 2996 36482
rect 2940 36418 2996 36430
rect 4172 36482 4228 37548
rect 4172 36430 4174 36482
rect 4226 36430 4228 36482
rect 4172 36418 4228 36430
rect 4284 37266 4340 37278
rect 4284 37214 4286 37266
rect 4338 37214 4340 37266
rect 4284 36484 4340 37214
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 2156 36082 2212 36092
rect 4284 36036 4340 36428
rect 4844 36708 4900 36718
rect 4844 36482 4900 36652
rect 4844 36430 4846 36482
rect 4898 36430 4900 36482
rect 4844 36418 4900 36430
rect 4956 36372 5012 37886
rect 6524 37938 6580 37950
rect 6524 37886 6526 37938
rect 6578 37886 6580 37938
rect 6188 37826 6244 37838
rect 6188 37774 6190 37826
rect 6242 37774 6244 37826
rect 5404 37268 5460 37278
rect 5404 37174 5460 37212
rect 5852 37268 5908 37278
rect 5292 36484 5348 36494
rect 4284 35980 4900 36036
rect 1820 34860 1988 34916
rect 2044 35810 2100 35822
rect 2044 35758 2046 35810
rect 2098 35758 2100 35810
rect 1820 33460 1876 34860
rect 1932 34690 1988 34702
rect 1932 34638 1934 34690
rect 1986 34638 1988 34690
rect 1932 34468 1988 34638
rect 1932 34402 1988 34412
rect 2044 34132 2100 35758
rect 2380 35810 2436 35822
rect 2380 35758 2382 35810
rect 2434 35758 2436 35810
rect 2380 34916 2436 35758
rect 4396 35812 4452 35822
rect 4396 35718 4452 35756
rect 4844 35810 4900 35980
rect 4844 35758 4846 35810
rect 4898 35758 4900 35810
rect 4844 35746 4900 35758
rect 4956 35812 5012 36316
rect 4956 35746 5012 35756
rect 5068 36370 5124 36382
rect 5068 36318 5070 36370
rect 5122 36318 5124 36370
rect 2604 35698 2660 35710
rect 2604 35646 2606 35698
rect 2658 35646 2660 35698
rect 2604 35588 2660 35646
rect 3948 35700 4004 35710
rect 2604 35522 2660 35532
rect 3164 35586 3220 35598
rect 3164 35534 3166 35586
rect 3218 35534 3220 35586
rect 3164 35028 3220 35534
rect 3612 35588 3668 35598
rect 3612 35494 3668 35532
rect 2380 34850 2436 34860
rect 2492 34972 3220 35028
rect 2268 34692 2324 34702
rect 2492 34692 2548 34972
rect 3388 34914 3444 34926
rect 3388 34862 3390 34914
rect 3442 34862 3444 34914
rect 2828 34804 2884 34814
rect 2044 34038 2100 34076
rect 2156 34690 2548 34692
rect 2156 34638 2270 34690
rect 2322 34638 2548 34690
rect 2156 34636 2548 34638
rect 2604 34692 2660 34702
rect 1820 33404 2100 33460
rect 1708 33292 1988 33348
rect 1820 33124 1876 33134
rect 1708 33122 1876 33124
rect 1708 33070 1822 33122
rect 1874 33070 1876 33122
rect 1708 33068 1876 33070
rect 1708 31220 1764 33068
rect 1820 33058 1876 33068
rect 1596 31164 1764 31220
rect 1820 32450 1876 32462
rect 1820 32398 1822 32450
rect 1874 32398 1876 32450
rect 1596 30772 1652 31164
rect 1708 30996 1764 31006
rect 1708 30902 1764 30940
rect 1596 30716 1764 30772
rect 1708 30210 1764 30716
rect 1708 30158 1710 30210
rect 1762 30158 1764 30210
rect 1708 29876 1764 30158
rect 1708 29810 1764 29820
rect 1820 29652 1876 32398
rect 1932 30996 1988 33292
rect 2044 33124 2100 33404
rect 2156 33348 2212 34636
rect 2268 34626 2324 34636
rect 2268 34468 2324 34478
rect 2324 34412 2436 34468
rect 2268 34402 2324 34412
rect 2156 33282 2212 33292
rect 2268 34244 2324 34254
rect 2268 33346 2324 34188
rect 2268 33294 2270 33346
rect 2322 33294 2324 33346
rect 2268 33282 2324 33294
rect 2268 33124 2324 33134
rect 2044 33068 2268 33124
rect 2268 32564 2324 33068
rect 2044 32562 2324 32564
rect 2044 32510 2270 32562
rect 2322 32510 2324 32562
rect 2044 32508 2324 32510
rect 2044 31890 2100 32508
rect 2268 32498 2324 32508
rect 2380 32228 2436 34412
rect 2604 34132 2660 34636
rect 2604 34130 2772 34132
rect 2604 34078 2606 34130
rect 2658 34078 2772 34130
rect 2604 34076 2772 34078
rect 2604 34066 2660 34076
rect 2492 33236 2548 33246
rect 2492 33142 2548 33180
rect 2492 32676 2548 32686
rect 2716 32676 2772 34076
rect 2828 34020 2884 34748
rect 2940 34802 2996 34814
rect 2940 34750 2942 34802
rect 2994 34750 2996 34802
rect 2940 34468 2996 34750
rect 2940 34402 2996 34412
rect 3388 34692 3444 34862
rect 3836 34692 3892 34702
rect 3388 34636 3836 34692
rect 3388 34244 3444 34636
rect 3836 34598 3892 34636
rect 3388 34178 3444 34188
rect 2828 33346 2884 33964
rect 2828 33294 2830 33346
rect 2882 33294 2884 33346
rect 2828 33282 2884 33294
rect 3052 34132 3108 34142
rect 2940 33234 2996 33246
rect 2940 33182 2942 33234
rect 2994 33182 2996 33234
rect 2828 33124 2884 33134
rect 2940 33124 2996 33182
rect 2884 33068 2996 33124
rect 2828 33058 2884 33068
rect 2828 32676 2884 32686
rect 2716 32674 2884 32676
rect 2716 32622 2830 32674
rect 2882 32622 2884 32674
rect 2716 32620 2884 32622
rect 2492 32582 2548 32620
rect 2828 32610 2884 32620
rect 2940 32340 2996 33068
rect 3052 32562 3108 34076
rect 3164 34020 3220 34030
rect 3220 33964 3332 34020
rect 3164 33954 3220 33964
rect 3052 32510 3054 32562
rect 3106 32510 3108 32562
rect 3052 32498 3108 32510
rect 2940 32284 3220 32340
rect 2380 32172 2548 32228
rect 2268 32004 2324 32014
rect 2268 31910 2324 31948
rect 2044 31838 2046 31890
rect 2098 31838 2100 31890
rect 2044 31826 2100 31838
rect 2492 31220 2548 32172
rect 2604 31556 2660 31566
rect 2604 31462 2660 31500
rect 2940 31554 2996 31566
rect 2940 31502 2942 31554
rect 2994 31502 2996 31554
rect 2044 31108 2100 31118
rect 2044 31014 2100 31052
rect 1932 30324 1988 30940
rect 2492 30994 2548 31164
rect 2492 30942 2494 30994
rect 2546 30942 2548 30994
rect 2492 30930 2548 30942
rect 2716 31106 2772 31118
rect 2716 31054 2718 31106
rect 2770 31054 2772 31106
rect 1932 30258 1988 30268
rect 2044 30436 2100 30446
rect 2044 30098 2100 30380
rect 2044 30046 2046 30098
rect 2098 30046 2100 30098
rect 2044 30034 2100 30046
rect 1708 29596 1876 29652
rect 2604 29876 2660 29886
rect 1372 29540 1428 29550
rect 1148 13794 1204 13804
rect 1260 20804 1316 20814
rect 1260 4788 1316 20748
rect 1372 16100 1428 29484
rect 1708 28642 1764 29596
rect 2044 29540 2100 29550
rect 2044 29446 2100 29484
rect 1708 28590 1710 28642
rect 1762 28590 1764 28642
rect 1708 26852 1764 28590
rect 1820 29426 1876 29438
rect 1820 29374 1822 29426
rect 1874 29374 1876 29426
rect 1820 28532 1876 29374
rect 2380 29428 2436 29438
rect 2380 29334 2436 29372
rect 1820 28466 1876 28476
rect 2044 28420 2100 28430
rect 2044 28418 2548 28420
rect 2044 28366 2046 28418
rect 2098 28366 2548 28418
rect 2044 28364 2548 28366
rect 2044 28354 2100 28364
rect 1708 26786 1764 26796
rect 2268 27746 2324 27758
rect 2268 27694 2270 27746
rect 2322 27694 2324 27746
rect 2268 26516 2324 27694
rect 2268 26450 2324 26460
rect 2156 26178 2212 26190
rect 2156 26126 2158 26178
rect 2210 26126 2212 26178
rect 2156 25620 2212 26126
rect 2156 25554 2212 25564
rect 2380 25844 2436 25854
rect 1820 25506 1876 25518
rect 1820 25454 1822 25506
rect 1874 25454 1876 25506
rect 1820 25060 1876 25454
rect 2044 25284 2100 25294
rect 2044 25190 2100 25228
rect 1820 25004 2324 25060
rect 1820 24948 1876 25004
rect 1820 24882 1876 24892
rect 2044 24836 2100 24846
rect 2044 24834 2212 24836
rect 2044 24782 2046 24834
rect 2098 24782 2212 24834
rect 2044 24780 2212 24782
rect 2044 24770 2100 24780
rect 1708 24722 1764 24734
rect 1708 24670 1710 24722
rect 1762 24670 1764 24722
rect 1708 24052 1764 24670
rect 1708 23986 1764 23996
rect 1932 23938 1988 23950
rect 1932 23886 1934 23938
rect 1986 23886 1988 23938
rect 1708 23714 1764 23726
rect 1708 23662 1710 23714
rect 1762 23662 1764 23714
rect 1596 21364 1652 21374
rect 1596 20804 1652 21308
rect 1708 20916 1764 23662
rect 1932 23156 1988 23886
rect 1932 23062 1988 23100
rect 1820 22930 1876 22942
rect 1820 22878 1822 22930
rect 1874 22878 1876 22930
rect 1820 22372 1876 22878
rect 2156 22708 2212 24780
rect 2268 23378 2324 25004
rect 2380 24834 2436 25788
rect 2380 24782 2382 24834
rect 2434 24782 2436 24834
rect 2380 24052 2436 24782
rect 2492 24276 2548 28364
rect 2604 27972 2660 29820
rect 2604 27906 2660 27916
rect 2604 26962 2660 26974
rect 2604 26910 2606 26962
rect 2658 26910 2660 26962
rect 2604 26516 2660 26910
rect 2716 26908 2772 31054
rect 2940 30772 2996 31502
rect 3164 31106 3220 32284
rect 3164 31054 3166 31106
rect 3218 31054 3220 31106
rect 3164 31042 3220 31054
rect 3276 32004 3332 33964
rect 3724 34018 3780 34030
rect 3724 33966 3726 34018
rect 3778 33966 3780 34018
rect 3500 33460 3556 33470
rect 3500 33366 3556 33404
rect 3612 32676 3668 32686
rect 3052 30772 3108 30782
rect 2940 30770 3108 30772
rect 2940 30718 3054 30770
rect 3106 30718 3108 30770
rect 2940 30716 3108 30718
rect 2940 30100 2996 30716
rect 3052 30706 3108 30716
rect 3276 30436 3332 31948
rect 3388 32338 3444 32350
rect 3388 32286 3390 32338
rect 3442 32286 3444 32338
rect 3388 31780 3444 32286
rect 3500 31892 3556 31902
rect 3500 31798 3556 31836
rect 3388 31714 3444 31724
rect 3612 31332 3668 32620
rect 3724 32004 3780 33966
rect 3724 31938 3780 31948
rect 3836 32450 3892 32462
rect 3836 32398 3838 32450
rect 3890 32398 3892 32450
rect 3836 31668 3892 32398
rect 3948 32116 4004 35644
rect 5068 35476 5124 36318
rect 5292 35698 5348 36428
rect 5740 36484 5796 36494
rect 5740 36390 5796 36428
rect 5852 36482 5908 37212
rect 5852 36430 5854 36482
rect 5906 36430 5908 36482
rect 5852 36418 5908 36430
rect 5964 37266 6020 37278
rect 5964 37214 5966 37266
rect 6018 37214 6020 37266
rect 5964 36596 6020 37214
rect 5964 36482 6020 36540
rect 5964 36430 5966 36482
rect 6018 36430 6020 36482
rect 5964 36418 6020 36430
rect 5292 35646 5294 35698
rect 5346 35646 5348 35698
rect 5292 35634 5348 35646
rect 6076 35588 6132 35598
rect 6076 35494 6132 35532
rect 5068 35410 5124 35420
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4284 35028 4340 35038
rect 4172 35026 4340 35028
rect 4172 34974 4286 35026
rect 4338 34974 4340 35026
rect 4172 34972 4340 34974
rect 6188 35028 6244 37774
rect 6412 37604 6468 37614
rect 6412 37266 6468 37548
rect 6412 37214 6414 37266
rect 6466 37214 6468 37266
rect 6412 37202 6468 37214
rect 6524 37492 6580 37886
rect 6748 37940 6804 38558
rect 6860 38276 6916 38286
rect 7084 38276 7140 38286
rect 6860 38274 7140 38276
rect 6860 38222 6862 38274
rect 6914 38222 7086 38274
rect 7138 38222 7140 38274
rect 6860 38220 7140 38222
rect 6860 38210 6916 38220
rect 7084 38210 7140 38220
rect 8092 38274 8148 38286
rect 8092 38222 8094 38274
rect 8146 38222 8148 38274
rect 7756 38164 7812 38174
rect 7756 38070 7812 38108
rect 7308 38052 7364 38062
rect 7308 37958 7364 37996
rect 6748 37938 7028 37940
rect 6748 37886 6750 37938
rect 6802 37886 7028 37938
rect 6748 37884 7028 37886
rect 6748 37874 6804 37884
rect 6300 37156 6356 37166
rect 6300 36596 6356 37100
rect 6524 37044 6580 37436
rect 6748 37380 6804 37390
rect 6748 37286 6804 37324
rect 6860 37156 6916 37166
rect 6860 37062 6916 37100
rect 6524 36978 6580 36988
rect 6412 36596 6468 36606
rect 6300 36540 6412 36596
rect 6300 35810 6356 36540
rect 6412 36530 6468 36540
rect 6972 36484 7028 37884
rect 7308 37266 7364 37278
rect 7308 37214 7310 37266
rect 7362 37214 7364 37266
rect 7308 36596 7364 37214
rect 8092 37268 8148 38222
rect 8876 38162 8932 38892
rect 8876 38110 8878 38162
rect 8930 38110 8932 38162
rect 8876 38098 8932 38110
rect 9436 38050 9492 38892
rect 9884 38164 9940 38174
rect 9436 37998 9438 38050
rect 9490 37998 9492 38050
rect 9436 37986 9492 37998
rect 9660 38162 9940 38164
rect 9660 38110 9886 38162
rect 9938 38110 9940 38162
rect 9660 38108 9940 38110
rect 8204 37940 8260 37950
rect 8204 37846 8260 37884
rect 9548 37940 9604 37950
rect 9548 37604 9604 37884
rect 8652 37492 8708 37502
rect 8204 37268 8260 37278
rect 8092 37266 8260 37268
rect 8092 37214 8206 37266
rect 8258 37214 8260 37266
rect 8092 37212 8260 37214
rect 7308 36530 7364 36540
rect 7756 37154 7812 37166
rect 7756 37102 7758 37154
rect 7810 37102 7812 37154
rect 7756 37044 7812 37102
rect 6972 36390 7028 36428
rect 6412 36260 6468 36270
rect 6412 36166 6468 36204
rect 7644 36258 7700 36270
rect 7644 36206 7646 36258
rect 7698 36206 7700 36258
rect 6860 35924 6916 35934
rect 6860 35830 6916 35868
rect 6300 35758 6302 35810
rect 6354 35758 6356 35810
rect 6300 35746 6356 35758
rect 7308 35812 7364 35822
rect 7308 35718 7364 35756
rect 6412 35698 6468 35710
rect 6412 35646 6414 35698
rect 6466 35646 6468 35698
rect 6412 35476 6468 35646
rect 6412 35410 6468 35420
rect 7644 35364 7700 36206
rect 7644 35298 7700 35308
rect 6188 34972 6468 35028
rect 4172 33012 4228 34972
rect 4284 34962 4340 34972
rect 4732 34802 4788 34814
rect 4732 34750 4734 34802
rect 4786 34750 4788 34802
rect 4732 34692 4788 34750
rect 4844 34804 4900 34814
rect 4844 34710 4900 34748
rect 6188 34804 6244 34814
rect 6188 34802 6356 34804
rect 6188 34750 6190 34802
rect 6242 34750 6356 34802
rect 6188 34748 6356 34750
rect 6188 34738 6244 34748
rect 5068 34692 5124 34702
rect 4732 34626 4788 34636
rect 4956 34690 5124 34692
rect 4956 34638 5070 34690
rect 5122 34638 5124 34690
rect 4956 34636 5124 34638
rect 4284 34242 4340 34254
rect 4284 34190 4286 34242
rect 4338 34190 4340 34242
rect 4284 33908 4340 34190
rect 4284 33572 4340 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4284 33516 4564 33572
rect 4396 33346 4452 33358
rect 4396 33294 4398 33346
rect 4450 33294 4452 33346
rect 4284 33012 4340 33022
rect 4172 32956 4284 33012
rect 4284 32946 4340 32956
rect 4396 32788 4452 33294
rect 4396 32722 4452 32732
rect 4284 32564 4340 32574
rect 4508 32564 4564 33516
rect 4844 33460 4900 33470
rect 4956 33460 5012 34636
rect 5068 34626 5124 34636
rect 5628 34690 5684 34702
rect 5628 34638 5630 34690
rect 5682 34638 5684 34690
rect 5628 34020 5684 34638
rect 6188 34468 6244 34478
rect 5628 33954 5684 33964
rect 5852 34130 5908 34142
rect 5852 34078 5854 34130
rect 5906 34078 5908 34130
rect 5852 33572 5908 34078
rect 6188 34130 6244 34412
rect 6188 34078 6190 34130
rect 6242 34078 6244 34130
rect 6188 34066 6244 34078
rect 6300 34132 6356 34748
rect 6300 34066 6356 34076
rect 5852 33506 5908 33516
rect 4844 33458 5012 33460
rect 4844 33406 4846 33458
rect 4898 33406 5012 33458
rect 4844 33404 5012 33406
rect 4844 33394 4900 33404
rect 4284 32562 4564 32564
rect 4284 32510 4286 32562
rect 4338 32510 4564 32562
rect 4284 32508 4564 32510
rect 4732 33346 4788 33358
rect 4732 33294 4734 33346
rect 4786 33294 4788 33346
rect 4284 32498 4340 32508
rect 4732 32340 4788 33294
rect 4956 33348 5012 33404
rect 4956 33282 5012 33292
rect 5628 33348 5684 33358
rect 5628 33254 5684 33292
rect 6300 33236 6356 33246
rect 5180 33124 5236 33134
rect 5180 33030 5236 33068
rect 5964 33122 6020 33134
rect 5964 33070 5966 33122
rect 6018 33070 6020 33122
rect 5292 32674 5348 32686
rect 5292 32622 5294 32674
rect 5346 32622 5348 32674
rect 3948 32050 4004 32060
rect 4284 32284 5012 32340
rect 4284 31778 4340 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4732 32004 4788 32014
rect 4284 31726 4286 31778
rect 4338 31726 4340 31778
rect 4284 31714 4340 31726
rect 4396 31778 4452 31790
rect 4396 31726 4398 31778
rect 4450 31726 4452 31778
rect 3836 31602 3892 31612
rect 4396 31332 4452 31726
rect 3164 30380 3332 30436
rect 3500 31276 4452 31332
rect 3052 30324 3108 30362
rect 3052 30258 3108 30268
rect 3164 30322 3220 30380
rect 3164 30270 3166 30322
rect 3218 30270 3220 30322
rect 3164 30258 3220 30270
rect 2940 30044 3220 30100
rect 2828 29988 2884 29998
rect 2828 29894 2884 29932
rect 3052 29876 3108 29886
rect 2940 29820 3052 29876
rect 2940 29650 2996 29820
rect 3052 29810 3108 29820
rect 2940 29598 2942 29650
rect 2994 29598 2996 29650
rect 2828 28642 2884 28654
rect 2828 28590 2830 28642
rect 2882 28590 2884 28642
rect 2828 28532 2884 28590
rect 2828 28466 2884 28476
rect 2940 27858 2996 29598
rect 2940 27806 2942 27858
rect 2994 27806 2996 27858
rect 2940 27794 2996 27806
rect 3164 27748 3220 30044
rect 3388 29426 3444 29438
rect 3388 29374 3390 29426
rect 3442 29374 3444 29426
rect 3388 29316 3444 29374
rect 3500 29316 3556 31276
rect 4732 31220 4788 31948
rect 4844 31890 4900 31902
rect 4844 31838 4846 31890
rect 4898 31838 4900 31890
rect 4844 31780 4900 31838
rect 4844 31714 4900 31724
rect 4732 31164 4900 31220
rect 3612 31108 3668 31118
rect 3612 30660 3668 31052
rect 4284 30994 4340 31006
rect 4284 30942 4286 30994
rect 4338 30942 4340 30994
rect 3836 30882 3892 30894
rect 3836 30830 3838 30882
rect 3890 30830 3892 30882
rect 3612 30604 3780 30660
rect 3612 30210 3668 30222
rect 3612 30158 3614 30210
rect 3666 30158 3668 30210
rect 3612 29988 3668 30158
rect 3612 29922 3668 29932
rect 3388 29260 3500 29316
rect 3500 29250 3556 29260
rect 3612 29428 3668 29438
rect 3500 29092 3556 29102
rect 3276 27972 3332 27982
rect 3276 27860 3332 27916
rect 3388 27860 3444 27870
rect 3276 27858 3444 27860
rect 3276 27806 3390 27858
rect 3442 27806 3444 27858
rect 3276 27804 3444 27806
rect 3388 27794 3444 27804
rect 3164 27692 3332 27748
rect 3164 27076 3220 27114
rect 3164 27010 3220 27020
rect 3276 26908 3332 27692
rect 3500 27636 3556 29036
rect 3612 28754 3668 29372
rect 3612 28702 3614 28754
rect 3666 28702 3668 28754
rect 3612 28690 3668 28702
rect 2716 26852 3108 26908
rect 2604 26450 2660 26460
rect 2604 26292 2660 26302
rect 2604 26198 2660 26236
rect 2716 24834 2772 24846
rect 2716 24782 2718 24834
rect 2770 24782 2772 24834
rect 2492 24220 2660 24276
rect 2492 24052 2548 24062
rect 2380 24050 2548 24052
rect 2380 23998 2494 24050
rect 2546 23998 2548 24050
rect 2380 23996 2548 23998
rect 2492 23986 2548 23996
rect 2268 23326 2270 23378
rect 2322 23326 2324 23378
rect 2268 23314 2324 23326
rect 2156 22652 2548 22708
rect 2492 22484 2548 22652
rect 2604 22596 2660 24220
rect 2716 23380 2772 24782
rect 2940 24052 2996 24062
rect 2940 23958 2996 23996
rect 2716 23314 2772 23324
rect 2716 23042 2772 23054
rect 2716 22990 2718 23042
rect 2770 22990 2772 23042
rect 2716 22930 2772 22990
rect 2716 22878 2718 22930
rect 2770 22878 2772 22930
rect 2716 22866 2772 22878
rect 2604 22540 2884 22596
rect 2492 22428 2772 22484
rect 1820 22278 1876 22316
rect 2380 22372 2436 22382
rect 2044 22148 2100 22158
rect 2044 22054 2100 22092
rect 2380 21810 2436 22316
rect 2716 22370 2772 22428
rect 2716 22318 2718 22370
rect 2770 22318 2772 22370
rect 2716 22306 2772 22318
rect 2380 21758 2382 21810
rect 2434 21758 2436 21810
rect 2044 21700 2100 21710
rect 2044 21606 2100 21644
rect 2268 21476 2324 21486
rect 1932 21420 2268 21476
rect 1708 20860 1876 20916
rect 1596 20748 1764 20804
rect 1708 20692 1764 20748
rect 1708 20626 1764 20636
rect 1708 20468 1764 20478
rect 1708 20130 1764 20412
rect 1708 20078 1710 20130
rect 1762 20078 1764 20130
rect 1708 19796 1764 20078
rect 1708 19730 1764 19740
rect 1708 19124 1764 19134
rect 1708 18676 1764 19068
rect 1708 18610 1764 18620
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 17780 1764 18398
rect 1708 17714 1764 17724
rect 1820 17666 1876 20860
rect 1932 18676 1988 21420
rect 2268 21410 2324 21420
rect 2380 20916 2436 21758
rect 2716 21586 2772 21598
rect 2716 21534 2718 21586
rect 2770 21534 2772 21586
rect 2716 21476 2772 21534
rect 2828 21588 2884 22540
rect 2940 22372 2996 22382
rect 3052 22372 3108 26852
rect 3164 26852 3332 26908
rect 3388 27580 3556 27636
rect 3612 27970 3668 27982
rect 3612 27918 3614 27970
rect 3666 27918 3668 27970
rect 3388 26962 3444 27580
rect 3388 26910 3390 26962
rect 3442 26910 3444 26962
rect 3388 26898 3444 26910
rect 3612 26908 3668 27918
rect 3500 26852 3668 26908
rect 3164 26290 3220 26852
rect 3164 26238 3166 26290
rect 3218 26238 3220 26290
rect 3164 26226 3220 26238
rect 3276 26516 3332 26526
rect 3276 25284 3332 26460
rect 3388 26180 3444 26190
rect 3388 25506 3444 26124
rect 3388 25454 3390 25506
rect 3442 25454 3444 25506
rect 3388 25442 3444 25454
rect 3388 25284 3444 25294
rect 3276 25228 3388 25284
rect 3164 25060 3220 25070
rect 3220 25004 3332 25060
rect 3164 24994 3220 25004
rect 3164 22372 3220 22382
rect 3052 22370 3220 22372
rect 3052 22318 3166 22370
rect 3218 22318 3220 22370
rect 3052 22316 3220 22318
rect 2940 21810 2996 22316
rect 3164 22306 3220 22316
rect 2940 21758 2942 21810
rect 2994 21758 2996 21810
rect 2940 21746 2996 21758
rect 3052 22146 3108 22158
rect 3052 22094 3054 22146
rect 3106 22094 3108 22146
rect 2828 21522 2884 21532
rect 2716 21410 2772 21420
rect 3052 21252 3108 22094
rect 3164 21812 3220 21822
rect 3276 21812 3332 25004
rect 3388 24722 3444 25228
rect 3388 24670 3390 24722
rect 3442 24670 3444 24722
rect 3388 24658 3444 24670
rect 3500 24388 3556 26852
rect 3612 24834 3668 24846
rect 3612 24782 3614 24834
rect 3666 24782 3668 24834
rect 3612 24500 3668 24782
rect 3612 24434 3668 24444
rect 3388 24332 3556 24388
rect 3388 22596 3444 24332
rect 3724 24276 3780 30604
rect 3836 29652 3892 30830
rect 3948 30436 4004 30446
rect 3948 29876 4004 30380
rect 4284 30436 4340 30942
rect 4732 30994 4788 31006
rect 4732 30942 4734 30994
rect 4786 30942 4788 30994
rect 4732 30884 4788 30942
rect 4732 30818 4788 30828
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4284 30370 4340 30380
rect 4508 30324 4564 30334
rect 4060 30100 4116 30110
rect 4060 30098 4452 30100
rect 4060 30046 4062 30098
rect 4114 30046 4452 30098
rect 4060 30044 4452 30046
rect 4060 30034 4116 30044
rect 3948 29820 4116 29876
rect 3836 29586 3892 29596
rect 3948 29428 4004 29438
rect 3836 29314 3892 29326
rect 3836 29262 3838 29314
rect 3890 29262 3892 29314
rect 3836 28644 3892 29262
rect 3836 28578 3892 28588
rect 3948 27860 4004 29372
rect 3612 24220 3780 24276
rect 3836 27858 4004 27860
rect 3836 27806 3950 27858
rect 4002 27806 4004 27858
rect 3836 27804 4004 27806
rect 3836 27076 3892 27804
rect 3948 27794 4004 27804
rect 3388 22530 3444 22540
rect 3500 24164 3556 24174
rect 3164 21810 3332 21812
rect 3164 21758 3166 21810
rect 3218 21758 3332 21810
rect 3164 21756 3332 21758
rect 3388 22370 3444 22382
rect 3388 22318 3390 22370
rect 3442 22318 3444 22370
rect 3164 21746 3220 21756
rect 2380 20850 2436 20860
rect 2828 21196 3108 21252
rect 3164 21588 3220 21598
rect 2716 20690 2772 20702
rect 2716 20638 2718 20690
rect 2770 20638 2772 20690
rect 2044 20578 2100 20590
rect 2044 20526 2046 20578
rect 2098 20526 2100 20578
rect 2044 20356 2100 20526
rect 2044 20300 2548 20356
rect 2044 20132 2100 20142
rect 2044 20130 2212 20132
rect 2044 20078 2046 20130
rect 2098 20078 2212 20130
rect 2044 20076 2212 20078
rect 2044 20066 2100 20076
rect 2156 19124 2212 20076
rect 2380 20020 2436 20030
rect 2380 19572 2436 19964
rect 2492 19796 2548 20300
rect 2716 20242 2772 20638
rect 2716 20190 2718 20242
rect 2770 20190 2772 20242
rect 2716 20178 2772 20190
rect 2828 20132 2884 21196
rect 2940 20916 2996 20926
rect 2940 20802 2996 20860
rect 2940 20750 2942 20802
rect 2994 20750 2996 20802
rect 2940 20738 2996 20750
rect 3052 20804 3108 20814
rect 3052 20710 3108 20748
rect 3164 20802 3220 21532
rect 3388 21588 3444 22318
rect 3276 21474 3332 21486
rect 3276 21422 3278 21474
rect 3330 21422 3332 21474
rect 3276 20916 3332 21422
rect 3276 20850 3332 20860
rect 3164 20750 3166 20802
rect 3218 20750 3220 20802
rect 3164 20738 3220 20750
rect 3388 20802 3444 21532
rect 3388 20750 3390 20802
rect 3442 20750 3444 20802
rect 3388 20738 3444 20750
rect 3164 20580 3220 20590
rect 3500 20580 3556 24108
rect 3612 21588 3668 24220
rect 3836 23154 3892 27020
rect 4060 26908 4116 29820
rect 4396 29764 4452 30044
rect 4508 30098 4564 30268
rect 4508 30046 4510 30098
rect 4562 30046 4564 30098
rect 4508 29764 4564 30046
rect 4284 29708 4564 29764
rect 4844 29988 4900 31164
rect 4172 29316 4228 29326
rect 4172 28642 4228 29260
rect 4284 29092 4340 29708
rect 4396 29428 4452 29438
rect 4396 29334 4452 29372
rect 4284 29026 4340 29036
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4172 28590 4174 28642
rect 4226 28590 4228 28642
rect 4172 28578 4228 28590
rect 4284 28644 4340 28654
rect 4284 26908 4340 28588
rect 4844 27972 4900 29932
rect 4956 29540 5012 32284
rect 5292 32116 5348 32622
rect 5292 32050 5348 32060
rect 5180 32004 5236 32014
rect 5180 31778 5236 31948
rect 5180 31726 5182 31778
rect 5234 31726 5236 31778
rect 5180 31714 5236 31726
rect 5628 31556 5684 31566
rect 5628 30994 5684 31500
rect 5964 31444 6020 33070
rect 6300 32562 6356 33180
rect 6300 32510 6302 32562
rect 6354 32510 6356 32562
rect 5964 31378 6020 31388
rect 6188 31778 6244 31790
rect 6188 31726 6190 31778
rect 6242 31726 6244 31778
rect 6188 31668 6244 31726
rect 5628 30942 5630 30994
rect 5682 30942 5684 30994
rect 5628 30930 5684 30942
rect 6076 30994 6132 31006
rect 6076 30942 6078 30994
rect 6130 30942 6132 30994
rect 5180 30882 5236 30894
rect 5180 30830 5182 30882
rect 5234 30830 5236 30882
rect 4956 27972 5012 29484
rect 5068 30210 5124 30222
rect 5068 30158 5070 30210
rect 5122 30158 5124 30210
rect 5068 28756 5124 30158
rect 5180 30212 5236 30830
rect 6076 30324 6132 30942
rect 6076 30258 6132 30268
rect 5180 30146 5236 30156
rect 6188 30100 6244 31612
rect 6300 30996 6356 32510
rect 6412 32228 6468 34972
rect 7756 34916 7812 36988
rect 8204 36484 8260 37212
rect 8540 37156 8596 37166
rect 8204 36418 8260 36428
rect 8428 37154 8596 37156
rect 8428 37102 8542 37154
rect 8594 37102 8596 37154
rect 8428 37100 8596 37102
rect 8092 36260 8148 36270
rect 8092 36166 8148 36204
rect 8204 35476 8260 35486
rect 7980 34916 8036 34926
rect 7756 34914 8036 34916
rect 7756 34862 7982 34914
rect 8034 34862 8036 34914
rect 7756 34860 8036 34862
rect 7980 34850 8036 34860
rect 8204 34914 8260 35420
rect 8204 34862 8206 34914
rect 8258 34862 8260 34914
rect 8204 34850 8260 34862
rect 8316 34916 8372 34926
rect 8428 34916 8484 37100
rect 8540 37090 8596 37100
rect 8540 36372 8596 36382
rect 8652 36372 8708 37436
rect 8540 36370 8708 36372
rect 8540 36318 8542 36370
rect 8594 36318 8708 36370
rect 8540 36316 8708 36318
rect 8540 36306 8596 36316
rect 8316 34914 8484 34916
rect 8316 34862 8318 34914
rect 8370 34862 8484 34914
rect 8316 34860 8484 34862
rect 8316 34850 8372 34860
rect 6524 34804 6580 34814
rect 6524 34710 6580 34748
rect 6860 34802 6916 34814
rect 6860 34750 6862 34802
rect 6914 34750 6916 34802
rect 6748 34244 6804 34254
rect 6860 34244 6916 34750
rect 8204 34468 8260 34478
rect 7868 34356 7924 34366
rect 7868 34262 7924 34300
rect 6748 34242 6916 34244
rect 6748 34190 6750 34242
rect 6802 34190 6916 34242
rect 6748 34188 6916 34190
rect 6748 34178 6804 34188
rect 6412 32162 6468 32172
rect 6748 33572 6804 33582
rect 6860 33572 6916 34188
rect 7868 33908 7924 33918
rect 6860 33516 7028 33572
rect 6748 32562 6804 33516
rect 6748 32510 6750 32562
rect 6802 32510 6804 32562
rect 6748 32116 6804 32510
rect 6524 32060 6804 32116
rect 6860 33346 6916 33358
rect 6860 33294 6862 33346
rect 6914 33294 6916 33346
rect 6860 33012 6916 33294
rect 6524 31892 6580 32060
rect 6412 31780 6468 31790
rect 6524 31780 6580 31836
rect 6412 31778 6580 31780
rect 6412 31726 6414 31778
rect 6466 31726 6580 31778
rect 6412 31724 6580 31726
rect 6636 31890 6692 31902
rect 6636 31838 6638 31890
rect 6690 31838 6692 31890
rect 6636 31780 6692 31838
rect 6412 31714 6468 31724
rect 6636 31714 6692 31724
rect 6860 31220 6916 32956
rect 6748 31164 6916 31220
rect 6972 33346 7028 33516
rect 7084 33460 7140 33470
rect 7140 33404 7252 33460
rect 7084 33366 7140 33404
rect 6972 33294 6974 33346
rect 7026 33294 7028 33346
rect 6524 30996 6580 31006
rect 6300 30994 6580 30996
rect 6300 30942 6526 30994
rect 6578 30942 6580 30994
rect 6300 30940 6580 30942
rect 6524 30884 6580 30940
rect 6524 30818 6580 30828
rect 6412 30324 6468 30334
rect 6412 30230 6468 30268
rect 6636 30212 6692 30222
rect 6636 30118 6692 30156
rect 6076 30044 6244 30100
rect 5068 28662 5124 28700
rect 5180 29540 5236 29550
rect 5068 27972 5124 27982
rect 4956 27970 5124 27972
rect 4956 27918 5070 27970
rect 5122 27918 5124 27970
rect 4956 27916 5124 27918
rect 4844 27906 4900 27916
rect 5068 27906 5124 27916
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4956 27188 5012 27198
rect 4956 27094 5012 27132
rect 5068 27076 5124 27086
rect 5068 26982 5124 27020
rect 3948 26852 4116 26908
rect 4172 26852 4340 26908
rect 3948 24164 4004 26852
rect 4060 26180 4116 26190
rect 4060 26086 4116 26124
rect 4060 24948 4116 24958
rect 4060 24854 4116 24892
rect 4172 24724 4228 26852
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4508 25620 4564 25630
rect 4564 25564 4676 25620
rect 4508 25554 4564 25564
rect 4620 25508 4676 25564
rect 4508 25396 4564 25406
rect 4172 24630 4228 24668
rect 4284 25340 4508 25396
rect 3948 24098 4004 24108
rect 4060 24500 4116 24510
rect 3948 23940 4004 23950
rect 3948 23846 4004 23884
rect 4060 23828 4116 24444
rect 4284 23938 4340 25340
rect 4508 25302 4564 25340
rect 4396 24724 4452 24734
rect 4620 24724 4676 25452
rect 4956 25618 5012 25630
rect 4956 25566 4958 25618
rect 5010 25566 5012 25618
rect 4956 24948 5012 25566
rect 5068 25620 5124 25630
rect 5068 25506 5124 25564
rect 5068 25454 5070 25506
rect 5122 25454 5124 25506
rect 5068 25442 5124 25454
rect 4956 24882 5012 24892
rect 4396 24722 4676 24724
rect 4396 24670 4398 24722
rect 4450 24670 4676 24722
rect 4396 24668 4676 24670
rect 4396 24658 4452 24668
rect 4620 24500 4676 24668
rect 4620 24434 4676 24444
rect 5068 24836 5124 24846
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4732 24052 4788 24062
rect 4732 24050 5012 24052
rect 4732 23998 4734 24050
rect 4786 23998 5012 24050
rect 4732 23996 5012 23998
rect 4732 23986 4788 23996
rect 4284 23886 4286 23938
rect 4338 23886 4340 23938
rect 4284 23874 4340 23886
rect 4172 23828 4228 23838
rect 4060 23772 4172 23828
rect 4172 23734 4228 23772
rect 4620 23828 4676 23838
rect 4620 23734 4676 23772
rect 3836 23102 3838 23154
rect 3890 23102 3892 23154
rect 3836 23090 3892 23102
rect 4732 23716 4788 23726
rect 4732 22932 4788 23660
rect 4844 23714 4900 23726
rect 4844 23662 4846 23714
rect 4898 23662 4900 23714
rect 4844 23604 4900 23662
rect 4844 23538 4900 23548
rect 4956 23156 5012 23996
rect 5068 23826 5124 24780
rect 5068 23774 5070 23826
rect 5122 23774 5124 23826
rect 5068 23762 5124 23774
rect 4956 23090 5012 23100
rect 4732 22876 4900 22932
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4172 22484 4228 22494
rect 4172 22390 4228 22428
rect 4284 22372 4340 22382
rect 4844 22372 4900 22876
rect 5068 22820 5124 22830
rect 5068 22594 5124 22764
rect 5068 22542 5070 22594
rect 5122 22542 5124 22594
rect 5068 22530 5124 22542
rect 4284 22278 4340 22316
rect 4732 22316 4900 22372
rect 3724 22260 3780 22270
rect 3724 22166 3780 22204
rect 3948 22146 4004 22158
rect 3948 22094 3950 22146
rect 4002 22094 4004 22146
rect 3948 22036 4004 22094
rect 4172 22148 4228 22158
rect 4172 22054 4228 22092
rect 3948 21970 4004 21980
rect 3836 21812 3892 21822
rect 3836 21718 3892 21756
rect 4732 21812 4788 22316
rect 4844 22148 4900 22158
rect 4844 22054 4900 22092
rect 4956 22146 5012 22158
rect 4956 22094 4958 22146
rect 5010 22094 5012 22146
rect 4732 21746 4788 21756
rect 4396 21700 4452 21710
rect 4284 21698 4452 21700
rect 4284 21646 4398 21698
rect 4450 21646 4452 21698
rect 4284 21644 4452 21646
rect 3724 21588 3780 21598
rect 3612 21586 3780 21588
rect 3612 21534 3726 21586
rect 3778 21534 3780 21586
rect 3612 21532 3780 21534
rect 3724 21522 3780 21532
rect 4284 21588 4340 21644
rect 4396 21634 4452 21644
rect 3836 21028 3892 21038
rect 3724 20972 3836 21028
rect 3724 20804 3780 20972
rect 3836 20962 3892 20972
rect 4284 20914 4340 21532
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4284 20862 4286 20914
rect 4338 20862 4340 20914
rect 4284 20850 4340 20862
rect 3164 20242 3220 20524
rect 3164 20190 3166 20242
rect 3218 20190 3220 20242
rect 3164 20178 3220 20190
rect 3388 20524 3556 20580
rect 3612 20802 3780 20804
rect 3612 20750 3726 20802
rect 3778 20750 3780 20802
rect 3612 20748 3780 20750
rect 2828 20066 2884 20076
rect 3052 19908 3108 19918
rect 2492 19740 2884 19796
rect 2380 19506 2436 19516
rect 2716 19236 2772 19246
rect 2492 19124 2548 19134
rect 2156 19122 2548 19124
rect 2156 19070 2494 19122
rect 2546 19070 2548 19122
rect 2156 19068 2548 19070
rect 2492 19058 2548 19068
rect 2044 19012 2100 19022
rect 2044 19010 2436 19012
rect 2044 18958 2046 19010
rect 2098 18958 2436 19010
rect 2044 18956 2436 18958
rect 2044 18946 2100 18956
rect 2268 18788 2324 18798
rect 2044 18676 2100 18686
rect 1932 18674 2100 18676
rect 1932 18622 2046 18674
rect 2098 18622 2100 18674
rect 1932 18620 2100 18622
rect 2044 18610 2100 18620
rect 2268 18004 2324 18732
rect 2380 18676 2436 18956
rect 2716 18900 2772 19180
rect 2716 18834 2772 18844
rect 2380 18610 2436 18620
rect 2716 18452 2772 18462
rect 2604 18450 2772 18452
rect 2604 18398 2718 18450
rect 2770 18398 2772 18450
rect 2604 18396 2772 18398
rect 2044 17948 2324 18004
rect 2380 18004 2436 18014
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1820 17602 1876 17614
rect 1932 17668 1988 17678
rect 1932 17574 1988 17612
rect 1932 17220 1988 17230
rect 1932 17106 1988 17164
rect 1932 17054 1934 17106
rect 1986 17054 1988 17106
rect 1932 17042 1988 17054
rect 1372 16034 1428 16044
rect 1708 16884 1764 16894
rect 1708 16098 1764 16828
rect 1820 16884 1876 16894
rect 1820 16882 1988 16884
rect 1820 16830 1822 16882
rect 1874 16830 1988 16882
rect 1820 16828 1988 16830
rect 1820 16818 1876 16828
rect 1708 16046 1710 16098
rect 1762 16046 1764 16098
rect 1484 15988 1540 15998
rect 1540 15932 1652 15988
rect 1484 15922 1540 15932
rect 1596 15428 1652 15932
rect 1708 15764 1764 16046
rect 1708 15698 1764 15708
rect 1708 15428 1764 15438
rect 1484 15426 1764 15428
rect 1484 15374 1710 15426
rect 1762 15374 1764 15426
rect 1484 15372 1764 15374
rect 1484 14420 1540 15372
rect 1708 15362 1764 15372
rect 1484 14354 1540 14364
rect 1708 14418 1764 14430
rect 1708 14366 1710 14418
rect 1762 14366 1764 14418
rect 1708 14196 1764 14366
rect 1932 14308 1988 16828
rect 2044 16770 2100 17948
rect 2380 17892 2436 17948
rect 2268 17836 2436 17892
rect 2268 17778 2324 17836
rect 2268 17726 2270 17778
rect 2322 17726 2324 17778
rect 2268 17714 2324 17726
rect 2380 17668 2436 17678
rect 2380 17666 2548 17668
rect 2380 17614 2382 17666
rect 2434 17614 2548 17666
rect 2380 17612 2548 17614
rect 2380 17602 2436 17612
rect 2156 17442 2212 17454
rect 2156 17390 2158 17442
rect 2210 17390 2212 17442
rect 2156 17108 2212 17390
rect 2156 17052 2436 17108
rect 2044 16718 2046 16770
rect 2098 16718 2100 16770
rect 2044 16706 2100 16718
rect 2156 16882 2212 16894
rect 2156 16830 2158 16882
rect 2210 16830 2212 16882
rect 2044 15988 2100 15998
rect 2156 15988 2212 16830
rect 2268 16882 2324 16894
rect 2268 16830 2270 16882
rect 2322 16830 2324 16882
rect 2268 16772 2324 16830
rect 2268 16706 2324 16716
rect 2044 15986 2212 15988
rect 2044 15934 2046 15986
rect 2098 15934 2212 15986
rect 2044 15932 2212 15934
rect 2044 15922 2100 15932
rect 2380 15876 2436 17052
rect 2492 16772 2548 17612
rect 2492 16706 2548 16716
rect 2156 15820 2436 15876
rect 2044 15540 2100 15550
rect 2156 15540 2212 15820
rect 2044 15538 2212 15540
rect 2044 15486 2046 15538
rect 2098 15486 2212 15538
rect 2044 15484 2212 15486
rect 2492 15764 2548 15774
rect 2044 15474 2100 15484
rect 2380 15316 2436 15326
rect 2380 15222 2436 15260
rect 2268 14756 2324 14766
rect 2044 14754 2324 14756
rect 2044 14702 2270 14754
rect 2322 14702 2324 14754
rect 2044 14700 2324 14702
rect 2044 14418 2100 14700
rect 2268 14690 2324 14700
rect 2492 14642 2548 15708
rect 2492 14590 2494 14642
rect 2546 14590 2548 14642
rect 2492 14578 2548 14590
rect 2044 14366 2046 14418
rect 2098 14366 2100 14418
rect 2044 14354 2100 14366
rect 2492 14420 2548 14430
rect 1708 14130 1764 14140
rect 1820 14252 1988 14308
rect 1708 13746 1764 13758
rect 1708 13694 1710 13746
rect 1762 13694 1764 13746
rect 1708 13636 1764 13694
rect 1708 13300 1764 13580
rect 1708 13234 1764 13244
rect 1708 12738 1764 12750
rect 1708 12686 1710 12738
rect 1762 12686 1764 12738
rect 1708 12404 1764 12686
rect 1708 12338 1764 12348
rect 1708 12178 1764 12190
rect 1708 12126 1710 12178
rect 1762 12126 1764 12178
rect 1708 12068 1764 12126
rect 1708 11508 1764 12012
rect 1708 11442 1764 11452
rect 1708 11282 1764 11294
rect 1708 11230 1710 11282
rect 1762 11230 1764 11282
rect 1708 11172 1764 11230
rect 1708 10612 1764 11116
rect 1708 10546 1764 10556
rect 1708 9716 1764 9726
rect 1820 9716 1876 14252
rect 2044 13972 2100 13982
rect 2044 13878 2100 13916
rect 2492 13970 2548 14364
rect 2492 13918 2494 13970
rect 2546 13918 2548 13970
rect 2492 13906 2548 13918
rect 2604 13636 2660 18396
rect 2716 18386 2772 18396
rect 2828 17554 2884 19740
rect 3052 19236 3108 19852
rect 3388 19796 3444 20524
rect 3500 20244 3556 20254
rect 3612 20244 3668 20748
rect 3724 20738 3780 20748
rect 3724 20580 3780 20590
rect 3780 20524 3892 20580
rect 3724 20514 3780 20524
rect 3500 20242 3668 20244
rect 3500 20190 3502 20242
rect 3554 20190 3668 20242
rect 3500 20188 3668 20190
rect 3500 20178 3556 20188
rect 3612 20020 3668 20030
rect 3668 19964 3780 20020
rect 3612 19954 3668 19964
rect 3388 19740 3668 19796
rect 3052 19234 3332 19236
rect 3052 19182 3054 19234
rect 3106 19182 3332 19234
rect 3052 19180 3332 19182
rect 3052 19170 3108 19180
rect 3052 18676 3108 18686
rect 3108 18620 3220 18676
rect 3052 18610 3108 18620
rect 2940 18564 2996 18574
rect 2940 18470 2996 18508
rect 3164 18562 3220 18620
rect 3164 18510 3166 18562
rect 3218 18510 3220 18562
rect 3164 18498 3220 18510
rect 3276 18674 3332 19180
rect 3276 18622 3278 18674
rect 3330 18622 3332 18674
rect 3052 18340 3108 18350
rect 2828 17502 2830 17554
rect 2882 17502 2884 17554
rect 2828 17490 2884 17502
rect 2940 18338 3108 18340
rect 2940 18286 3054 18338
rect 3106 18286 3108 18338
rect 2940 18284 3108 18286
rect 2828 16994 2884 17006
rect 2828 16942 2830 16994
rect 2882 16942 2884 16994
rect 2828 16212 2884 16942
rect 2716 16156 2884 16212
rect 2716 15538 2772 16156
rect 2716 15486 2718 15538
rect 2770 15486 2772 15538
rect 2716 15474 2772 15486
rect 2828 15986 2884 15998
rect 2828 15934 2830 15986
rect 2882 15934 2884 15986
rect 2828 15316 2884 15934
rect 2716 15260 2884 15316
rect 2716 14754 2772 15260
rect 2940 15204 2996 18284
rect 3052 18274 3108 18284
rect 3276 17668 3332 18622
rect 3276 17574 3332 17612
rect 3500 19234 3556 19246
rect 3500 19182 3502 19234
rect 3554 19182 3556 19234
rect 3164 16882 3220 16894
rect 3164 16830 3166 16882
rect 3218 16830 3220 16882
rect 3164 16772 3220 16830
rect 3164 15988 3220 16716
rect 3276 16324 3332 16334
rect 3276 16100 3332 16268
rect 3276 16098 3444 16100
rect 3276 16046 3278 16098
rect 3330 16046 3444 16098
rect 3276 16044 3444 16046
rect 3276 16034 3332 16044
rect 3164 15922 3220 15932
rect 3276 15540 3332 15550
rect 2716 14702 2718 14754
rect 2770 14702 2772 14754
rect 2716 14690 2772 14702
rect 2828 15148 2996 15204
rect 3052 15538 3332 15540
rect 3052 15486 3278 15538
rect 3330 15486 3332 15538
rect 3052 15484 3332 15486
rect 2828 14644 2884 15148
rect 3052 15092 3108 15484
rect 3276 15474 3332 15484
rect 3164 15314 3220 15326
rect 3388 15316 3444 16044
rect 3500 15764 3556 19182
rect 3612 16882 3668 19740
rect 3724 18452 3780 19964
rect 3836 19012 3892 20524
rect 4956 20244 5012 22094
rect 5180 21140 5236 29484
rect 5628 28644 5684 28654
rect 5628 28550 5684 28588
rect 5740 28532 5796 28542
rect 5740 27076 5796 28476
rect 6076 27636 6132 30044
rect 5740 27010 5796 27020
rect 5964 27580 6132 27636
rect 6188 29652 6244 29662
rect 6188 28530 6244 29596
rect 6188 28478 6190 28530
rect 6242 28478 6244 28530
rect 5516 26962 5572 26974
rect 5516 26910 5518 26962
rect 5570 26910 5572 26962
rect 5292 26402 5348 26414
rect 5292 26350 5294 26402
rect 5346 26350 5348 26402
rect 5292 25284 5348 26350
rect 5292 23154 5348 25228
rect 5516 25396 5572 26910
rect 5964 26908 6020 27580
rect 6188 26908 6244 28478
rect 6412 29428 6468 29438
rect 6748 29428 6804 31164
rect 6860 30996 6916 31006
rect 6860 30902 6916 30940
rect 6972 30436 7028 33294
rect 6972 30370 7028 30380
rect 7084 31668 7140 31678
rect 6972 29652 7028 29662
rect 6972 29538 7028 29596
rect 6972 29486 6974 29538
rect 7026 29486 7028 29538
rect 6972 29474 7028 29486
rect 6412 29426 6804 29428
rect 6412 29374 6414 29426
rect 6466 29374 6804 29426
rect 6412 29372 6804 29374
rect 6412 28532 6468 29372
rect 6412 28466 6468 28476
rect 6748 28756 6804 28766
rect 6636 28418 6692 28430
rect 6636 28366 6638 28418
rect 6690 28366 6692 28418
rect 6524 27972 6580 27982
rect 6524 27074 6580 27916
rect 6524 27022 6526 27074
rect 6578 27022 6580 27074
rect 6524 27010 6580 27022
rect 5852 26852 6020 26908
rect 6076 26852 6244 26908
rect 5852 25620 5908 26852
rect 5516 23266 5572 25340
rect 5740 25564 5852 25620
rect 5628 24948 5684 24958
rect 5628 24276 5684 24892
rect 5740 24834 5796 25564
rect 5852 25526 5908 25564
rect 5964 26290 6020 26302
rect 5964 26238 5966 26290
rect 6018 26238 6020 26290
rect 5964 26180 6020 26238
rect 5740 24782 5742 24834
rect 5794 24782 5796 24834
rect 5740 24770 5796 24782
rect 5964 25506 6020 26124
rect 5964 25454 5966 25506
rect 6018 25454 6020 25506
rect 5852 24724 5908 24734
rect 5628 24220 5796 24276
rect 5628 23938 5684 23950
rect 5628 23886 5630 23938
rect 5682 23886 5684 23938
rect 5628 23828 5684 23886
rect 5628 23762 5684 23772
rect 5740 23492 5796 24220
rect 5852 23826 5908 24668
rect 5964 24722 6020 25454
rect 6076 24836 6132 26852
rect 6636 26628 6692 28366
rect 6636 26562 6692 26572
rect 6524 26404 6580 26414
rect 6748 26404 6804 28700
rect 6524 26402 6804 26404
rect 6524 26350 6526 26402
rect 6578 26350 6804 26402
rect 6524 26348 6804 26350
rect 6524 26338 6580 26348
rect 6188 25508 6244 25518
rect 6244 25452 6468 25508
rect 6188 25414 6244 25452
rect 6412 25060 6468 25452
rect 6524 25396 6580 25406
rect 6524 25282 6580 25340
rect 6524 25230 6526 25282
rect 6578 25230 6580 25282
rect 6524 25218 6580 25230
rect 6636 25284 6692 25294
rect 6412 25004 6580 25060
rect 6076 24770 6132 24780
rect 6412 24836 6468 24846
rect 6412 24742 6468 24780
rect 5964 24670 5966 24722
rect 6018 24670 6020 24722
rect 5964 24658 6020 24670
rect 6524 24722 6580 25004
rect 6524 24670 6526 24722
rect 6578 24670 6580 24722
rect 6524 24658 6580 24670
rect 6636 23938 6692 25228
rect 6636 23886 6638 23938
rect 6690 23886 6692 23938
rect 6636 23874 6692 23886
rect 5852 23774 5854 23826
rect 5906 23774 5908 23826
rect 5852 23762 5908 23774
rect 6636 23716 6692 23726
rect 6636 23622 6692 23660
rect 6972 23716 7028 23726
rect 5964 23492 6020 23502
rect 5740 23436 5964 23492
rect 5516 23214 5518 23266
rect 5570 23214 5572 23266
rect 5516 23202 5572 23214
rect 5292 23102 5294 23154
rect 5346 23102 5348 23154
rect 5292 23090 5348 23102
rect 5964 22594 6020 23436
rect 6860 23380 6916 23390
rect 6636 23324 6860 23380
rect 6412 23268 6468 23278
rect 6076 22930 6132 22942
rect 6076 22878 6078 22930
rect 6130 22878 6132 22930
rect 6076 22820 6132 22878
rect 6076 22754 6132 22764
rect 5964 22542 5966 22594
rect 6018 22542 6020 22594
rect 5964 22530 6020 22542
rect 5740 22372 5796 22382
rect 5740 22258 5796 22316
rect 5740 22206 5742 22258
rect 5794 22206 5796 22258
rect 5740 22148 5796 22206
rect 6412 22372 6468 23212
rect 6412 22258 6468 22316
rect 6412 22206 6414 22258
rect 6466 22206 6468 22258
rect 6412 22194 6468 22206
rect 6636 22594 6692 23324
rect 6860 23286 6916 23324
rect 6636 22542 6638 22594
rect 6690 22542 6692 22594
rect 5740 22082 5796 22092
rect 5852 22146 5908 22158
rect 5852 22094 5854 22146
rect 5906 22094 5908 22146
rect 5180 21074 5236 21084
rect 5516 22036 5572 22046
rect 5516 21698 5572 21980
rect 5516 21646 5518 21698
rect 5570 21646 5572 21698
rect 5180 20692 5236 20702
rect 5180 20598 5236 20636
rect 4844 20188 5012 20244
rect 5516 20356 5572 21646
rect 5852 21700 5908 22094
rect 6524 22146 6580 22158
rect 6524 22094 6526 22146
rect 6578 22094 6580 22146
rect 5852 21634 5908 21644
rect 6188 21812 6244 21822
rect 6524 21812 6580 22094
rect 5852 20802 5908 20814
rect 5852 20750 5854 20802
rect 5906 20750 5908 20802
rect 5852 20692 5908 20750
rect 6188 20802 6244 21756
rect 6412 21756 6580 21812
rect 6188 20750 6190 20802
rect 6242 20750 6244 20802
rect 6188 20738 6244 20750
rect 6300 21586 6356 21598
rect 6300 21534 6302 21586
rect 6354 21534 6356 21586
rect 5852 20626 5908 20636
rect 6076 20578 6132 20590
rect 6076 20526 6078 20578
rect 6130 20526 6132 20578
rect 6076 20356 6132 20526
rect 5516 20300 6132 20356
rect 4060 19908 4116 19918
rect 4396 19908 4452 19918
rect 4060 19906 4340 19908
rect 4060 19854 4062 19906
rect 4114 19854 4340 19906
rect 4060 19852 4340 19854
rect 4060 19842 4116 19852
rect 3836 18946 3892 18956
rect 3948 19234 4004 19246
rect 3948 19182 3950 19234
rect 4002 19182 4004 19234
rect 3948 18564 4004 19182
rect 4284 19124 4340 19852
rect 4396 19814 4452 19852
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4844 19236 4900 20188
rect 5404 20132 5460 20142
rect 5404 20038 5460 20076
rect 4956 20020 5012 20030
rect 4956 19926 5012 19964
rect 5292 20018 5348 20030
rect 5292 19966 5294 20018
rect 5346 19966 5348 20018
rect 5292 19236 5348 19966
rect 4844 19180 5012 19236
rect 4396 19124 4452 19134
rect 4284 19122 4452 19124
rect 4284 19070 4398 19122
rect 4450 19070 4452 19122
rect 4284 19068 4452 19070
rect 4172 19010 4228 19022
rect 4172 18958 4174 19010
rect 4226 18958 4228 19010
rect 4172 18676 4228 18958
rect 4172 18610 4228 18620
rect 3836 18452 3892 18462
rect 3724 18450 3892 18452
rect 3724 18398 3838 18450
rect 3890 18398 3892 18450
rect 3724 18396 3892 18398
rect 3836 18386 3892 18396
rect 3612 16830 3614 16882
rect 3666 16830 3668 16882
rect 3612 16818 3668 16830
rect 3724 17666 3780 17678
rect 3724 17614 3726 17666
rect 3778 17614 3780 17666
rect 3724 16212 3780 17614
rect 3836 17668 3892 17678
rect 3836 17442 3892 17612
rect 3836 17390 3838 17442
rect 3890 17390 3892 17442
rect 3836 17378 3892 17390
rect 3948 17444 4004 18508
rect 4060 17444 4116 17454
rect 3948 17442 4228 17444
rect 3948 17390 4062 17442
rect 4114 17390 4228 17442
rect 3948 17388 4228 17390
rect 4060 17378 4116 17388
rect 3836 17108 3892 17118
rect 3836 17014 3892 17052
rect 4060 17108 4116 17118
rect 3948 16996 4004 17006
rect 3724 16146 3780 16156
rect 3836 16884 3892 16894
rect 3612 16100 3668 16110
rect 3612 16006 3668 16044
rect 3836 15874 3892 16828
rect 3836 15822 3838 15874
rect 3890 15822 3892 15874
rect 3836 15810 3892 15822
rect 3612 15764 3668 15774
rect 3500 15708 3612 15764
rect 3612 15698 3668 15708
rect 3948 15540 4004 16940
rect 4060 15874 4116 17052
rect 4172 16100 4228 17388
rect 4284 17108 4340 19068
rect 4396 19058 4452 19068
rect 4844 19012 4900 19022
rect 4844 18918 4900 18956
rect 4508 18564 4564 18574
rect 4508 18470 4564 18508
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4620 17780 4676 17790
rect 4620 17686 4676 17724
rect 4284 17042 4340 17052
rect 4732 17108 4788 17118
rect 4956 17108 5012 19180
rect 5292 19170 5348 19180
rect 5068 18564 5124 18574
rect 5068 18470 5124 18508
rect 5404 18340 5460 18350
rect 5516 18340 5572 20300
rect 6188 20244 6244 20254
rect 5628 20020 5684 20030
rect 5628 19926 5684 19964
rect 6076 19906 6132 19918
rect 6076 19854 6078 19906
rect 6130 19854 6132 19906
rect 6076 19794 6132 19854
rect 6076 19742 6078 19794
rect 6130 19742 6132 19794
rect 6076 19730 6132 19742
rect 5740 19124 5796 19134
rect 5740 19030 5796 19068
rect 5852 18564 5908 18574
rect 5852 18450 5908 18508
rect 5852 18398 5854 18450
rect 5906 18398 5908 18450
rect 5852 18386 5908 18398
rect 5404 18338 5572 18340
rect 5404 18286 5406 18338
rect 5458 18286 5572 18338
rect 5404 18284 5572 18286
rect 5292 17892 5348 17902
rect 4956 17052 5236 17108
rect 4732 17014 4788 17052
rect 4508 16882 4564 16894
rect 4508 16830 4510 16882
rect 4562 16830 4564 16882
rect 4508 16772 4564 16830
rect 4956 16882 5012 16894
rect 4956 16830 4958 16882
rect 5010 16830 5012 16882
rect 4508 16706 4564 16716
rect 4844 16772 4900 16782
rect 4844 16678 4900 16716
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4620 16210 4676 16222
rect 4620 16158 4622 16210
rect 4674 16158 4676 16210
rect 4172 16044 4340 16100
rect 4060 15822 4062 15874
rect 4114 15822 4116 15874
rect 4060 15810 4116 15822
rect 4172 15764 4228 15774
rect 3836 15484 4004 15540
rect 4060 15652 4116 15662
rect 3500 15428 3556 15438
rect 3836 15428 3892 15484
rect 3500 15426 3892 15428
rect 3500 15374 3502 15426
rect 3554 15374 3892 15426
rect 3500 15372 3892 15374
rect 3500 15362 3556 15372
rect 3164 15262 3166 15314
rect 3218 15262 3220 15314
rect 3164 15204 3220 15262
rect 3276 15260 3444 15316
rect 3276 15204 3332 15260
rect 3164 15148 3332 15204
rect 3052 15036 3220 15092
rect 2828 14578 2884 14588
rect 2940 14980 2996 14990
rect 2940 14642 2996 14924
rect 2940 14590 2942 14642
rect 2994 14590 2996 14642
rect 2940 14578 2996 14590
rect 3052 14868 3108 14878
rect 1932 13580 2660 13636
rect 2940 13636 2996 13646
rect 1932 10052 1988 13580
rect 2940 13542 2996 13580
rect 2044 13412 2100 13422
rect 2044 12850 2100 13356
rect 3052 13300 3108 14812
rect 2044 12798 2046 12850
rect 2098 12798 2100 12850
rect 2044 12786 2100 12798
rect 2156 13244 3108 13300
rect 2044 12404 2100 12414
rect 2156 12404 2212 13244
rect 3164 13188 3220 15036
rect 3388 14532 3444 15260
rect 3948 15314 4004 15326
rect 3948 15262 3950 15314
rect 4002 15262 4004 15314
rect 3836 14756 3892 14766
rect 3836 14662 3892 14700
rect 3724 14532 3780 14542
rect 3388 14530 3780 14532
rect 3388 14478 3726 14530
rect 3778 14478 3780 14530
rect 3388 14476 3780 14478
rect 3724 14466 3780 14476
rect 3388 14306 3444 14318
rect 3388 14254 3390 14306
rect 3442 14254 3444 14306
rect 3388 14196 3444 14254
rect 3388 14130 3444 14140
rect 3836 14306 3892 14318
rect 3836 14254 3838 14306
rect 3890 14254 3892 14306
rect 3836 13972 3892 14254
rect 3836 13906 3892 13916
rect 2044 12402 2212 12404
rect 2044 12350 2046 12402
rect 2098 12350 2212 12402
rect 2044 12348 2212 12350
rect 2268 13132 3220 13188
rect 2044 12338 2100 12348
rect 2044 11284 2100 11294
rect 2268 11284 2324 13132
rect 2492 12738 2548 12750
rect 2492 12686 2494 12738
rect 2546 12686 2548 12738
rect 2492 12404 2548 12686
rect 2492 12338 2548 12348
rect 2492 12068 2548 12078
rect 2492 11974 2548 12012
rect 2044 11282 2324 11284
rect 2044 11230 2046 11282
rect 2098 11230 2324 11282
rect 2044 11228 2324 11230
rect 2044 11218 2100 11228
rect 2492 11172 2548 11182
rect 2492 11078 2548 11116
rect 1932 9996 2100 10052
rect 1708 9714 1876 9716
rect 1708 9662 1710 9714
rect 1762 9662 1876 9714
rect 1708 9660 1876 9662
rect 1932 9826 1988 9838
rect 1932 9774 1934 9826
rect 1986 9774 1988 9826
rect 1932 9716 1988 9774
rect 1708 9650 1764 9660
rect 1932 9650 1988 9660
rect 2044 9492 2100 9996
rect 2492 9716 2548 9726
rect 2492 9622 2548 9660
rect 1932 9436 2100 9492
rect 1708 9042 1764 9054
rect 1708 8990 1710 9042
rect 1762 8990 1764 9042
rect 1708 8820 1764 8990
rect 1708 8754 1764 8764
rect 1708 8146 1764 8158
rect 1708 8094 1710 8146
rect 1762 8094 1764 8146
rect 1708 7924 1764 8094
rect 1708 7858 1764 7868
rect 1708 7474 1764 7486
rect 1708 7422 1710 7474
rect 1762 7422 1764 7474
rect 1708 7028 1764 7422
rect 1708 6962 1764 6972
rect 1708 6578 1764 6590
rect 1708 6526 1710 6578
rect 1762 6526 1764 6578
rect 1708 6132 1764 6526
rect 1708 6066 1764 6076
rect 1708 5906 1764 5918
rect 1708 5854 1710 5906
rect 1762 5854 1764 5906
rect 1708 5796 1764 5854
rect 1932 5908 1988 9436
rect 2044 9268 2100 9278
rect 2044 9174 2100 9212
rect 2492 8930 2548 8942
rect 2492 8878 2494 8930
rect 2546 8878 2548 8930
rect 2492 8820 2548 8878
rect 2492 8754 2548 8764
rect 3948 8428 4004 15262
rect 4060 11396 4116 15596
rect 4060 11330 4116 11340
rect 4172 8428 4228 15708
rect 4284 15426 4340 16044
rect 4284 15374 4286 15426
rect 4338 15374 4340 15426
rect 4284 15362 4340 15374
rect 4620 15988 4676 16158
rect 4620 15316 4676 15932
rect 4620 15250 4676 15260
rect 4844 16212 4900 16222
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 3724 8372 4004 8428
rect 4060 8372 4228 8428
rect 2044 8148 2100 8158
rect 2044 8054 2100 8092
rect 2492 8034 2548 8046
rect 2492 7982 2494 8034
rect 2546 7982 2548 8034
rect 2492 7924 2548 7982
rect 2492 7858 2548 7868
rect 2044 7700 2100 7710
rect 2044 7606 2100 7644
rect 2044 7476 2100 7486
rect 2044 6578 2100 7420
rect 2492 7362 2548 7374
rect 2492 7310 2494 7362
rect 2546 7310 2548 7362
rect 2492 7028 2548 7310
rect 2492 6962 2548 6972
rect 2044 6526 2046 6578
rect 2098 6526 2100 6578
rect 2044 6514 2100 6526
rect 2492 6466 2548 6478
rect 2492 6414 2494 6466
rect 2546 6414 2548 6466
rect 2156 6356 2212 6366
rect 2044 6132 2100 6142
rect 2156 6132 2212 6300
rect 2044 6130 2212 6132
rect 2044 6078 2046 6130
rect 2098 6078 2212 6130
rect 2044 6076 2212 6078
rect 2492 6132 2548 6414
rect 3724 6356 3780 8372
rect 4060 7476 4116 8372
rect 4844 7700 4900 16156
rect 4956 15204 5012 16830
rect 5068 16882 5124 16894
rect 5068 16830 5070 16882
rect 5122 16830 5124 16882
rect 5068 16324 5124 16830
rect 5068 16258 5124 16268
rect 5068 16100 5124 16110
rect 5180 16100 5236 17052
rect 5068 16098 5180 16100
rect 5068 16046 5070 16098
rect 5122 16046 5180 16098
rect 5068 16044 5180 16046
rect 5068 16034 5124 16044
rect 5180 16006 5236 16044
rect 4956 15138 5012 15148
rect 5292 14756 5348 17836
rect 5404 17332 5460 18284
rect 5404 17266 5460 17276
rect 5628 16324 5684 16334
rect 5628 15986 5684 16268
rect 5852 16100 5908 16110
rect 5852 16006 5908 16044
rect 5628 15934 5630 15986
rect 5682 15934 5684 15986
rect 5628 15922 5684 15934
rect 6076 15876 6132 15886
rect 6076 15314 6132 15820
rect 6188 15426 6244 20188
rect 6188 15374 6190 15426
rect 6242 15374 6244 15426
rect 6188 15362 6244 15374
rect 6300 15428 6356 21534
rect 6412 21028 6468 21756
rect 6636 21700 6692 22542
rect 6972 22484 7028 23660
rect 6972 22418 7028 22428
rect 6412 20962 6468 20972
rect 6524 21644 6692 21700
rect 6412 19908 6468 19918
rect 6412 19814 6468 19852
rect 6524 19794 6580 21644
rect 6636 21476 6692 21486
rect 6636 20802 6692 21420
rect 6636 20750 6638 20802
rect 6690 20750 6692 20802
rect 6636 20738 6692 20750
rect 6860 20804 6916 20814
rect 6860 20802 7028 20804
rect 6860 20750 6862 20802
rect 6914 20750 7028 20802
rect 6860 20748 7028 20750
rect 6860 20738 6916 20748
rect 6524 19742 6526 19794
rect 6578 19742 6580 19794
rect 6524 19730 6580 19742
rect 6972 19906 7028 20748
rect 6972 19854 6974 19906
rect 7026 19854 7028 19906
rect 6972 19348 7028 19854
rect 6972 19282 7028 19292
rect 6860 17666 6916 17678
rect 6860 17614 6862 17666
rect 6914 17614 6916 17666
rect 6860 16884 6916 17614
rect 7084 17108 7140 31612
rect 7196 30098 7252 33404
rect 7756 33122 7812 33134
rect 7756 33070 7758 33122
rect 7810 33070 7812 33122
rect 7756 33012 7812 33070
rect 7756 32946 7812 32956
rect 7868 32676 7924 33852
rect 7756 32674 7924 32676
rect 7756 32622 7870 32674
rect 7922 32622 7924 32674
rect 7756 32620 7924 32622
rect 7420 31778 7476 31790
rect 7420 31726 7422 31778
rect 7474 31726 7476 31778
rect 7420 31444 7476 31726
rect 7756 31778 7812 32620
rect 7868 32610 7924 32620
rect 7756 31726 7758 31778
rect 7810 31726 7812 31778
rect 7756 31714 7812 31726
rect 7868 31892 7924 31902
rect 7868 31778 7924 31836
rect 7868 31726 7870 31778
rect 7922 31726 7924 31778
rect 7868 31714 7924 31726
rect 7420 31378 7476 31388
rect 7868 31556 7924 31566
rect 7868 31218 7924 31500
rect 7868 31166 7870 31218
rect 7922 31166 7924 31218
rect 7868 31154 7924 31166
rect 7532 30884 7588 30894
rect 7196 30046 7198 30098
rect 7250 30046 7252 30098
rect 7196 28642 7252 30046
rect 7196 28590 7198 28642
rect 7250 28590 7252 28642
rect 7196 28578 7252 28590
rect 7308 30324 7364 30334
rect 7196 27748 7252 27758
rect 7196 27654 7252 27692
rect 7308 27074 7364 30268
rect 7532 27860 7588 30828
rect 8204 30324 8260 34412
rect 8428 34132 8484 34860
rect 8428 34038 8484 34076
rect 8652 35364 8708 35374
rect 8652 35028 8708 35308
rect 8652 33346 8708 34972
rect 8764 34916 8820 34926
rect 8764 34822 8820 34860
rect 8876 34244 8932 34254
rect 9548 34244 9604 37548
rect 8876 34242 9604 34244
rect 8876 34190 8878 34242
rect 8930 34190 9604 34242
rect 8876 34188 9604 34190
rect 8876 34178 8932 34188
rect 9548 34130 9604 34188
rect 9548 34078 9550 34130
rect 9602 34078 9604 34130
rect 8652 33294 8654 33346
rect 8706 33294 8708 33346
rect 8652 33282 8708 33294
rect 8764 34018 8820 34030
rect 8764 33966 8766 34018
rect 8818 33966 8820 34018
rect 8316 32786 8372 32798
rect 8316 32734 8318 32786
rect 8370 32734 8372 32786
rect 8316 32340 8372 32734
rect 8316 32274 8372 32284
rect 8652 31780 8708 31790
rect 8428 31778 8708 31780
rect 8428 31726 8654 31778
rect 8706 31726 8708 31778
rect 8428 31724 8708 31726
rect 8204 30258 8260 30268
rect 8316 31444 8372 31454
rect 7868 30212 7924 30222
rect 7868 29764 7924 30156
rect 8092 29988 8148 29998
rect 8092 29986 8260 29988
rect 8092 29934 8094 29986
rect 8146 29934 8260 29986
rect 8092 29932 8260 29934
rect 8092 29922 8148 29932
rect 7644 29428 7700 29438
rect 7644 28754 7700 29372
rect 7756 29316 7812 29326
rect 7756 29222 7812 29260
rect 7644 28702 7646 28754
rect 7698 28702 7700 28754
rect 7644 28690 7700 28702
rect 7756 28756 7812 28766
rect 7644 27860 7700 27870
rect 7532 27858 7700 27860
rect 7532 27806 7646 27858
rect 7698 27806 7700 27858
rect 7532 27804 7700 27806
rect 7644 27794 7700 27804
rect 7308 27022 7310 27074
rect 7362 27022 7364 27074
rect 7308 26908 7364 27022
rect 7196 26852 7364 26908
rect 7756 26962 7812 28700
rect 7756 26910 7758 26962
rect 7810 26910 7812 26962
rect 7756 26898 7812 26910
rect 7868 27074 7924 29708
rect 8092 28756 8148 28766
rect 8092 28662 8148 28700
rect 7868 27022 7870 27074
rect 7922 27022 7924 27074
rect 7532 26852 7588 26862
rect 7196 26404 7252 26852
rect 7420 26850 7588 26852
rect 7420 26798 7534 26850
rect 7586 26798 7588 26850
rect 7420 26796 7588 26798
rect 7196 26338 7252 26348
rect 7308 26628 7364 26638
rect 7308 25508 7364 26572
rect 7308 25394 7364 25452
rect 7308 25342 7310 25394
rect 7362 25342 7364 25394
rect 7308 25330 7364 25342
rect 7420 25284 7476 26796
rect 7532 26786 7588 26796
rect 7868 26290 7924 27022
rect 7868 26238 7870 26290
rect 7922 26238 7924 26290
rect 7868 26226 7924 26238
rect 7980 28532 8036 28542
rect 7980 26068 8036 28476
rect 8092 27188 8148 27198
rect 8092 26404 8148 27132
rect 8204 26628 8260 29932
rect 8316 29316 8372 31388
rect 8428 31108 8484 31724
rect 8652 31714 8708 31724
rect 8540 31556 8596 31566
rect 8596 31500 8708 31556
rect 8540 31490 8596 31500
rect 8428 31052 8596 31108
rect 8428 30882 8484 30894
rect 8428 30830 8430 30882
rect 8482 30830 8484 30882
rect 8428 30324 8484 30830
rect 8428 30258 8484 30268
rect 8540 29540 8596 31052
rect 8652 30434 8708 31500
rect 8764 30548 8820 33966
rect 9212 33458 9268 33470
rect 9212 33406 9214 33458
rect 9266 33406 9268 33458
rect 8876 31780 8932 31790
rect 8876 31686 8932 31724
rect 8764 30492 8932 30548
rect 8652 30382 8654 30434
rect 8706 30382 8708 30434
rect 8652 30370 8708 30382
rect 8764 30322 8820 30334
rect 8764 30270 8766 30322
rect 8818 30270 8820 30322
rect 8652 30212 8708 30222
rect 8764 30212 8820 30270
rect 8708 30156 8820 30212
rect 8652 30146 8708 30156
rect 8876 29764 8932 30492
rect 8988 30436 9044 30446
rect 8988 30342 9044 30380
rect 9100 30212 9156 30222
rect 9100 30118 9156 30156
rect 8876 29708 9044 29764
rect 8764 29652 8820 29662
rect 8764 29558 8820 29596
rect 8316 27970 8372 29260
rect 8428 29484 8596 29540
rect 8876 29538 8932 29550
rect 8876 29486 8878 29538
rect 8930 29486 8932 29538
rect 8428 28420 8484 29484
rect 8652 29428 8708 29438
rect 8428 28354 8484 28364
rect 8540 29372 8652 29428
rect 8316 27918 8318 27970
rect 8370 27918 8372 27970
rect 8316 27906 8372 27918
rect 8540 27858 8596 29372
rect 8652 29334 8708 29372
rect 8876 29316 8932 29486
rect 8876 29250 8932 29260
rect 8988 28754 9044 29708
rect 9212 28868 9268 33406
rect 9548 33236 9604 34078
rect 9548 33170 9604 33180
rect 9660 32116 9716 38108
rect 9884 38098 9940 38108
rect 11004 38164 11060 38174
rect 11004 38070 11060 38108
rect 11788 38162 11844 38174
rect 11788 38110 11790 38162
rect 11842 38110 11844 38162
rect 10444 37828 10500 37838
rect 9996 37826 10500 37828
rect 9996 37774 10446 37826
rect 10498 37774 10500 37826
rect 9996 37772 10500 37774
rect 9996 37156 10052 37772
rect 10444 37762 10500 37772
rect 9996 36482 10052 37100
rect 9996 36430 9998 36482
rect 10050 36430 10052 36482
rect 9996 36418 10052 36430
rect 10220 37378 10276 37390
rect 11116 37380 11172 37390
rect 10220 37326 10222 37378
rect 10274 37326 10276 37378
rect 10220 37268 10276 37326
rect 11004 37378 11172 37380
rect 11004 37326 11118 37378
rect 11170 37326 11172 37378
rect 11004 37324 11172 37326
rect 10108 35812 10164 35822
rect 9996 35810 10164 35812
rect 9996 35758 10110 35810
rect 10162 35758 10164 35810
rect 9996 35756 10164 35758
rect 9772 34132 9828 34142
rect 9996 34132 10052 35756
rect 10108 35746 10164 35756
rect 9828 34076 10052 34132
rect 10220 34802 10276 37212
rect 10780 37266 10836 37278
rect 10780 37214 10782 37266
rect 10834 37214 10836 37266
rect 10780 35028 10836 37214
rect 11004 37044 11060 37324
rect 11116 37314 11172 37324
rect 11004 36372 11060 36988
rect 11340 37154 11396 37166
rect 11340 37102 11342 37154
rect 11394 37102 11396 37154
rect 11004 36370 11284 36372
rect 11004 36318 11006 36370
rect 11058 36318 11284 36370
rect 11004 36316 11284 36318
rect 11004 36306 11060 36316
rect 11004 35700 11060 35710
rect 11004 35606 11060 35644
rect 11228 35698 11284 36316
rect 11228 35646 11230 35698
rect 11282 35646 11284 35698
rect 11228 35634 11284 35646
rect 10780 34914 10836 34972
rect 10780 34862 10782 34914
rect 10834 34862 10836 34914
rect 10780 34850 10836 34862
rect 10220 34750 10222 34802
rect 10274 34750 10276 34802
rect 9772 34038 9828 34076
rect 10108 33906 10164 33918
rect 10108 33854 10110 33906
rect 10162 33854 10164 33906
rect 10108 33348 10164 33854
rect 9996 32564 10052 32574
rect 10108 32564 10164 33292
rect 10220 33346 10276 34750
rect 10220 33294 10222 33346
rect 10274 33294 10276 33346
rect 10220 33282 10276 33294
rect 10892 34802 10948 34814
rect 10892 34750 10894 34802
rect 10946 34750 10948 34802
rect 10332 33236 10388 33246
rect 10332 33142 10388 33180
rect 10780 33124 10836 33134
rect 10780 32674 10836 33068
rect 10780 32622 10782 32674
rect 10834 32622 10836 32674
rect 10780 32610 10836 32622
rect 9996 32562 10388 32564
rect 9996 32510 9998 32562
rect 10050 32510 10388 32562
rect 9996 32508 10388 32510
rect 9996 32498 10052 32508
rect 10108 32340 10164 32350
rect 9996 32228 10052 32238
rect 9660 32060 9940 32116
rect 9436 31666 9492 31678
rect 9436 31614 9438 31666
rect 9490 31614 9492 31666
rect 9436 30100 9492 31614
rect 9436 30034 9492 30044
rect 9548 31668 9604 31678
rect 9548 29988 9604 31612
rect 9548 29894 9604 29932
rect 9772 31554 9828 31566
rect 9772 31502 9774 31554
rect 9826 31502 9828 31554
rect 9772 29540 9828 31502
rect 9884 30884 9940 32060
rect 9996 31444 10052 32172
rect 10108 32002 10164 32284
rect 10108 31950 10110 32002
rect 10162 31950 10164 32002
rect 10108 31938 10164 31950
rect 10332 31890 10388 32508
rect 10332 31838 10334 31890
rect 10386 31838 10388 31890
rect 10332 31826 10388 31838
rect 10444 32450 10500 32462
rect 10444 32398 10446 32450
rect 10498 32398 10500 32450
rect 9996 31378 10052 31388
rect 10220 30996 10276 31006
rect 10444 30996 10500 32398
rect 10220 30902 10276 30940
rect 10332 30940 10500 30996
rect 10668 31554 10724 31566
rect 10668 31502 10670 31554
rect 10722 31502 10724 31554
rect 9884 30818 9940 30828
rect 9996 30882 10052 30894
rect 9996 30830 9998 30882
rect 10050 30830 10052 30882
rect 9996 30772 10052 30830
rect 10220 30772 10276 30782
rect 9996 30716 10220 30772
rect 9996 30324 10052 30334
rect 9996 30230 10052 30268
rect 9772 29474 9828 29484
rect 9884 30210 9940 30222
rect 9884 30158 9886 30210
rect 9938 30158 9940 30210
rect 9884 30100 9940 30158
rect 9548 29428 9604 29438
rect 8988 28702 8990 28754
rect 9042 28702 9044 28754
rect 8540 27806 8542 27858
rect 8594 27806 8596 27858
rect 8540 27794 8596 27806
rect 8876 28642 8932 28654
rect 8876 28590 8878 28642
rect 8930 28590 8932 28642
rect 8876 28082 8932 28590
rect 8876 28030 8878 28082
rect 8930 28030 8932 28082
rect 8876 26908 8932 28030
rect 8764 26852 8932 26908
rect 8428 26628 8484 26638
rect 8204 26572 8428 26628
rect 8428 26514 8484 26572
rect 8428 26462 8430 26514
rect 8482 26462 8484 26514
rect 8428 26450 8484 26462
rect 8092 26348 8260 26404
rect 8092 26180 8148 26190
rect 8092 26086 8148 26124
rect 7644 26012 8036 26068
rect 7644 25506 7700 26012
rect 7644 25454 7646 25506
rect 7698 25454 7700 25506
rect 7644 25442 7700 25454
rect 7420 25218 7476 25228
rect 7532 25282 7588 25294
rect 7532 25230 7534 25282
rect 7586 25230 7588 25282
rect 7532 24724 7588 25230
rect 7756 25284 7812 25294
rect 7756 25190 7812 25228
rect 7532 24658 7588 24668
rect 7420 24612 7476 24622
rect 7308 23826 7364 23838
rect 7308 23774 7310 23826
rect 7362 23774 7364 23826
rect 7308 21924 7364 23774
rect 7420 23826 7476 24556
rect 8092 24610 8148 24622
rect 8092 24558 8094 24610
rect 8146 24558 8148 24610
rect 7644 24500 7700 24510
rect 7644 23938 7700 24444
rect 8092 24388 8148 24558
rect 8092 24322 8148 24332
rect 7644 23886 7646 23938
rect 7698 23886 7700 23938
rect 7644 23874 7700 23886
rect 7868 24052 7924 24062
rect 7420 23774 7422 23826
rect 7474 23774 7476 23826
rect 7420 23762 7476 23774
rect 7756 23156 7812 23166
rect 7756 23062 7812 23100
rect 7420 23044 7476 23054
rect 7420 22950 7476 22988
rect 7532 22708 7588 22718
rect 7308 21858 7364 21868
rect 7420 22146 7476 22158
rect 7420 22094 7422 22146
rect 7474 22094 7476 22146
rect 7196 21588 7252 21598
rect 7196 20914 7252 21532
rect 7308 21588 7364 21598
rect 7420 21588 7476 22094
rect 7308 21586 7476 21588
rect 7308 21534 7310 21586
rect 7362 21534 7476 21586
rect 7308 21532 7476 21534
rect 7308 21140 7364 21532
rect 7308 21074 7364 21084
rect 7196 20862 7198 20914
rect 7250 20862 7252 20914
rect 7196 20850 7252 20862
rect 7196 20578 7252 20590
rect 7196 20526 7198 20578
rect 7250 20526 7252 20578
rect 7196 20020 7252 20526
rect 7420 20020 7476 20030
rect 7196 20018 7476 20020
rect 7196 19966 7422 20018
rect 7474 19966 7476 20018
rect 7196 19964 7476 19966
rect 7420 19954 7476 19964
rect 7196 19796 7252 19806
rect 7532 19796 7588 22652
rect 7756 20916 7812 20926
rect 7644 20802 7700 20814
rect 7644 20750 7646 20802
rect 7698 20750 7700 20802
rect 7644 20244 7700 20750
rect 7644 20178 7700 20188
rect 7756 20130 7812 20860
rect 7868 20244 7924 23996
rect 8204 23826 8260 26348
rect 8764 26402 8820 26852
rect 8988 26740 9044 28702
rect 9100 28812 9268 28868
rect 9324 29372 9548 29428
rect 9884 29428 9940 30044
rect 9996 29428 10052 29438
rect 9884 29372 9996 29428
rect 9100 26908 9156 28812
rect 9324 28420 9380 29372
rect 9548 29334 9604 29372
rect 9996 29334 10052 29372
rect 9884 28866 9940 28878
rect 9884 28814 9886 28866
rect 9938 28814 9940 28866
rect 9772 28644 9828 28654
rect 9212 28364 9380 28420
rect 9660 28420 9716 28430
rect 9212 27186 9268 28364
rect 9212 27134 9214 27186
rect 9266 27134 9268 27186
rect 9212 27122 9268 27134
rect 9660 26908 9716 28364
rect 9772 27858 9828 28588
rect 9772 27806 9774 27858
rect 9826 27806 9828 27858
rect 9772 27074 9828 27806
rect 9772 27022 9774 27074
rect 9826 27022 9828 27074
rect 9772 27010 9828 27022
rect 9100 26852 9268 26908
rect 9660 26852 9828 26908
rect 8988 26674 9044 26684
rect 8764 26350 8766 26402
rect 8818 26350 8820 26402
rect 8764 26338 8820 26350
rect 8876 26402 8932 26414
rect 8876 26350 8878 26402
rect 8930 26350 8932 26402
rect 8876 26180 8932 26350
rect 9100 26292 9156 26302
rect 8540 26124 8932 26180
rect 8988 26290 9156 26292
rect 8988 26238 9102 26290
rect 9154 26238 9156 26290
rect 8988 26236 9156 26238
rect 8204 23774 8206 23826
rect 8258 23774 8260 23826
rect 8204 23380 8260 23774
rect 8204 23314 8260 23324
rect 8316 24724 8372 24734
rect 8316 23266 8372 24668
rect 8428 23940 8484 23950
rect 8428 23846 8484 23884
rect 8316 23214 8318 23266
rect 8370 23214 8372 23266
rect 8316 23202 8372 23214
rect 8092 23154 8148 23166
rect 8092 23102 8094 23154
rect 8146 23102 8148 23154
rect 8092 22932 8148 23102
rect 7980 22484 8036 22494
rect 8092 22484 8148 22876
rect 7980 22482 8148 22484
rect 7980 22430 7982 22482
rect 8034 22430 8148 22482
rect 7980 22428 8148 22430
rect 8540 22820 8596 26124
rect 8652 25060 8708 25070
rect 8652 24498 8708 25004
rect 8876 24948 8932 24958
rect 8876 24854 8932 24892
rect 8764 24612 8820 24622
rect 8764 24518 8820 24556
rect 8652 24446 8654 24498
rect 8706 24446 8708 24498
rect 8652 23044 8708 24446
rect 8876 23044 8932 23054
rect 8652 22988 8876 23044
rect 7980 22418 8036 22428
rect 8540 22370 8596 22764
rect 8876 22820 8932 22988
rect 8876 22754 8932 22764
rect 8540 22318 8542 22370
rect 8594 22318 8596 22370
rect 8540 22306 8596 22318
rect 8764 22594 8820 22606
rect 8764 22542 8766 22594
rect 8818 22542 8820 22594
rect 8316 21812 8372 21822
rect 8316 21026 8372 21756
rect 8652 21588 8708 21598
rect 8652 21494 8708 21532
rect 8316 20974 8318 21026
rect 8370 20974 8372 21026
rect 8316 20962 8372 20974
rect 8204 20804 8260 20814
rect 8204 20710 8260 20748
rect 7868 20188 8148 20244
rect 7756 20078 7758 20130
rect 7810 20078 7812 20130
rect 7756 20066 7812 20078
rect 7980 20020 8036 20030
rect 7196 19794 7588 19796
rect 7196 19742 7198 19794
rect 7250 19742 7588 19794
rect 7196 19740 7588 19742
rect 7868 20018 8036 20020
rect 7868 19966 7982 20018
rect 8034 19966 8036 20018
rect 7868 19964 8036 19966
rect 7196 19730 7252 19740
rect 7868 18788 7924 19964
rect 7980 19954 8036 19964
rect 8092 18788 8148 20188
rect 8764 20130 8820 22542
rect 8988 22372 9044 26236
rect 9100 26226 9156 26236
rect 9212 25618 9268 26852
rect 9436 26740 9492 26750
rect 9212 25566 9214 25618
rect 9266 25566 9268 25618
rect 9100 25284 9156 25294
rect 9100 23380 9156 25228
rect 9212 24276 9268 25566
rect 9212 24210 9268 24220
rect 9324 26516 9380 26526
rect 9100 23324 9268 23380
rect 9100 23156 9156 23166
rect 9100 23062 9156 23100
rect 8988 22306 9044 22316
rect 9100 20802 9156 20814
rect 9100 20750 9102 20802
rect 9154 20750 9156 20802
rect 8988 20690 9044 20702
rect 8988 20638 8990 20690
rect 9042 20638 9044 20690
rect 8876 20244 8932 20254
rect 8988 20244 9044 20638
rect 8876 20242 9044 20244
rect 8876 20190 8878 20242
rect 8930 20190 9044 20242
rect 8876 20188 9044 20190
rect 8876 20178 8932 20188
rect 8764 20078 8766 20130
rect 8818 20078 8820 20130
rect 8204 19908 8260 19918
rect 8204 19906 8484 19908
rect 8204 19854 8206 19906
rect 8258 19854 8484 19906
rect 8204 19852 8484 19854
rect 8204 19842 8260 19852
rect 7308 18732 7924 18788
rect 7980 18732 8372 18788
rect 7196 17108 7252 17118
rect 7084 17052 7196 17108
rect 7196 17014 7252 17052
rect 7308 17106 7364 18732
rect 7980 18676 8036 18732
rect 7532 18620 8036 18676
rect 7532 18562 7588 18620
rect 7532 18510 7534 18562
rect 7586 18510 7588 18562
rect 7532 18498 7588 18510
rect 7308 17054 7310 17106
rect 7362 17054 7364 17106
rect 7308 17042 7364 17054
rect 7420 18450 7476 18462
rect 7420 18398 7422 18450
rect 7474 18398 7476 18450
rect 6860 16818 6916 16828
rect 7420 16772 7476 18398
rect 7532 18228 7588 18238
rect 7532 18134 7588 18172
rect 8092 17780 8148 17790
rect 7868 16996 7924 17006
rect 7868 16902 7924 16940
rect 8092 16994 8148 17724
rect 8316 17554 8372 18732
rect 8316 17502 8318 17554
rect 8370 17502 8372 17554
rect 8316 17490 8372 17502
rect 8092 16942 8094 16994
rect 8146 16942 8148 16994
rect 8092 16930 8148 16942
rect 8316 17332 8372 17342
rect 7756 16884 7812 16894
rect 7756 16790 7812 16828
rect 8316 16882 8372 17276
rect 8316 16830 8318 16882
rect 8370 16830 8372 16882
rect 8316 16818 8372 16830
rect 7420 16706 7476 16716
rect 7868 16436 7924 16446
rect 7868 16098 7924 16380
rect 7868 16046 7870 16098
rect 7922 16046 7924 16098
rect 7868 16034 7924 16046
rect 8204 15988 8260 15998
rect 8204 15894 8260 15932
rect 7980 15874 8036 15886
rect 7980 15822 7982 15874
rect 8034 15822 8036 15874
rect 7980 15764 8036 15822
rect 7980 15698 8036 15708
rect 6300 15372 6468 15428
rect 6076 15262 6078 15314
rect 6130 15262 6132 15314
rect 6076 15250 6132 15262
rect 6412 15148 6468 15372
rect 5292 14690 5348 14700
rect 6300 15092 6468 15148
rect 6972 15426 7028 15438
rect 6972 15374 6974 15426
rect 7026 15374 7028 15426
rect 6300 9268 6356 15092
rect 6972 13748 7028 15374
rect 7196 15316 7252 15326
rect 7196 15222 7252 15260
rect 6972 13682 7028 13692
rect 8428 11788 8484 19852
rect 8764 18788 8820 20078
rect 8988 20018 9044 20030
rect 8988 19966 8990 20018
rect 9042 19966 9044 20018
rect 8876 19908 8932 19918
rect 8988 19908 9044 19966
rect 8932 19852 9044 19908
rect 9100 19908 9156 20750
rect 8876 19346 8932 19852
rect 9100 19842 9156 19852
rect 8876 19294 8878 19346
rect 8930 19294 8932 19346
rect 8876 19282 8932 19294
rect 9212 18788 9268 23324
rect 9324 19236 9380 26460
rect 9436 23380 9492 26684
rect 9548 26180 9604 26190
rect 9548 25506 9604 26124
rect 9548 25454 9550 25506
rect 9602 25454 9604 25506
rect 9548 24722 9604 25454
rect 9548 24670 9550 24722
rect 9602 24670 9604 24722
rect 9548 24658 9604 24670
rect 9772 24052 9828 26852
rect 9884 25060 9940 28814
rect 9996 26404 10052 26414
rect 9996 25284 10052 26348
rect 9996 25218 10052 25228
rect 9884 24994 9940 25004
rect 9436 23314 9492 23324
rect 9548 23996 9828 24052
rect 9884 24834 9940 24846
rect 9884 24782 9886 24834
rect 9938 24782 9940 24834
rect 9548 20802 9604 23996
rect 9884 23492 9940 24782
rect 10220 24836 10276 30716
rect 10332 30548 10388 30940
rect 10332 30482 10388 30492
rect 10444 30772 10500 30782
rect 10668 30772 10724 31502
rect 10892 30884 10948 34750
rect 11228 33236 11284 33246
rect 11004 32338 11060 32350
rect 11004 32286 11006 32338
rect 11058 32286 11060 32338
rect 11004 32004 11060 32286
rect 11004 31938 11060 31948
rect 11228 32338 11284 33180
rect 11228 32286 11230 32338
rect 11282 32286 11284 32338
rect 11116 31892 11172 31902
rect 10892 30828 11060 30884
rect 10444 30770 10724 30772
rect 10444 30718 10446 30770
rect 10498 30718 10724 30770
rect 10444 30716 10724 30718
rect 10780 30772 10836 30782
rect 10780 30770 10948 30772
rect 10780 30718 10782 30770
rect 10834 30718 10948 30770
rect 10780 30716 10948 30718
rect 10444 30212 10500 30716
rect 10780 30706 10836 30716
rect 10444 30146 10500 30156
rect 10556 30436 10612 30446
rect 10444 29428 10500 29438
rect 10332 29314 10388 29326
rect 10332 29262 10334 29314
rect 10386 29262 10388 29314
rect 10332 29092 10388 29262
rect 10332 29026 10388 29036
rect 10444 28642 10500 29372
rect 10444 28590 10446 28642
rect 10498 28590 10500 28642
rect 10332 28308 10388 28318
rect 10332 26908 10388 28252
rect 10444 27074 10500 28590
rect 10444 27022 10446 27074
rect 10498 27022 10500 27074
rect 10444 27010 10500 27022
rect 10556 27076 10612 30380
rect 10668 29986 10724 29998
rect 10668 29934 10670 29986
rect 10722 29934 10724 29986
rect 10668 29316 10724 29934
rect 10780 29316 10836 29326
rect 10668 29314 10836 29316
rect 10668 29262 10782 29314
rect 10834 29262 10836 29314
rect 10668 29260 10836 29262
rect 10668 28756 10724 29260
rect 10780 29250 10836 29260
rect 10724 28700 10836 28756
rect 10668 28690 10724 28700
rect 10668 27746 10724 27758
rect 10668 27694 10670 27746
rect 10722 27694 10724 27746
rect 10668 27300 10724 27694
rect 10668 27234 10724 27244
rect 10668 27076 10724 27086
rect 10556 27020 10668 27076
rect 10668 27010 10724 27020
rect 10332 26852 10724 26908
rect 10668 24948 10724 26852
rect 10780 26068 10836 28700
rect 10892 26908 10948 30716
rect 11004 30548 11060 30828
rect 11116 30772 11172 31836
rect 11228 31668 11284 32286
rect 11228 31602 11284 31612
rect 11340 31332 11396 37102
rect 11564 36594 11620 36606
rect 11564 36542 11566 36594
rect 11618 36542 11620 36594
rect 11452 33684 11508 33694
rect 11452 33236 11508 33628
rect 11452 33142 11508 33180
rect 11452 32340 11508 32350
rect 11452 32246 11508 32284
rect 11564 31556 11620 36542
rect 11788 35700 11844 38110
rect 12348 38050 12404 38062
rect 12348 37998 12350 38050
rect 12402 37998 12404 38050
rect 12348 36820 12404 37998
rect 12572 38052 12628 41200
rect 15932 38276 15988 41200
rect 15932 38210 15988 38220
rect 17164 38276 17220 38286
rect 17164 38182 17220 38220
rect 12572 37986 12628 37996
rect 13132 38164 13188 38174
rect 13132 38050 13188 38108
rect 13132 37998 13134 38050
rect 13186 37998 13188 38050
rect 13132 37986 13188 37998
rect 13692 38164 13748 38174
rect 13356 37938 13412 37950
rect 13356 37886 13358 37938
rect 13410 37886 13412 37938
rect 11788 35634 11844 35644
rect 11900 36764 12348 36820
rect 11900 36708 11956 36764
rect 12348 36754 12404 36764
rect 12684 37266 12740 37278
rect 12684 37214 12686 37266
rect 12738 37214 12740 37266
rect 11676 35586 11732 35598
rect 11676 35534 11678 35586
rect 11730 35534 11732 35586
rect 11676 31780 11732 35534
rect 11788 34804 11844 34814
rect 11788 34242 11844 34748
rect 11788 34190 11790 34242
rect 11842 34190 11844 34242
rect 11788 34178 11844 34190
rect 11900 34242 11956 36652
rect 11900 34190 11902 34242
rect 11954 34190 11956 34242
rect 11900 34178 11956 34190
rect 12012 36484 12068 36494
rect 12012 34242 12068 36428
rect 12236 36482 12292 36494
rect 12236 36430 12238 36482
rect 12290 36430 12292 36482
rect 12236 35476 12292 36430
rect 12572 35700 12628 35710
rect 12684 35700 12740 37214
rect 13356 37044 13412 37886
rect 13468 37940 13524 37950
rect 13468 37846 13524 37884
rect 13468 37492 13524 37502
rect 13468 37266 13524 37436
rect 13468 37214 13470 37266
rect 13522 37214 13524 37266
rect 13468 37202 13524 37214
rect 13692 37268 13748 38108
rect 14252 38052 14308 38062
rect 14252 37958 14308 37996
rect 15036 38052 15092 38062
rect 15036 37958 15092 37996
rect 13916 37828 13972 37838
rect 13916 37826 14420 37828
rect 13916 37774 13918 37826
rect 13970 37774 14420 37826
rect 13916 37772 14420 37774
rect 13916 37762 13972 37772
rect 13692 37266 13860 37268
rect 13692 37214 13694 37266
rect 13746 37214 13860 37266
rect 13692 37212 13860 37214
rect 13692 37202 13748 37212
rect 13356 36978 13412 36988
rect 12796 36596 12852 36606
rect 12796 36482 12852 36540
rect 12796 36430 12798 36482
rect 12850 36430 12852 36482
rect 12796 36418 12852 36430
rect 12908 36484 12964 36494
rect 12628 35644 12852 35700
rect 12572 35606 12628 35644
rect 12236 34692 12292 35420
rect 12796 34914 12852 35644
rect 12796 34862 12798 34914
rect 12850 34862 12852 34914
rect 12796 34850 12852 34862
rect 12908 34804 12964 36428
rect 13692 36484 13748 36494
rect 13692 35810 13748 36428
rect 13804 36482 13860 37212
rect 14140 37154 14196 37166
rect 14140 37102 14142 37154
rect 14194 37102 14196 37154
rect 13804 36430 13806 36482
rect 13858 36430 13860 36482
rect 13804 36372 13860 36430
rect 13804 36306 13860 36316
rect 13916 37042 13972 37054
rect 13916 36990 13918 37042
rect 13970 36990 13972 37042
rect 13692 35758 13694 35810
rect 13746 35758 13748 35810
rect 13692 35746 13748 35758
rect 12908 34710 12964 34748
rect 12236 34636 12628 34692
rect 12012 34190 12014 34242
rect 12066 34190 12068 34242
rect 12012 34178 12068 34190
rect 12460 34020 12516 34030
rect 12460 33926 12516 33964
rect 11788 33348 11844 33358
rect 11844 33292 12292 33348
rect 11788 33254 11844 33292
rect 12012 33122 12068 33134
rect 12012 33070 12014 33122
rect 12066 33070 12068 33122
rect 12012 32452 12068 33070
rect 12236 32786 12292 33292
rect 12236 32734 12238 32786
rect 12290 32734 12292 32786
rect 12236 32722 12292 32734
rect 12460 32900 12516 32910
rect 12460 32786 12516 32844
rect 12460 32734 12462 32786
rect 12514 32734 12516 32786
rect 12460 32722 12516 32734
rect 12124 32674 12180 32686
rect 12124 32622 12126 32674
rect 12178 32622 12180 32674
rect 12124 32564 12180 32622
rect 12124 32508 12404 32564
rect 12012 32396 12292 32452
rect 11900 32340 11956 32350
rect 11900 32338 12180 32340
rect 11900 32286 11902 32338
rect 11954 32286 12180 32338
rect 11900 32284 12180 32286
rect 11900 32274 11956 32284
rect 11676 31724 11844 31780
rect 11676 31556 11732 31566
rect 11564 31500 11676 31556
rect 11676 31462 11732 31500
rect 11116 30706 11172 30716
rect 11228 31276 11396 31332
rect 11004 30492 11172 30548
rect 11004 30324 11060 30334
rect 11004 29426 11060 30268
rect 11004 29374 11006 29426
rect 11058 29374 11060 29426
rect 11004 28756 11060 29374
rect 11116 28868 11172 30492
rect 11228 29988 11284 31276
rect 11340 31108 11396 31118
rect 11340 30436 11396 31052
rect 11340 30370 11396 30380
rect 11452 30996 11508 31006
rect 11676 30996 11732 31006
rect 11452 30210 11508 30940
rect 11452 30158 11454 30210
rect 11506 30158 11508 30210
rect 11452 30146 11508 30158
rect 11564 30994 11732 30996
rect 11564 30942 11678 30994
rect 11730 30942 11732 30994
rect 11564 30940 11732 30942
rect 11228 29932 11508 29988
rect 11228 29316 11284 29326
rect 11228 29222 11284 29260
rect 11340 29204 11396 29214
rect 11116 28812 11284 28868
rect 11060 28700 11172 28756
rect 11004 28690 11060 28700
rect 11116 27858 11172 28700
rect 11228 28308 11284 28812
rect 11228 28242 11284 28252
rect 11116 27806 11118 27858
rect 11170 27806 11172 27858
rect 11116 27794 11172 27806
rect 11228 28082 11284 28094
rect 11228 28030 11230 28082
rect 11282 28030 11284 28082
rect 11228 27300 11284 28030
rect 11340 27858 11396 29148
rect 11452 28644 11508 29932
rect 11452 28550 11508 28588
rect 11564 28532 11620 30940
rect 11676 30930 11732 30940
rect 11676 29314 11732 29326
rect 11676 29262 11678 29314
rect 11730 29262 11732 29314
rect 11676 29204 11732 29262
rect 11676 29138 11732 29148
rect 11564 28466 11620 28476
rect 11340 27806 11342 27858
rect 11394 27806 11396 27858
rect 11340 27794 11396 27806
rect 11116 27244 11284 27300
rect 11340 27300 11396 27310
rect 10892 26852 11060 26908
rect 10780 26002 10836 26012
rect 10892 26178 10948 26190
rect 10892 26126 10894 26178
rect 10946 26126 10948 26178
rect 10668 24892 10836 24948
rect 10220 24780 10612 24836
rect 10220 24610 10276 24622
rect 10220 24558 10222 24610
rect 10274 24558 10276 24610
rect 9996 24276 10052 24286
rect 10052 24220 10164 24276
rect 9996 24210 10052 24220
rect 9884 23426 9940 23436
rect 10108 23938 10164 24220
rect 10108 23886 10110 23938
rect 10162 23886 10164 23938
rect 9660 23156 9716 23166
rect 9716 23100 10052 23156
rect 9660 23090 9716 23100
rect 9772 22932 9828 22942
rect 9772 22370 9828 22876
rect 9772 22318 9774 22370
rect 9826 22318 9828 22370
rect 9772 22306 9828 22318
rect 9996 21810 10052 23100
rect 10108 23042 10164 23886
rect 10220 23604 10276 24558
rect 10220 23538 10276 23548
rect 10332 23826 10388 23838
rect 10332 23774 10334 23826
rect 10386 23774 10388 23826
rect 10220 23268 10276 23278
rect 10220 23154 10276 23212
rect 10220 23102 10222 23154
rect 10274 23102 10276 23154
rect 10220 23090 10276 23102
rect 10108 22990 10110 23042
rect 10162 22990 10164 23042
rect 10108 22932 10164 22990
rect 10108 22876 10276 22932
rect 10220 22370 10276 22876
rect 10220 22318 10222 22370
rect 10274 22318 10276 22370
rect 10220 22306 10276 22318
rect 9996 21758 9998 21810
rect 10050 21758 10052 21810
rect 9996 21746 10052 21758
rect 10108 22148 10164 22158
rect 10108 21810 10164 22092
rect 10108 21758 10110 21810
rect 10162 21758 10164 21810
rect 10108 21746 10164 21758
rect 9548 20750 9550 20802
rect 9602 20750 9604 20802
rect 9548 20738 9604 20750
rect 9660 21698 9716 21710
rect 9660 21646 9662 21698
rect 9714 21646 9716 21698
rect 9660 21588 9716 21646
rect 9660 20804 9716 21532
rect 9884 21588 9940 21598
rect 9884 21586 10052 21588
rect 9884 21534 9886 21586
rect 9938 21534 10052 21586
rect 9884 21532 10052 21534
rect 9884 21522 9940 21532
rect 9660 20748 9940 20804
rect 9772 20580 9828 20590
rect 9660 20524 9772 20580
rect 9548 19236 9604 19246
rect 9324 19180 9548 19236
rect 9548 19142 9604 19180
rect 9324 19012 9380 19022
rect 9324 18918 9380 18956
rect 8764 18722 8820 18732
rect 8988 18732 9268 18788
rect 8876 18676 8932 18686
rect 8764 17668 8820 17678
rect 8764 17574 8820 17612
rect 8652 17108 8708 17118
rect 8652 17014 8708 17052
rect 8540 15876 8596 15886
rect 8540 15782 8596 15820
rect 8652 15764 8708 15774
rect 8652 15538 8708 15708
rect 8652 15486 8654 15538
rect 8706 15486 8708 15538
rect 8652 15474 8708 15486
rect 8092 11732 8484 11788
rect 8092 11620 8148 11732
rect 8092 11554 8148 11564
rect 8876 11508 8932 18620
rect 8988 18452 9044 18732
rect 8988 18358 9044 18396
rect 8988 17108 9044 17118
rect 8988 17014 9044 17052
rect 8988 16884 9044 16894
rect 8988 15986 9044 16828
rect 8988 15934 8990 15986
rect 9042 15934 9044 15986
rect 8988 15922 9044 15934
rect 8988 15540 9044 15550
rect 9100 15540 9156 18732
rect 9548 18676 9604 18686
rect 9436 18620 9548 18676
rect 9436 17554 9492 18620
rect 9548 18610 9604 18620
rect 9548 18452 9604 18462
rect 9548 18358 9604 18396
rect 9436 17502 9438 17554
rect 9490 17502 9492 17554
rect 9436 17490 9492 17502
rect 9660 17556 9716 20524
rect 9772 20486 9828 20524
rect 9772 20244 9828 20254
rect 9772 19684 9828 20188
rect 9884 20132 9940 20748
rect 9884 19906 9940 20076
rect 9884 19854 9886 19906
rect 9938 19854 9940 19906
rect 9884 19842 9940 19854
rect 9772 19628 9940 19684
rect 9772 19010 9828 19022
rect 9772 18958 9774 19010
rect 9826 18958 9828 19010
rect 9772 18452 9828 18958
rect 9772 18386 9828 18396
rect 9884 17778 9940 19628
rect 9884 17726 9886 17778
rect 9938 17726 9940 17778
rect 9884 17714 9940 17726
rect 9660 17500 9940 17556
rect 9660 17108 9716 17118
rect 9660 16882 9716 17052
rect 9660 16830 9662 16882
rect 9714 16830 9716 16882
rect 9660 16818 9716 16830
rect 9436 16436 9492 16446
rect 9212 15988 9268 15998
rect 9212 15894 9268 15932
rect 8988 15538 9156 15540
rect 8988 15486 8990 15538
rect 9042 15486 9156 15538
rect 8988 15484 9156 15486
rect 8988 15474 9044 15484
rect 9100 15148 9156 15484
rect 9436 15316 9492 16380
rect 9548 16100 9604 16110
rect 9548 16098 9716 16100
rect 9548 16046 9550 16098
rect 9602 16046 9716 16098
rect 9548 16044 9716 16046
rect 9548 16034 9604 16044
rect 9548 15316 9604 15326
rect 9436 15314 9604 15316
rect 9436 15262 9550 15314
rect 9602 15262 9604 15314
rect 9436 15260 9604 15262
rect 9548 15250 9604 15260
rect 9660 15148 9716 16044
rect 9884 15986 9940 17500
rect 9996 16772 10052 21532
rect 10220 20690 10276 20702
rect 10220 20638 10222 20690
rect 10274 20638 10276 20690
rect 10220 20468 10276 20638
rect 10108 20412 10220 20468
rect 10108 18452 10164 20412
rect 10220 20402 10276 20412
rect 10332 20244 10388 23774
rect 10444 23492 10500 23502
rect 10444 22482 10500 23436
rect 10444 22430 10446 22482
rect 10498 22430 10500 22482
rect 10444 22418 10500 22430
rect 10556 21812 10612 24780
rect 10668 24724 10724 24734
rect 10668 24630 10724 24668
rect 10780 24388 10836 24892
rect 10668 24332 10836 24388
rect 10668 22036 10724 24332
rect 10780 24164 10836 24174
rect 10780 24050 10836 24108
rect 10780 23998 10782 24050
rect 10834 23998 10836 24050
rect 10780 23986 10836 23998
rect 10668 21970 10724 21980
rect 10780 23380 10836 23390
rect 10556 21756 10724 21812
rect 10444 21586 10500 21598
rect 10444 21534 10446 21586
rect 10498 21534 10500 21586
rect 10444 20802 10500 21534
rect 10444 20750 10446 20802
rect 10498 20750 10500 20802
rect 10444 20580 10500 20750
rect 10444 20514 10500 20524
rect 10556 21588 10612 21598
rect 10108 18358 10164 18396
rect 10220 20188 10388 20244
rect 10444 20356 10500 20366
rect 10220 17108 10276 20188
rect 10332 20020 10388 20030
rect 10444 20020 10500 20300
rect 10556 20242 10612 21532
rect 10556 20190 10558 20242
rect 10610 20190 10612 20242
rect 10556 20178 10612 20190
rect 10332 20018 10500 20020
rect 10332 19966 10334 20018
rect 10386 19966 10500 20018
rect 10332 19964 10500 19966
rect 10332 19012 10388 19964
rect 10332 18946 10388 18956
rect 10444 19010 10500 19022
rect 10444 18958 10446 19010
rect 10498 18958 10500 19010
rect 10332 17108 10388 17118
rect 10220 17106 10388 17108
rect 10220 17054 10334 17106
rect 10386 17054 10388 17106
rect 10220 17052 10388 17054
rect 10332 17042 10388 17052
rect 9996 16678 10052 16716
rect 10108 16996 10164 17006
rect 9884 15934 9886 15986
rect 9938 15934 9940 15986
rect 9884 15316 9940 15934
rect 9996 15988 10052 15998
rect 10108 15988 10164 16940
rect 10444 16884 10500 18958
rect 10556 18676 10612 18686
rect 10556 18582 10612 18620
rect 10556 17890 10612 17902
rect 10556 17838 10558 17890
rect 10610 17838 10612 17890
rect 10556 17444 10612 17838
rect 10668 17668 10724 21756
rect 10780 20804 10836 23324
rect 10892 21364 10948 26126
rect 11004 26180 11060 26852
rect 11004 25732 11060 26124
rect 11004 25666 11060 25676
rect 11004 25506 11060 25518
rect 11004 25454 11006 25506
rect 11058 25454 11060 25506
rect 11004 22484 11060 25454
rect 11116 23380 11172 27244
rect 11228 27076 11284 27086
rect 11228 23940 11284 27020
rect 11228 23874 11284 23884
rect 11340 23380 11396 27244
rect 11676 27298 11732 27310
rect 11676 27246 11678 27298
rect 11730 27246 11732 27298
rect 11564 26292 11620 26302
rect 11564 26198 11620 26236
rect 11676 24948 11732 27246
rect 11788 27074 11844 31724
rect 12012 31556 12068 31566
rect 12012 31462 12068 31500
rect 12124 30994 12180 32284
rect 12124 30942 12126 30994
rect 12178 30942 12180 30994
rect 12124 30930 12180 30942
rect 11900 30100 11956 30110
rect 11900 30006 11956 30044
rect 12236 29988 12292 32396
rect 12348 31892 12404 32508
rect 12348 31826 12404 31836
rect 12348 31554 12404 31566
rect 12348 31502 12350 31554
rect 12402 31502 12404 31554
rect 12348 30996 12404 31502
rect 12348 30930 12404 30940
rect 12572 30772 12628 34636
rect 13692 34690 13748 34702
rect 13692 34638 13694 34690
rect 13746 34638 13748 34690
rect 13580 34020 13636 34030
rect 13580 33346 13636 33964
rect 13580 33294 13582 33346
rect 13634 33294 13636 33346
rect 13580 33282 13636 33294
rect 13580 33124 13636 33134
rect 13580 32786 13636 33068
rect 13580 32734 13582 32786
rect 13634 32734 13636 32786
rect 12796 32562 12852 32574
rect 12796 32510 12798 32562
rect 12850 32510 12852 32562
rect 12796 31892 12852 32510
rect 13580 32452 13636 32734
rect 13692 32788 13748 34638
rect 13804 34132 13860 34142
rect 13916 34132 13972 36990
rect 14140 36708 14196 37102
rect 14140 36642 14196 36652
rect 14252 36932 14308 36942
rect 14252 36594 14308 36876
rect 14252 36542 14254 36594
rect 14306 36542 14308 36594
rect 14028 36484 14084 36494
rect 14028 36390 14084 36428
rect 14252 36148 14308 36542
rect 14252 36082 14308 36092
rect 13804 34130 13916 34132
rect 13804 34078 13806 34130
rect 13858 34078 13916 34130
rect 13804 34076 13916 34078
rect 13804 34066 13860 34076
rect 13916 34038 13972 34076
rect 14028 35586 14084 35598
rect 14028 35534 14030 35586
rect 14082 35534 14084 35586
rect 14028 33572 14084 35534
rect 14252 35028 14308 35038
rect 14252 34934 14308 34972
rect 14140 33908 14196 33918
rect 14140 33814 14196 33852
rect 14028 33506 14084 33516
rect 14028 33346 14084 33358
rect 14028 33294 14030 33346
rect 14082 33294 14084 33346
rect 14028 32788 14084 33294
rect 14364 33124 14420 37772
rect 14588 37826 14644 37838
rect 14588 37774 14590 37826
rect 14642 37774 14644 37826
rect 14588 36932 14644 37774
rect 14700 37492 14756 37502
rect 14700 37398 14756 37436
rect 15260 37154 15316 37166
rect 15260 37102 15262 37154
rect 15314 37102 15316 37154
rect 15260 37044 15316 37102
rect 19292 37156 19348 41200
rect 22652 38276 22708 41200
rect 22652 38210 22708 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 19516 38052 19572 38062
rect 19516 37958 19572 37996
rect 19964 38052 20020 38062
rect 24556 38052 24612 38062
rect 19964 37958 20020 37996
rect 23660 38050 24612 38052
rect 23660 37998 24558 38050
rect 24610 37998 24612 38050
rect 23660 37996 24612 37998
rect 21308 37940 21364 37950
rect 21308 37846 21364 37884
rect 20972 37828 21028 37838
rect 20972 37734 21028 37772
rect 21644 37828 21700 37838
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 21644 37266 21700 37772
rect 23660 37490 23716 37996
rect 24556 37986 24612 37996
rect 23660 37438 23662 37490
rect 23714 37438 23716 37490
rect 23660 37426 23716 37438
rect 26012 37492 26068 41200
rect 29372 41076 29428 41200
rect 29708 41188 29764 41244
rect 29596 41132 29764 41188
rect 29596 41076 29652 41132
rect 29372 41020 29652 41076
rect 30044 38274 30100 41244
rect 32704 41200 32816 42000
rect 36064 41200 36176 42000
rect 39424 41200 39536 42000
rect 30044 38222 30046 38274
rect 30098 38222 30100 38274
rect 30044 38210 30100 38222
rect 32732 38276 32788 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 32732 38210 32788 38220
rect 33852 38276 33908 38286
rect 33852 38182 33908 38220
rect 36092 38276 36148 41200
rect 36092 38210 36148 38220
rect 37324 38276 37380 38286
rect 37324 38182 37380 38220
rect 28700 38052 28756 38062
rect 26012 37426 26068 37436
rect 27244 37492 27300 37502
rect 27244 37398 27300 37436
rect 25900 37378 25956 37390
rect 25900 37326 25902 37378
rect 25954 37326 25956 37378
rect 23324 37268 23380 37278
rect 21644 37214 21646 37266
rect 21698 37214 21700 37266
rect 21644 37202 21700 37214
rect 23212 37266 23380 37268
rect 23212 37214 23326 37266
rect 23378 37214 23380 37266
rect 23212 37212 23380 37214
rect 19740 37156 19796 37166
rect 19292 37154 19796 37156
rect 19292 37102 19742 37154
rect 19794 37102 19796 37154
rect 19292 37100 19796 37102
rect 19740 37090 19796 37100
rect 15260 36988 15652 37044
rect 14588 36876 14756 36932
rect 14700 36484 14756 36876
rect 14700 36418 14756 36428
rect 15148 36820 15204 36830
rect 15148 36482 15204 36764
rect 15260 36708 15316 36718
rect 15260 36596 15316 36652
rect 15260 36594 15540 36596
rect 15260 36542 15262 36594
rect 15314 36542 15540 36594
rect 15260 36540 15540 36542
rect 15260 36530 15316 36540
rect 15148 36430 15150 36482
rect 15202 36430 15204 36482
rect 15148 36418 15204 36430
rect 14588 36372 14644 36382
rect 14588 35698 14644 36316
rect 15260 36372 15316 36382
rect 15260 36278 15316 36316
rect 14588 35646 14590 35698
rect 14642 35646 14644 35698
rect 14588 35634 14644 35646
rect 14700 36258 14756 36270
rect 14700 36206 14702 36258
rect 14754 36206 14756 36258
rect 14700 35308 14756 36206
rect 14588 35252 14756 35308
rect 14588 33684 14644 35252
rect 15484 34802 15540 36540
rect 15596 36148 15652 36988
rect 16716 36596 16772 36606
rect 16604 36594 16772 36596
rect 16604 36542 16718 36594
rect 16770 36542 16772 36594
rect 16604 36540 16772 36542
rect 16380 36482 16436 36494
rect 16380 36430 16382 36482
rect 16434 36430 16436 36482
rect 15596 36082 15652 36092
rect 16044 36148 16100 36158
rect 16044 35812 16100 36092
rect 16156 35812 16212 35822
rect 16044 35810 16212 35812
rect 16044 35758 16158 35810
rect 16210 35758 16212 35810
rect 16044 35756 16212 35758
rect 16044 34914 16100 35756
rect 16156 35746 16212 35756
rect 16044 34862 16046 34914
rect 16098 34862 16100 34914
rect 16044 34850 16100 34862
rect 16380 34916 16436 36430
rect 16380 34822 16436 34860
rect 16492 35364 16548 35374
rect 15484 34750 15486 34802
rect 15538 34750 15540 34802
rect 15484 34738 15540 34750
rect 16492 34356 16548 35308
rect 16380 34300 16548 34356
rect 14700 34132 14756 34170
rect 14700 33796 14756 34076
rect 16044 34132 16100 34142
rect 16044 34038 16100 34076
rect 15260 34020 15316 34030
rect 15708 34020 15764 34030
rect 15260 34018 15652 34020
rect 15260 33966 15262 34018
rect 15314 33966 15652 34018
rect 15260 33964 15652 33966
rect 15260 33954 15316 33964
rect 15148 33908 15204 33918
rect 14700 33740 15092 33796
rect 14588 33628 14980 33684
rect 14700 33124 14756 33134
rect 14364 33122 14756 33124
rect 14364 33070 14702 33122
rect 14754 33070 14756 33122
rect 14364 33068 14756 33070
rect 14028 32732 14308 32788
rect 13692 32722 13748 32732
rect 14140 32564 14196 32574
rect 14140 32470 14196 32508
rect 13580 32396 13972 32452
rect 12796 31826 12852 31836
rect 13244 31892 13300 31902
rect 13020 31780 13076 31790
rect 13020 31218 13076 31724
rect 13020 31166 13022 31218
rect 13074 31166 13076 31218
rect 13020 31154 13076 31166
rect 13244 31106 13300 31836
rect 13916 31778 13972 32396
rect 14252 32340 14308 32732
rect 13916 31726 13918 31778
rect 13970 31726 13972 31778
rect 13916 31714 13972 31726
rect 14140 32284 14308 32340
rect 14588 32452 14644 33068
rect 14700 33058 14756 33068
rect 13244 31054 13246 31106
rect 13298 31054 13300 31106
rect 13244 31042 13300 31054
rect 13356 31556 13412 31566
rect 12348 30716 12628 30772
rect 12908 30994 12964 31006
rect 12908 30942 12910 30994
rect 12962 30942 12964 30994
rect 12908 30884 12964 30942
rect 12348 30098 12404 30716
rect 12348 30046 12350 30098
rect 12402 30046 12404 30098
rect 12348 30034 12404 30046
rect 12460 30212 12516 30222
rect 12460 30098 12516 30156
rect 12460 30046 12462 30098
rect 12514 30046 12516 30098
rect 12460 30034 12516 30046
rect 12572 30098 12628 30110
rect 12572 30046 12574 30098
rect 12626 30046 12628 30098
rect 12124 29764 12180 29774
rect 11900 29428 11956 29438
rect 11900 29334 11956 29372
rect 12124 29426 12180 29708
rect 12124 29374 12126 29426
rect 12178 29374 12180 29426
rect 12124 29362 12180 29374
rect 12236 29428 12292 29932
rect 12572 29876 12628 30046
rect 12908 29988 12964 30828
rect 12572 29810 12628 29820
rect 12684 29932 12964 29988
rect 12684 29540 12740 29932
rect 13244 29764 13300 29774
rect 12572 29484 12740 29540
rect 12796 29540 12852 29550
rect 12348 29428 12404 29438
rect 12236 29426 12404 29428
rect 12236 29374 12350 29426
rect 12402 29374 12404 29426
rect 12236 29372 12404 29374
rect 12348 29362 12404 29372
rect 12012 29316 12068 29326
rect 12012 29222 12068 29260
rect 12460 29092 12516 29102
rect 11900 28756 11956 28766
rect 11900 28662 11956 28700
rect 12460 28756 12516 29036
rect 12236 28420 12292 28430
rect 12236 27970 12292 28364
rect 12236 27918 12238 27970
rect 12290 27918 12292 27970
rect 12236 27906 12292 27918
rect 12460 27858 12516 28700
rect 12460 27806 12462 27858
rect 12514 27806 12516 27858
rect 12460 27794 12516 27806
rect 12572 27636 12628 29484
rect 12796 29204 12852 29484
rect 13244 29426 13300 29708
rect 13244 29374 13246 29426
rect 13298 29374 13300 29426
rect 13244 29316 13300 29374
rect 13244 29250 13300 29260
rect 12460 27580 12628 27636
rect 12684 29148 12852 29204
rect 11788 27022 11790 27074
rect 11842 27022 11844 27074
rect 11788 26964 11844 27022
rect 11788 26898 11844 26908
rect 12348 27186 12404 27198
rect 12348 27134 12350 27186
rect 12402 27134 12404 27186
rect 12124 26516 12180 26526
rect 11788 25508 11844 25518
rect 11788 25414 11844 25452
rect 11676 24882 11732 24892
rect 11788 24834 11844 24846
rect 11788 24782 11790 24834
rect 11842 24782 11844 24834
rect 11788 24162 11844 24782
rect 12124 24276 12180 26460
rect 12348 24388 12404 27134
rect 12348 24322 12404 24332
rect 11788 24110 11790 24162
rect 11842 24110 11844 24162
rect 11788 24098 11844 24110
rect 11900 24220 12180 24276
rect 11676 23940 11732 23950
rect 11676 23938 11844 23940
rect 11676 23886 11678 23938
rect 11730 23886 11844 23938
rect 11676 23884 11844 23886
rect 11676 23874 11732 23884
rect 11116 23314 11172 23324
rect 11228 23324 11396 23380
rect 11452 23492 11508 23502
rect 11116 23044 11172 23054
rect 11116 22950 11172 22988
rect 11228 22932 11284 23324
rect 11228 22866 11284 22876
rect 11340 23156 11396 23166
rect 11004 22418 11060 22428
rect 11004 22148 11060 22158
rect 11004 21586 11060 22092
rect 11004 21534 11006 21586
rect 11058 21534 11060 21586
rect 11004 21522 11060 21534
rect 11228 21364 11284 21374
rect 10892 21308 11228 21364
rect 11228 21298 11284 21308
rect 11228 21028 11284 21038
rect 10780 20748 11060 20804
rect 10780 20580 10836 20590
rect 10780 20486 10836 20524
rect 10780 20132 10836 20142
rect 10780 20038 10836 20076
rect 10892 20018 10948 20030
rect 10892 19966 10894 20018
rect 10946 19966 10948 20018
rect 10780 19124 10836 19134
rect 10780 19030 10836 19068
rect 10892 19012 10948 19966
rect 11004 19348 11060 20748
rect 11228 19684 11284 20972
rect 11340 20020 11396 23100
rect 11452 20802 11508 23436
rect 11564 22148 11620 22158
rect 11564 21698 11620 22092
rect 11676 21812 11732 21822
rect 11676 21718 11732 21756
rect 11564 21646 11566 21698
rect 11618 21646 11620 21698
rect 11564 21634 11620 21646
rect 11452 20750 11454 20802
rect 11506 20750 11508 20802
rect 11452 20738 11508 20750
rect 11564 21364 11620 21374
rect 11564 20578 11620 21308
rect 11676 21364 11732 21374
rect 11788 21364 11844 23884
rect 11676 21362 11844 21364
rect 11676 21310 11678 21362
rect 11730 21310 11844 21362
rect 11676 21308 11844 21310
rect 11676 21298 11732 21308
rect 11788 20580 11844 20590
rect 11564 20526 11566 20578
rect 11618 20526 11620 20578
rect 11452 20020 11508 20030
rect 11340 20018 11508 20020
rect 11340 19966 11454 20018
rect 11506 19966 11508 20018
rect 11340 19964 11508 19966
rect 11452 19954 11508 19964
rect 11228 19628 11508 19684
rect 11340 19460 11396 19470
rect 11340 19348 11396 19404
rect 11004 19292 11396 19348
rect 11004 19234 11060 19292
rect 11004 19182 11006 19234
rect 11058 19182 11060 19234
rect 11004 19170 11060 19182
rect 11340 19234 11396 19292
rect 11340 19182 11342 19234
rect 11394 19182 11396 19234
rect 11228 19124 11284 19134
rect 11116 19068 11228 19124
rect 11004 19012 11060 19022
rect 10892 18956 11004 19012
rect 10780 18900 10836 18910
rect 10836 18844 10948 18900
rect 10780 18834 10836 18844
rect 10668 17612 10836 17668
rect 10668 17444 10724 17454
rect 10556 17442 10724 17444
rect 10556 17390 10670 17442
rect 10722 17390 10724 17442
rect 10556 17388 10724 17390
rect 10668 17378 10724 17388
rect 10668 17108 10724 17118
rect 10444 16818 10500 16828
rect 10556 16994 10612 17006
rect 10556 16942 10558 16994
rect 10610 16942 10612 16994
rect 10444 16100 10500 16110
rect 10444 16006 10500 16044
rect 9996 15986 10164 15988
rect 9996 15934 9998 15986
rect 10050 15934 10164 15986
rect 9996 15932 10164 15934
rect 9996 15922 10052 15932
rect 9996 15316 10052 15326
rect 9884 15314 10052 15316
rect 9884 15262 9998 15314
rect 10050 15262 10052 15314
rect 9884 15260 10052 15262
rect 9996 15250 10052 15260
rect 9100 15092 9380 15148
rect 9324 14642 9380 15092
rect 9324 14590 9326 14642
rect 9378 14590 9380 14642
rect 9324 14578 9380 14590
rect 9548 15092 9716 15148
rect 9548 14308 9604 15092
rect 10108 14644 10164 15932
rect 10220 15988 10276 15998
rect 10220 15894 10276 15932
rect 10556 15764 10612 16942
rect 10668 16994 10724 17052
rect 10668 16942 10670 16994
rect 10722 16942 10724 16994
rect 10668 16930 10724 16942
rect 10556 15698 10612 15708
rect 10668 16772 10724 16782
rect 10668 15314 10724 16716
rect 10668 15262 10670 15314
rect 10722 15262 10724 15314
rect 10668 15148 10724 15262
rect 10332 15092 10724 15148
rect 10780 16100 10836 17612
rect 10780 15876 10836 16044
rect 10220 14644 10276 14654
rect 10108 14642 10276 14644
rect 10108 14590 10222 14642
rect 10274 14590 10276 14642
rect 10108 14588 10276 14590
rect 10220 14578 10276 14588
rect 9884 14308 9940 14318
rect 9548 14252 9884 14308
rect 9884 14214 9940 14252
rect 10332 13972 10388 15092
rect 10780 14754 10836 15820
rect 10892 15764 10948 18844
rect 11004 18450 11060 18956
rect 11004 18398 11006 18450
rect 11058 18398 11060 18450
rect 11004 18386 11060 18398
rect 11004 17444 11060 17454
rect 11004 16210 11060 17388
rect 11004 16158 11006 16210
rect 11058 16158 11060 16210
rect 11004 16146 11060 16158
rect 10892 15708 11060 15764
rect 10892 15540 10948 15550
rect 10892 15446 10948 15484
rect 10780 14702 10782 14754
rect 10834 14702 10836 14754
rect 10780 14642 10836 14702
rect 10780 14590 10782 14642
rect 10834 14590 10836 14642
rect 10780 14578 10836 14590
rect 11004 15428 11060 15708
rect 10332 13878 10388 13916
rect 11004 13970 11060 15372
rect 11116 15148 11172 19068
rect 11228 19058 11284 19068
rect 11340 18004 11396 19182
rect 11228 17892 11284 17902
rect 11340 17892 11396 17948
rect 11228 17890 11396 17892
rect 11228 17838 11230 17890
rect 11282 17838 11396 17890
rect 11228 17836 11396 17838
rect 11228 17826 11284 17836
rect 11228 17668 11284 17678
rect 11284 17612 11396 17668
rect 11228 17574 11284 17612
rect 11228 16996 11284 17006
rect 11228 16902 11284 16940
rect 11340 16100 11396 17612
rect 11452 16996 11508 19628
rect 11564 18562 11620 20526
rect 11676 20578 11844 20580
rect 11676 20526 11790 20578
rect 11842 20526 11844 20578
rect 11676 20524 11844 20526
rect 11676 20130 11732 20524
rect 11788 20514 11844 20524
rect 11900 20132 11956 24220
rect 12460 24164 12516 27580
rect 12684 26908 12740 29148
rect 13132 29092 13188 29102
rect 13356 29092 13412 31500
rect 14140 31108 14196 32284
rect 14140 31042 14196 31052
rect 14252 31554 14308 31566
rect 14252 31502 14254 31554
rect 14306 31502 14308 31554
rect 13692 30996 13748 31006
rect 13580 29986 13636 29998
rect 13580 29934 13582 29986
rect 13634 29934 13636 29986
rect 13580 29764 13636 29934
rect 13580 29698 13636 29708
rect 13692 29540 13748 30940
rect 14140 30770 14196 30782
rect 14140 30718 14142 30770
rect 14194 30718 14196 30770
rect 14140 30210 14196 30718
rect 14252 30436 14308 31502
rect 14364 30882 14420 30894
rect 14364 30830 14366 30882
rect 14418 30830 14420 30882
rect 14364 30770 14420 30830
rect 14364 30718 14366 30770
rect 14418 30718 14420 30770
rect 14364 30706 14420 30718
rect 14252 30370 14308 30380
rect 14140 30158 14142 30210
rect 14194 30158 14196 30210
rect 13692 29474 13748 29484
rect 13916 29540 13972 29550
rect 13580 29316 13636 29326
rect 12908 27748 12964 27758
rect 12796 27634 12852 27646
rect 12796 27582 12798 27634
rect 12850 27582 12852 27634
rect 12796 27076 12852 27582
rect 12796 27010 12852 27020
rect 12012 24108 12516 24164
rect 12572 26852 12740 26908
rect 12796 26908 12852 26918
rect 12012 20244 12068 24108
rect 12124 23940 12180 23950
rect 12124 23938 12292 23940
rect 12124 23886 12126 23938
rect 12178 23886 12292 23938
rect 12124 23884 12292 23886
rect 12124 23874 12180 23884
rect 12124 22932 12180 22942
rect 12124 22148 12180 22876
rect 12236 22370 12292 23884
rect 12236 22318 12238 22370
rect 12290 22318 12292 22370
rect 12236 22306 12292 22318
rect 12460 23154 12516 23166
rect 12460 23102 12462 23154
rect 12514 23102 12516 23154
rect 12460 22260 12516 23102
rect 12572 22820 12628 26852
rect 12796 25506 12852 26852
rect 12908 26068 12964 27692
rect 13020 26628 13076 26638
rect 13020 26290 13076 26572
rect 13020 26238 13022 26290
rect 13074 26238 13076 26290
rect 13020 26226 13076 26238
rect 13132 26292 13188 29036
rect 13132 26226 13188 26236
rect 13244 29036 13412 29092
rect 13468 29260 13580 29316
rect 13468 29092 13524 29260
rect 13580 29222 13636 29260
rect 13244 26404 13300 29036
rect 13468 29026 13524 29036
rect 13916 28980 13972 29484
rect 14028 29428 14084 29438
rect 14028 29334 14084 29372
rect 13804 28924 13972 28980
rect 13692 28644 13748 28654
rect 13804 28644 13860 28924
rect 14140 28756 14196 30158
rect 14364 30324 14420 30334
rect 14364 29650 14420 30268
rect 14588 29764 14644 32396
rect 14700 30884 14756 30894
rect 14700 30790 14756 30828
rect 14588 29698 14644 29708
rect 14700 30100 14756 30110
rect 14364 29598 14366 29650
rect 14418 29598 14420 29650
rect 14364 29586 14420 29598
rect 13692 28642 13860 28644
rect 13692 28590 13694 28642
rect 13746 28590 13860 28642
rect 13692 28588 13860 28590
rect 14028 28700 14196 28756
rect 14252 29426 14308 29438
rect 14252 29374 14254 29426
rect 14306 29374 14308 29426
rect 13692 28578 13748 28588
rect 14028 28532 14084 28700
rect 14252 28644 14308 29374
rect 14476 29426 14532 29438
rect 14476 29374 14478 29426
rect 14530 29374 14532 29426
rect 13244 26290 13300 26348
rect 13244 26238 13246 26290
rect 13298 26238 13300 26290
rect 13244 26226 13300 26238
rect 13356 28420 13412 28430
rect 12908 26012 13076 26068
rect 12908 25620 12964 25630
rect 12908 25526 12964 25564
rect 12796 25454 12798 25506
rect 12850 25454 12852 25506
rect 12796 25442 12852 25454
rect 12908 25172 12964 25182
rect 12684 24722 12740 24734
rect 12684 24670 12686 24722
rect 12738 24670 12740 24722
rect 12684 24500 12740 24670
rect 12684 24434 12740 24444
rect 12572 22754 12628 22764
rect 12684 23940 12740 23950
rect 12572 22372 12628 22382
rect 12684 22372 12740 23884
rect 12572 22370 12740 22372
rect 12572 22318 12574 22370
rect 12626 22318 12740 22370
rect 12572 22316 12740 22318
rect 12796 23938 12852 23950
rect 12796 23886 12798 23938
rect 12850 23886 12852 23938
rect 12572 22306 12628 22316
rect 12124 22092 12292 22148
rect 12124 21700 12180 21710
rect 12124 21476 12180 21644
rect 12124 21382 12180 21420
rect 12236 20914 12292 22092
rect 12460 21812 12516 22204
rect 12796 22036 12852 23886
rect 12908 23826 12964 25116
rect 12908 23774 12910 23826
rect 12962 23774 12964 23826
rect 12908 23762 12964 23774
rect 12460 21746 12516 21756
rect 12572 21980 12852 22036
rect 12908 22820 12964 22830
rect 12572 21588 12628 21980
rect 12908 21924 12964 22764
rect 12684 21812 12740 21822
rect 12908 21812 12964 21868
rect 12684 21810 12964 21812
rect 12684 21758 12686 21810
rect 12738 21758 12964 21810
rect 12684 21756 12964 21758
rect 12684 21746 12740 21756
rect 13020 21588 13076 26012
rect 13356 25172 13412 28364
rect 13580 28418 13636 28430
rect 13580 28366 13582 28418
rect 13634 28366 13636 28418
rect 13580 28196 13636 28366
rect 13580 28130 13636 28140
rect 14028 28418 14084 28476
rect 14028 28366 14030 28418
rect 14082 28366 14084 28418
rect 13692 27972 13748 27982
rect 13692 27878 13748 27916
rect 13468 27858 13524 27870
rect 13468 27806 13470 27858
rect 13522 27806 13524 27858
rect 13468 26404 13524 27806
rect 14028 27748 14084 28366
rect 14140 28588 14308 28644
rect 14364 29092 14420 29102
rect 14140 28196 14196 28588
rect 14140 28130 14196 28140
rect 14252 28420 14308 28430
rect 14028 27682 14084 27692
rect 13580 27412 13636 27422
rect 13580 26516 13636 27356
rect 13804 27188 13860 27198
rect 14028 27188 14084 27198
rect 13580 26450 13636 26460
rect 13692 27186 14028 27188
rect 13692 27134 13806 27186
rect 13858 27134 14028 27186
rect 13692 27132 14028 27134
rect 13468 26338 13524 26348
rect 13580 26290 13636 26302
rect 13580 26238 13582 26290
rect 13634 26238 13636 26290
rect 13580 26180 13636 26238
rect 13580 25732 13636 26124
rect 13580 25666 13636 25676
rect 13468 25284 13524 25294
rect 13468 25190 13524 25228
rect 13356 25106 13412 25116
rect 13468 23828 13524 23838
rect 13244 23604 13300 23614
rect 13244 23154 13300 23548
rect 13244 23102 13246 23154
rect 13298 23102 13300 23154
rect 13244 22932 13300 23102
rect 13244 22866 13300 22876
rect 12572 21522 12628 21532
rect 12684 21586 13076 21588
rect 12684 21534 13022 21586
rect 13074 21534 13076 21586
rect 12684 21532 13076 21534
rect 12236 20862 12238 20914
rect 12290 20862 12292 20914
rect 12236 20850 12292 20862
rect 12684 20914 12740 21532
rect 13020 21522 13076 21532
rect 13244 21924 13300 21934
rect 13244 21586 13300 21868
rect 13244 21534 13246 21586
rect 13298 21534 13300 21586
rect 13244 21522 13300 21534
rect 12684 20862 12686 20914
rect 12738 20862 12740 20914
rect 12012 20188 12180 20244
rect 11676 20078 11678 20130
rect 11730 20078 11732 20130
rect 11676 20066 11732 20078
rect 11788 20130 11956 20132
rect 11788 20078 11902 20130
rect 11954 20078 11956 20130
rect 11788 20076 11956 20078
rect 11564 18510 11566 18562
rect 11618 18510 11620 18562
rect 11564 18498 11620 18510
rect 11564 17442 11620 17454
rect 11564 17390 11566 17442
rect 11618 17390 11620 17442
rect 11564 17108 11620 17390
rect 11564 17014 11620 17052
rect 11676 17108 11732 17118
rect 11788 17108 11844 20076
rect 11900 20066 11956 20076
rect 12012 20018 12068 20030
rect 12012 19966 12014 20018
rect 12066 19966 12068 20018
rect 11900 19234 11956 19246
rect 11900 19182 11902 19234
rect 11954 19182 11956 19234
rect 11900 19012 11956 19182
rect 11900 18946 11956 18956
rect 12012 17892 12068 19966
rect 12012 17826 12068 17836
rect 12012 17668 12068 17678
rect 12124 17668 12180 20188
rect 12460 20132 12516 20142
rect 12460 20038 12516 20076
rect 12348 19460 12404 19470
rect 12348 19346 12404 19404
rect 12348 19294 12350 19346
rect 12402 19294 12404 19346
rect 12348 19282 12404 19294
rect 12348 18788 12404 18798
rect 12348 18450 12404 18732
rect 12348 18398 12350 18450
rect 12402 18398 12404 18450
rect 12348 18386 12404 18398
rect 12068 17612 12180 17668
rect 12348 17666 12404 17678
rect 12348 17614 12350 17666
rect 12402 17614 12404 17666
rect 12012 17574 12068 17612
rect 12348 17108 12404 17614
rect 11676 17106 11844 17108
rect 11676 17054 11678 17106
rect 11730 17054 11844 17106
rect 11676 17052 11844 17054
rect 12124 17052 12404 17108
rect 12572 17442 12628 17454
rect 12572 17390 12574 17442
rect 12626 17390 12628 17442
rect 11676 17042 11732 17052
rect 11452 16930 11508 16940
rect 11788 16884 11844 16894
rect 12124 16884 12180 17052
rect 12572 16996 12628 17390
rect 12572 16930 12628 16940
rect 11788 16882 12180 16884
rect 11788 16830 11790 16882
rect 11842 16830 12180 16882
rect 11788 16828 12180 16830
rect 12236 16882 12292 16894
rect 12236 16830 12238 16882
rect 12290 16830 12292 16882
rect 11788 16436 11844 16828
rect 11676 16380 11844 16436
rect 11676 16212 11732 16380
rect 12236 16324 12292 16830
rect 12460 16884 12516 16894
rect 12460 16324 12516 16828
rect 12684 16660 12740 20862
rect 12796 21252 12852 21262
rect 12796 20242 12852 21196
rect 13468 20692 13524 23772
rect 13580 22484 13636 22522
rect 13580 22418 13636 22428
rect 13580 22258 13636 22270
rect 13580 22206 13582 22258
rect 13634 22206 13636 22258
rect 13580 21700 13636 22206
rect 13580 21634 13636 21644
rect 13580 21362 13636 21374
rect 13580 21310 13582 21362
rect 13634 21310 13636 21362
rect 13580 21028 13636 21310
rect 13580 20962 13636 20972
rect 13468 20626 13524 20636
rect 12796 20190 12798 20242
rect 12850 20190 12852 20242
rect 12796 19124 12852 20190
rect 13356 20018 13412 20030
rect 13356 19966 13358 20018
rect 13410 19966 13412 20018
rect 12908 19236 12964 19246
rect 12908 19142 12964 19180
rect 12796 17554 12852 19068
rect 13356 18788 13412 19966
rect 13580 19346 13636 19358
rect 13580 19294 13582 19346
rect 13634 19294 13636 19346
rect 13580 18788 13636 19294
rect 13692 19236 13748 27132
rect 13804 27122 13860 27132
rect 14028 27122 14084 27132
rect 14252 27074 14308 28364
rect 14364 27748 14420 29036
rect 14476 28644 14532 29374
rect 14588 29426 14644 29438
rect 14588 29374 14590 29426
rect 14642 29374 14644 29426
rect 14588 29316 14644 29374
rect 14588 29250 14644 29260
rect 14700 29092 14756 30044
rect 14924 29652 14980 33628
rect 15036 33346 15092 33740
rect 15036 33294 15038 33346
rect 15090 33294 15092 33346
rect 15036 33282 15092 33294
rect 15036 33124 15092 33134
rect 15036 32564 15092 33068
rect 15148 33012 15204 33852
rect 15596 33684 15652 33964
rect 15708 33926 15764 33964
rect 15596 33628 15764 33684
rect 15596 33460 15652 33470
rect 15596 33366 15652 33404
rect 15260 33236 15316 33246
rect 15260 33142 15316 33180
rect 15484 33124 15540 33134
rect 15484 33030 15540 33068
rect 15596 33122 15652 33134
rect 15596 33070 15598 33122
rect 15650 33070 15652 33122
rect 15148 32956 15316 33012
rect 15036 31332 15092 32508
rect 15148 31668 15204 31678
rect 15148 31574 15204 31612
rect 15036 31266 15092 31276
rect 15148 31108 15204 31118
rect 15148 31014 15204 31052
rect 15148 30548 15204 30558
rect 15036 29652 15092 29662
rect 14924 29650 15092 29652
rect 14924 29598 15038 29650
rect 15090 29598 15092 29650
rect 14924 29596 15092 29598
rect 15148 29652 15204 30492
rect 15260 30210 15316 32956
rect 15596 32900 15652 33070
rect 15484 32844 15652 32900
rect 15372 32788 15428 32798
rect 15372 32562 15428 32732
rect 15372 32510 15374 32562
rect 15426 32510 15428 32562
rect 15372 31948 15428 32510
rect 15484 32452 15540 32844
rect 15484 32386 15540 32396
rect 15596 32674 15652 32686
rect 15596 32622 15598 32674
rect 15650 32622 15652 32674
rect 15596 32004 15652 32622
rect 15372 31892 15540 31948
rect 15596 31938 15652 31948
rect 15372 31778 15428 31790
rect 15372 31726 15374 31778
rect 15426 31726 15428 31778
rect 15372 31668 15428 31726
rect 15372 31602 15428 31612
rect 15260 30158 15262 30210
rect 15314 30158 15316 30210
rect 15260 30146 15316 30158
rect 15372 30212 15428 30222
rect 15484 30212 15540 31892
rect 15708 31780 15764 33628
rect 16268 33572 16324 33582
rect 16044 33346 16100 33358
rect 16044 33294 16046 33346
rect 16098 33294 16100 33346
rect 16044 32228 16100 33294
rect 16268 33346 16324 33516
rect 16268 33294 16270 33346
rect 16322 33294 16324 33346
rect 16268 33282 16324 33294
rect 16380 33348 16436 34300
rect 16492 34132 16548 34142
rect 16492 34038 16548 34076
rect 16492 33348 16548 33358
rect 16380 33346 16548 33348
rect 16380 33294 16494 33346
rect 16546 33294 16548 33346
rect 16380 33292 16548 33294
rect 16380 33124 16436 33134
rect 16380 33030 16436 33068
rect 16492 32900 16548 33292
rect 16268 32844 16548 32900
rect 16268 32564 16324 32844
rect 16492 32676 16548 32686
rect 16268 32508 16436 32564
rect 16268 32340 16324 32350
rect 16268 32246 16324 32284
rect 16044 31892 16100 32172
rect 16044 31826 16100 31836
rect 16268 32004 16324 32014
rect 16268 31890 16324 31948
rect 16268 31838 16270 31890
rect 16322 31838 16324 31890
rect 16268 31826 16324 31838
rect 15708 31778 15988 31780
rect 15708 31726 15710 31778
rect 15762 31726 15988 31778
rect 15708 31724 15988 31726
rect 15708 31714 15764 31724
rect 15596 31668 15652 31678
rect 15596 31218 15652 31612
rect 15932 31332 15988 31724
rect 16044 31666 16100 31678
rect 16044 31614 16046 31666
rect 16098 31614 16100 31666
rect 16044 31556 16100 31614
rect 16044 31490 16100 31500
rect 16380 31668 16436 32508
rect 16492 32340 16548 32620
rect 16604 32564 16660 36540
rect 16716 36530 16772 36540
rect 17276 36484 17332 36494
rect 17276 36482 17444 36484
rect 17276 36430 17278 36482
rect 17330 36430 17444 36482
rect 17276 36428 17444 36430
rect 17276 36418 17332 36428
rect 17388 35698 17444 36428
rect 17388 35646 17390 35698
rect 17442 35646 17444 35698
rect 17388 35588 17444 35646
rect 17388 35522 17444 35532
rect 17500 36258 17556 36270
rect 17500 36206 17502 36258
rect 17554 36206 17556 36258
rect 16940 34914 16996 34926
rect 16940 34862 16942 34914
rect 16994 34862 16996 34914
rect 16828 34242 16884 34254
rect 16828 34190 16830 34242
rect 16882 34190 16884 34242
rect 16716 33348 16772 33358
rect 16828 33348 16884 34190
rect 16716 33346 16884 33348
rect 16716 33294 16718 33346
rect 16770 33294 16884 33346
rect 16716 33292 16884 33294
rect 16716 33282 16772 33292
rect 16828 32788 16884 33292
rect 16828 32674 16884 32732
rect 16828 32622 16830 32674
rect 16882 32622 16884 32674
rect 16828 32610 16884 32622
rect 16604 32508 16772 32564
rect 16604 32340 16660 32350
rect 16492 32338 16660 32340
rect 16492 32286 16606 32338
rect 16658 32286 16660 32338
rect 16492 32284 16660 32286
rect 16604 32274 16660 32284
rect 15932 31276 16100 31332
rect 15596 31166 15598 31218
rect 15650 31166 15652 31218
rect 15596 31154 15652 31166
rect 15932 31108 15988 31118
rect 15820 31106 15988 31108
rect 15820 31054 15934 31106
rect 15986 31054 15988 31106
rect 15820 31052 15988 31054
rect 15596 30212 15652 30222
rect 15484 30210 15652 30212
rect 15484 30158 15598 30210
rect 15650 30158 15652 30210
rect 15484 30156 15652 30158
rect 15260 29652 15316 29662
rect 15148 29650 15316 29652
rect 15148 29598 15262 29650
rect 15314 29598 15316 29650
rect 15148 29596 15316 29598
rect 14924 29540 14980 29596
rect 15036 29586 15092 29596
rect 14924 29474 14980 29484
rect 15148 29428 15204 29438
rect 15148 29334 15204 29372
rect 15260 29204 15316 29596
rect 15260 29138 15316 29148
rect 14700 29026 14756 29036
rect 15372 28756 15428 30156
rect 15596 30146 15652 30156
rect 15596 29426 15652 29438
rect 15596 29374 15598 29426
rect 15650 29374 15652 29426
rect 15596 29316 15652 29374
rect 14588 28644 14644 28654
rect 15260 28644 15316 28654
rect 15372 28644 15428 28700
rect 14476 28642 15092 28644
rect 14476 28590 14590 28642
rect 14642 28590 15092 28642
rect 14476 28588 15092 28590
rect 14588 28578 14644 28588
rect 14924 28420 14980 28430
rect 14700 28418 14980 28420
rect 14700 28366 14926 28418
rect 14978 28366 14980 28418
rect 14700 28364 14980 28366
rect 14364 27682 14420 27692
rect 14588 27746 14644 27758
rect 14588 27694 14590 27746
rect 14642 27694 14644 27746
rect 14252 27022 14254 27074
rect 14306 27022 14308 27074
rect 14252 26516 14308 27022
rect 14476 26852 14532 26862
rect 14252 26290 14308 26460
rect 14252 26238 14254 26290
rect 14306 26238 14308 26290
rect 14252 26226 14308 26238
rect 14364 26796 14476 26852
rect 13916 25620 13972 25630
rect 13804 25618 13972 25620
rect 13804 25566 13918 25618
rect 13970 25566 13972 25618
rect 13804 25564 13972 25566
rect 13804 22484 13860 25564
rect 13916 25554 13972 25564
rect 14028 25508 14084 25518
rect 14028 25396 14084 25452
rect 13804 22370 13860 22428
rect 13804 22318 13806 22370
rect 13858 22318 13860 22370
rect 13804 22306 13860 22318
rect 13916 25340 14084 25396
rect 13916 23154 13972 25340
rect 14364 24834 14420 26796
rect 14476 26786 14532 26796
rect 14476 26068 14532 26078
rect 14476 25618 14532 26012
rect 14476 25566 14478 25618
rect 14530 25566 14532 25618
rect 14476 25554 14532 25566
rect 14588 25172 14644 27694
rect 14364 24782 14366 24834
rect 14418 24782 14420 24834
rect 14364 24770 14420 24782
rect 14476 25116 14644 25172
rect 14252 24724 14308 24734
rect 14028 24612 14084 24622
rect 14028 24518 14084 24556
rect 14140 23940 14196 23950
rect 14140 23604 14196 23884
rect 14140 23538 14196 23548
rect 13916 23102 13918 23154
rect 13970 23102 13972 23154
rect 13916 22148 13972 23102
rect 13804 22092 13972 22148
rect 13804 21364 13860 22092
rect 13804 21298 13860 21308
rect 13916 21924 13972 21934
rect 13804 20802 13860 20814
rect 13804 20750 13806 20802
rect 13858 20750 13860 20802
rect 13804 20356 13860 20750
rect 13804 20290 13860 20300
rect 13916 20018 13972 21868
rect 14028 21700 14084 21710
rect 14028 21252 14084 21644
rect 14028 21186 14084 21196
rect 14140 21588 14196 21598
rect 14140 20468 14196 21532
rect 13916 19966 13918 20018
rect 13970 19966 13972 20018
rect 13916 19954 13972 19966
rect 14028 20412 14196 20468
rect 14028 19796 14084 20412
rect 13692 19170 13748 19180
rect 13916 19740 14084 19796
rect 13916 19122 13972 19740
rect 14028 19572 14084 19582
rect 14028 19236 14084 19516
rect 14028 19142 14084 19180
rect 13916 19070 13918 19122
rect 13970 19070 13972 19122
rect 13916 19058 13972 19070
rect 13356 18732 13636 18788
rect 12796 17502 12798 17554
rect 12850 17502 12852 17554
rect 12796 17490 12852 17502
rect 13020 17668 13076 17678
rect 13020 16882 13076 17612
rect 13356 17332 13412 18732
rect 14028 18452 14084 18462
rect 13580 17780 13636 17818
rect 13580 17714 13636 17724
rect 13468 17668 13524 17678
rect 13468 17574 13524 17612
rect 14028 17666 14084 18396
rect 14028 17614 14030 17666
rect 14082 17614 14084 17666
rect 13692 17444 13748 17454
rect 13692 17442 13972 17444
rect 13692 17390 13694 17442
rect 13746 17390 13972 17442
rect 13692 17388 13972 17390
rect 13692 17378 13748 17388
rect 13356 17266 13412 17276
rect 13020 16830 13022 16882
rect 13074 16830 13076 16882
rect 13020 16818 13076 16830
rect 13468 17108 13524 17118
rect 13468 16882 13524 17052
rect 13468 16830 13470 16882
rect 13522 16830 13524 16882
rect 12684 16604 13076 16660
rect 12460 16268 12628 16324
rect 12236 16258 12292 16268
rect 11340 16098 11508 16100
rect 11340 16046 11342 16098
rect 11394 16046 11508 16098
rect 11340 16044 11508 16046
rect 11340 16034 11396 16044
rect 11228 15428 11284 15438
rect 11228 15334 11284 15372
rect 11116 15092 11396 15148
rect 11228 14644 11284 14654
rect 11340 14644 11396 15092
rect 11452 14980 11508 16044
rect 11676 15874 11732 16156
rect 11788 16100 11844 16110
rect 11788 16006 11844 16044
rect 12236 16098 12292 16110
rect 12236 16046 12238 16098
rect 12290 16046 12292 16098
rect 12236 15988 12292 16046
rect 12460 16100 12516 16110
rect 12460 16006 12516 16044
rect 12236 15922 12292 15932
rect 11676 15822 11678 15874
rect 11730 15822 11732 15874
rect 11676 15540 11732 15822
rect 11900 15876 11956 15886
rect 11900 15782 11956 15820
rect 12572 15876 12628 16268
rect 12572 15810 12628 15820
rect 12796 15874 12852 15886
rect 12796 15822 12798 15874
rect 12850 15822 12852 15874
rect 11676 15474 11732 15484
rect 12572 15316 12628 15326
rect 11676 15204 11732 15242
rect 12572 15222 12628 15260
rect 11676 15138 11732 15148
rect 12796 15092 12852 15822
rect 13020 15540 13076 16604
rect 12908 15428 12964 15438
rect 12908 15334 12964 15372
rect 12796 15026 12852 15036
rect 11452 14924 11844 14980
rect 11228 14642 11396 14644
rect 11228 14590 11230 14642
rect 11282 14590 11396 14642
rect 11228 14588 11396 14590
rect 11676 14754 11732 14766
rect 11676 14702 11678 14754
rect 11730 14702 11732 14754
rect 11676 14642 11732 14702
rect 11676 14590 11678 14642
rect 11730 14590 11732 14642
rect 11228 14578 11284 14588
rect 11676 14578 11732 14590
rect 11788 14308 11844 14924
rect 13020 14642 13076 15484
rect 13244 16324 13300 16334
rect 13244 16100 13300 16268
rect 13468 16210 13524 16830
rect 13916 16882 13972 17388
rect 14028 17108 14084 17614
rect 14140 18450 14196 18462
rect 14140 18398 14142 18450
rect 14194 18398 14196 18450
rect 14140 17780 14196 18398
rect 14140 17444 14196 17724
rect 14140 17378 14196 17388
rect 14252 17220 14308 24668
rect 14476 23156 14532 25116
rect 14476 23090 14532 23100
rect 14588 24948 14644 24958
rect 14364 22484 14420 22494
rect 14420 22428 14532 22484
rect 14364 22418 14420 22428
rect 14364 20916 14420 20926
rect 14364 20690 14420 20860
rect 14364 20638 14366 20690
rect 14418 20638 14420 20690
rect 14364 20626 14420 20638
rect 14028 17042 14084 17052
rect 14140 17164 14308 17220
rect 14364 20130 14420 20142
rect 14364 20078 14366 20130
rect 14418 20078 14420 20130
rect 13916 16830 13918 16882
rect 13970 16830 13972 16882
rect 13468 16158 13470 16210
rect 13522 16158 13524 16210
rect 13468 16146 13524 16158
rect 13580 16660 13636 16670
rect 13244 15538 13300 16044
rect 13244 15486 13246 15538
rect 13298 15486 13300 15538
rect 13244 15474 13300 15486
rect 13468 15316 13524 15326
rect 13580 15316 13636 16604
rect 13916 16548 13972 16830
rect 14140 16660 14196 17164
rect 14364 16996 14420 20078
rect 14476 19684 14532 22428
rect 14588 20018 14644 24892
rect 14700 23940 14756 28364
rect 14924 28354 14980 28364
rect 14924 27972 14980 27982
rect 15036 27972 15092 28588
rect 15260 28642 15428 28644
rect 15260 28590 15262 28642
rect 15314 28590 15428 28642
rect 15260 28588 15428 28590
rect 15484 29314 15652 29316
rect 15484 29262 15598 29314
rect 15650 29262 15652 29314
rect 15484 29260 15652 29262
rect 15260 28578 15316 28588
rect 15484 28532 15540 29260
rect 15596 29250 15652 29260
rect 15708 29204 15764 29214
rect 15708 28868 15764 29148
rect 14924 27970 15092 27972
rect 14924 27918 14926 27970
rect 14978 27918 15092 27970
rect 14924 27916 15092 27918
rect 14924 27906 14980 27916
rect 14812 27858 14868 27870
rect 14812 27806 14814 27858
rect 14866 27806 14868 27858
rect 14812 27188 14868 27806
rect 14812 27074 14868 27132
rect 14812 27022 14814 27074
rect 14866 27022 14868 27074
rect 14812 27010 14868 27022
rect 14924 27748 14980 27758
rect 14924 26908 14980 27692
rect 15036 27188 15092 27916
rect 15036 27122 15092 27132
rect 15372 28476 15540 28532
rect 15596 28812 15764 28868
rect 15148 27076 15204 27114
rect 15148 27010 15204 27020
rect 14924 26852 15092 26908
rect 15148 26852 15204 26862
rect 15036 26796 15148 26852
rect 15148 26786 15204 26796
rect 15372 26628 15428 28476
rect 15484 28308 15540 28318
rect 15484 28082 15540 28252
rect 15484 28030 15486 28082
rect 15538 28030 15540 28082
rect 15484 28018 15540 28030
rect 15484 27636 15540 27646
rect 15484 27300 15540 27580
rect 15484 27234 15540 27244
rect 15596 26908 15652 28812
rect 15708 28532 15764 28542
rect 15708 28438 15764 28476
rect 15820 27970 15876 31052
rect 15932 31042 15988 31052
rect 15932 30212 15988 30222
rect 15932 30118 15988 30156
rect 16044 29876 16100 31276
rect 16380 30660 16436 31612
rect 16604 31778 16660 31790
rect 16604 31726 16606 31778
rect 16658 31726 16660 31778
rect 16492 31554 16548 31566
rect 16492 31502 16494 31554
rect 16546 31502 16548 31554
rect 16492 31162 16548 31502
rect 16604 31332 16660 31726
rect 16716 31668 16772 32508
rect 16940 32116 16996 34862
rect 17500 34356 17556 36206
rect 19836 36092 20100 36102
rect 19628 36036 19684 36046
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 17836 35586 17892 35598
rect 17836 35534 17838 35586
rect 17890 35534 17892 35586
rect 17836 35364 17892 35534
rect 17836 35298 17892 35308
rect 19628 34356 19684 35980
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 17500 34300 18004 34356
rect 19628 34300 20020 34356
rect 17948 34244 18004 34300
rect 18060 34244 18116 34254
rect 17948 34242 18116 34244
rect 17948 34190 18062 34242
rect 18114 34190 18116 34242
rect 17948 34188 18116 34190
rect 17836 34130 17892 34142
rect 17836 34078 17838 34130
rect 17890 34078 17892 34130
rect 17612 33570 17668 33582
rect 17612 33518 17614 33570
rect 17666 33518 17668 33570
rect 17052 33460 17108 33470
rect 17052 33346 17108 33404
rect 17052 33294 17054 33346
rect 17106 33294 17108 33346
rect 17052 33282 17108 33294
rect 17276 33122 17332 33134
rect 17276 33070 17278 33122
rect 17330 33070 17332 33122
rect 17276 32900 17332 33070
rect 17500 33124 17556 33134
rect 17500 33030 17556 33068
rect 17276 32834 17332 32844
rect 17388 32676 17444 32686
rect 17388 32582 17444 32620
rect 16940 32060 17108 32116
rect 16940 31892 16996 31902
rect 16940 31778 16996 31836
rect 16940 31726 16942 31778
rect 16994 31726 16996 31778
rect 16940 31714 16996 31726
rect 16716 31612 16884 31668
rect 16604 31266 16660 31276
rect 16492 31110 16494 31162
rect 16546 31110 16548 31162
rect 16492 31098 16548 31110
rect 16604 31106 16660 31118
rect 16604 31054 16606 31106
rect 16658 31054 16660 31106
rect 16604 30996 16660 31054
rect 16380 30594 16436 30604
rect 16492 30940 16660 30996
rect 16044 29810 16100 29820
rect 16380 30436 16436 30446
rect 16380 29652 16436 30380
rect 16492 30324 16548 30940
rect 16716 30884 16772 30894
rect 16604 30772 16660 30782
rect 16716 30772 16772 30828
rect 16604 30770 16772 30772
rect 16604 30718 16606 30770
rect 16658 30718 16772 30770
rect 16604 30716 16772 30718
rect 16604 30706 16660 30716
rect 16492 30258 16548 30268
rect 16492 29876 16548 29886
rect 16548 29820 16660 29876
rect 16492 29810 16548 29820
rect 16492 29652 16548 29662
rect 16380 29650 16548 29652
rect 16380 29598 16494 29650
rect 16546 29598 16548 29650
rect 16380 29596 16548 29598
rect 15820 27918 15822 27970
rect 15874 27918 15876 27970
rect 15708 27860 15764 27870
rect 15708 27300 15764 27804
rect 15708 27234 15764 27244
rect 15596 26852 15764 26908
rect 15148 26572 15428 26628
rect 15484 26740 15540 26750
rect 14812 25508 14868 25518
rect 14812 25414 14868 25452
rect 15148 24724 15204 26572
rect 15372 26404 15428 26414
rect 15484 26404 15540 26684
rect 15372 26402 15540 26404
rect 15372 26350 15374 26402
rect 15426 26350 15540 26402
rect 15372 26348 15540 26350
rect 15372 25284 15428 26348
rect 15260 25228 15372 25284
rect 15260 24946 15316 25228
rect 15372 25218 15428 25228
rect 15596 26292 15652 26302
rect 15260 24894 15262 24946
rect 15314 24894 15316 24946
rect 15260 24882 15316 24894
rect 15372 24948 15428 24958
rect 15372 24854 15428 24892
rect 15148 24668 15316 24724
rect 14700 23846 14756 23884
rect 14924 24052 14980 24062
rect 14924 23714 14980 23996
rect 14924 23662 14926 23714
rect 14978 23662 14980 23714
rect 14924 23650 14980 23662
rect 15036 23266 15092 23278
rect 15036 23214 15038 23266
rect 15090 23214 15092 23266
rect 14924 23156 14980 23166
rect 14924 22370 14980 23100
rect 14924 22318 14926 22370
rect 14978 22318 14980 22370
rect 14924 22306 14980 22318
rect 14812 22148 14868 22158
rect 15036 22148 15092 23214
rect 14868 22092 15092 22148
rect 14812 22054 14868 22092
rect 14700 21140 14756 21150
rect 14700 20916 14756 21084
rect 14700 20850 14756 20860
rect 15148 20804 15204 20814
rect 15148 20710 15204 20748
rect 14588 19966 14590 20018
rect 14642 19966 14644 20018
rect 14588 19796 14644 19966
rect 14700 20020 14756 20030
rect 14924 20020 14980 20030
rect 14700 20018 14980 20020
rect 14700 19966 14702 20018
rect 14754 19966 14926 20018
rect 14978 19966 14980 20018
rect 14700 19964 14980 19966
rect 14700 19954 14756 19964
rect 14924 19954 14980 19964
rect 15148 20020 15204 20030
rect 15148 19926 15204 19964
rect 14588 19740 14980 19796
rect 14476 19628 14756 19684
rect 14700 19124 14756 19628
rect 14588 19122 14756 19124
rect 14588 19070 14702 19122
rect 14754 19070 14756 19122
rect 14588 19068 14756 19070
rect 14588 18452 14644 19068
rect 14700 19058 14756 19068
rect 14812 19236 14868 19246
rect 14588 18386 14644 18396
rect 14700 18562 14756 18574
rect 14700 18510 14702 18562
rect 14754 18510 14756 18562
rect 14588 17444 14644 17454
rect 14588 17350 14644 17388
rect 14700 17108 14756 18510
rect 14364 16930 14420 16940
rect 14476 17052 14756 17108
rect 14140 16594 14196 16604
rect 14252 16882 14308 16894
rect 14252 16830 14254 16882
rect 14306 16830 14308 16882
rect 13916 16482 13972 16492
rect 14028 16324 14084 16334
rect 14252 16324 14308 16830
rect 14028 16322 14308 16324
rect 14028 16270 14030 16322
rect 14082 16270 14308 16322
rect 14028 16268 14308 16270
rect 13692 16212 13748 16222
rect 13692 16118 13748 16156
rect 13916 15540 13972 15550
rect 13916 15446 13972 15484
rect 13524 15260 13636 15316
rect 13468 15222 13524 15260
rect 14028 14980 14084 16268
rect 14476 15540 14532 17052
rect 14364 15484 14532 15540
rect 14588 16882 14644 16894
rect 14588 16830 14590 16882
rect 14642 16830 14644 16882
rect 14588 16324 14644 16830
rect 14700 16884 14756 16894
rect 14700 16790 14756 16828
rect 14364 15204 14420 15484
rect 14476 15316 14532 15326
rect 14476 15222 14532 15260
rect 14364 15138 14420 15148
rect 14028 14914 14084 14924
rect 14252 14756 14308 14766
rect 13020 14590 13022 14642
rect 13074 14590 13076 14642
rect 13020 14578 13076 14590
rect 14140 14700 14252 14756
rect 13580 14530 13636 14542
rect 13580 14478 13582 14530
rect 13634 14478 13636 14530
rect 12236 14308 12292 14318
rect 11788 14306 12292 14308
rect 11788 14254 12238 14306
rect 12290 14254 12292 14306
rect 11788 14252 12292 14254
rect 12236 14196 12292 14252
rect 12236 14130 12292 14140
rect 11004 13918 11006 13970
rect 11058 13918 11060 13970
rect 11004 13906 11060 13918
rect 12796 13860 12852 13870
rect 12796 13766 12852 13804
rect 13244 13860 13300 13870
rect 13580 13860 13636 14478
rect 14028 14532 14084 14542
rect 14028 14438 14084 14476
rect 14028 13972 14084 13982
rect 14140 13972 14196 14700
rect 14252 14690 14308 14700
rect 14028 13970 14196 13972
rect 14028 13918 14030 13970
rect 14082 13918 14196 13970
rect 14028 13916 14196 13918
rect 14588 13972 14644 16268
rect 14700 15988 14756 15998
rect 14700 15894 14756 15932
rect 14812 15764 14868 19180
rect 14924 17666 14980 19740
rect 15260 19348 15316 24668
rect 15596 24722 15652 26236
rect 15596 24670 15598 24722
rect 15650 24670 15652 24722
rect 15596 24658 15652 24670
rect 15372 23940 15428 23950
rect 15372 23938 15540 23940
rect 15372 23886 15374 23938
rect 15426 23886 15540 23938
rect 15372 23884 15540 23886
rect 15372 23874 15428 23884
rect 15372 22260 15428 22270
rect 15372 21474 15428 22204
rect 15372 21422 15374 21474
rect 15426 21422 15428 21474
rect 15372 21410 15428 21422
rect 15484 19458 15540 23884
rect 15708 22596 15764 26852
rect 15820 24724 15876 27918
rect 15932 29540 15988 29550
rect 15932 26964 15988 29484
rect 16044 29314 16100 29326
rect 16044 29262 16046 29314
rect 16098 29262 16100 29314
rect 16044 29204 16100 29262
rect 16380 29314 16436 29596
rect 16492 29586 16548 29596
rect 16604 29428 16660 29820
rect 16380 29262 16382 29314
rect 16434 29262 16436 29314
rect 16380 29250 16436 29262
rect 16492 29372 16660 29428
rect 16044 29138 16100 29148
rect 16044 28530 16100 28542
rect 16044 28478 16046 28530
rect 16098 28478 16100 28530
rect 16044 27860 16100 28478
rect 16492 28532 16548 29372
rect 16604 29204 16660 29214
rect 16604 28980 16660 29148
rect 16604 28642 16660 28924
rect 16604 28590 16606 28642
rect 16658 28590 16660 28642
rect 16604 28578 16660 28590
rect 16492 28466 16548 28476
rect 16268 28308 16324 28318
rect 16268 28082 16324 28252
rect 16268 28030 16270 28082
rect 16322 28030 16324 28082
rect 16268 28018 16324 28030
rect 16044 27766 16100 27804
rect 16380 27858 16436 27870
rect 16380 27806 16382 27858
rect 16434 27806 16436 27858
rect 16268 27748 16324 27758
rect 16268 27654 16324 27692
rect 15932 26898 15988 26908
rect 16044 27300 16100 27310
rect 15932 25508 15988 25518
rect 15932 25414 15988 25452
rect 16044 24834 16100 27244
rect 16380 25844 16436 27806
rect 16604 27860 16660 27870
rect 16604 27074 16660 27804
rect 16604 27022 16606 27074
rect 16658 27022 16660 27074
rect 16492 26852 16548 26862
rect 16492 26758 16548 26796
rect 16492 26404 16548 26414
rect 16492 26290 16548 26348
rect 16492 26238 16494 26290
rect 16546 26238 16548 26290
rect 16492 26226 16548 26238
rect 16044 24782 16046 24834
rect 16098 24782 16100 24834
rect 16044 24770 16100 24782
rect 16156 25788 16436 25844
rect 15932 24724 15988 24734
rect 15820 24722 15988 24724
rect 15820 24670 15934 24722
rect 15986 24670 15988 24722
rect 15820 24668 15988 24670
rect 15820 24388 15876 24398
rect 15820 23826 15876 24332
rect 15820 23774 15822 23826
rect 15874 23774 15876 23826
rect 15820 23762 15876 23774
rect 15708 22530 15764 22540
rect 15820 22484 15876 22494
rect 15820 22270 15876 22428
rect 15820 22218 15822 22270
rect 15874 22218 15876 22270
rect 15820 22206 15876 22218
rect 15708 21588 15764 21598
rect 15932 21588 15988 24668
rect 16156 23940 16212 25788
rect 16156 23266 16212 23884
rect 16156 23214 16158 23266
rect 16210 23214 16212 23266
rect 16156 23202 16212 23214
rect 16268 24948 16324 24958
rect 15708 21586 15988 21588
rect 15708 21534 15710 21586
rect 15762 21534 15988 21586
rect 15708 21532 15988 21534
rect 16044 22484 16100 22494
rect 15708 20356 15764 21532
rect 15708 20290 15764 20300
rect 15932 21364 15988 21374
rect 15932 20690 15988 21308
rect 15932 20638 15934 20690
rect 15986 20638 15988 20690
rect 15708 19906 15764 19918
rect 15708 19854 15710 19906
rect 15762 19854 15764 19906
rect 15708 19796 15764 19854
rect 15708 19730 15764 19740
rect 15484 19406 15486 19458
rect 15538 19406 15540 19458
rect 15484 19394 15540 19406
rect 15596 19684 15652 19694
rect 15372 19348 15428 19358
rect 15260 19346 15428 19348
rect 15260 19294 15374 19346
rect 15426 19294 15428 19346
rect 15260 19292 15428 19294
rect 15148 18564 15204 18574
rect 14924 17614 14926 17666
rect 14978 17614 14980 17666
rect 14924 17602 14980 17614
rect 15036 18340 15092 18350
rect 15036 17444 15092 18284
rect 15148 18116 15204 18508
rect 15260 18340 15316 19292
rect 15372 19282 15428 19292
rect 15260 18274 15316 18284
rect 15372 19124 15428 19134
rect 15148 18060 15316 18116
rect 15148 17556 15204 17566
rect 15148 17462 15204 17500
rect 14924 16884 14980 16894
rect 15036 16884 15092 17388
rect 14924 16882 15092 16884
rect 14924 16830 14926 16882
rect 14978 16830 15092 16882
rect 14924 16828 15092 16830
rect 15148 16882 15204 16894
rect 15148 16830 15150 16882
rect 15202 16830 15204 16882
rect 14924 16818 14980 16828
rect 15148 16772 15204 16830
rect 15148 16706 15204 16716
rect 15260 16770 15316 18060
rect 15372 17666 15428 19068
rect 15372 17614 15374 17666
rect 15426 17614 15428 17666
rect 15372 17602 15428 17614
rect 15596 18674 15652 19628
rect 15596 18622 15598 18674
rect 15650 18622 15652 18674
rect 15596 17666 15652 18622
rect 15708 19458 15764 19470
rect 15708 19406 15710 19458
rect 15762 19406 15764 19458
rect 15708 18116 15764 19406
rect 15932 19124 15988 20638
rect 16044 19460 16100 22428
rect 16156 22372 16212 22382
rect 16156 22278 16212 22316
rect 16268 22148 16324 24892
rect 16380 23828 16436 23838
rect 16380 22260 16436 23772
rect 16492 23154 16548 23166
rect 16492 23102 16494 23154
rect 16546 23102 16548 23154
rect 16492 22484 16548 23102
rect 16492 22418 16548 22428
rect 16380 22204 16548 22260
rect 16268 22092 16436 22148
rect 16268 21812 16324 21822
rect 16156 20804 16212 20814
rect 16156 20710 16212 20748
rect 16268 20018 16324 21756
rect 16380 21364 16436 22092
rect 16380 21298 16436 21308
rect 16380 20356 16436 20366
rect 16380 20130 16436 20300
rect 16380 20078 16382 20130
rect 16434 20078 16436 20130
rect 16380 20066 16436 20078
rect 16268 19966 16270 20018
rect 16322 19966 16324 20018
rect 16268 19954 16324 19966
rect 16044 19404 16212 19460
rect 15932 19058 15988 19068
rect 15820 18340 15876 18350
rect 15820 18246 15876 18284
rect 16044 18228 16100 18238
rect 16044 18134 16100 18172
rect 15708 18060 15876 18116
rect 15708 17892 15764 17902
rect 15708 17778 15764 17836
rect 15708 17726 15710 17778
rect 15762 17726 15764 17778
rect 15708 17714 15764 17726
rect 15596 17614 15598 17666
rect 15650 17614 15652 17666
rect 15596 17602 15652 17614
rect 15372 17444 15428 17454
rect 15372 17106 15428 17388
rect 15708 17220 15764 17230
rect 15372 17054 15374 17106
rect 15426 17054 15428 17106
rect 15372 17042 15428 17054
rect 15596 17108 15652 17118
rect 15596 17014 15652 17052
rect 15260 16718 15262 16770
rect 15314 16718 15316 16770
rect 15260 16706 15316 16718
rect 15596 16660 15652 16670
rect 15484 16604 15596 16660
rect 15484 16548 15540 16604
rect 15596 16594 15652 16604
rect 15260 16492 15540 16548
rect 15260 16210 15316 16492
rect 15260 16158 15262 16210
rect 15314 16158 15316 16210
rect 15260 16146 15316 16158
rect 15372 16212 15428 16222
rect 14924 16100 14980 16110
rect 14924 16006 14980 16044
rect 14700 15708 14868 15764
rect 15148 15874 15204 15886
rect 15148 15822 15150 15874
rect 15202 15822 15204 15874
rect 14700 14642 14756 15708
rect 15148 15540 15204 15822
rect 15148 15474 15204 15484
rect 15260 15874 15316 15886
rect 15260 15822 15262 15874
rect 15314 15822 15316 15874
rect 14812 15428 14868 15438
rect 14812 15334 14868 15372
rect 15260 14756 15316 15822
rect 15372 15314 15428 16156
rect 15708 16098 15764 17164
rect 15820 17108 15876 18060
rect 16156 17668 16212 19404
rect 16380 19234 16436 19246
rect 16380 19182 16382 19234
rect 16434 19182 16436 19234
rect 16380 18900 16436 19182
rect 16380 18834 16436 18844
rect 16492 18452 16548 22204
rect 16604 22148 16660 27022
rect 16716 27076 16772 27086
rect 16716 26514 16772 27020
rect 16716 26462 16718 26514
rect 16770 26462 16772 26514
rect 16716 26450 16772 26462
rect 16716 23378 16772 23390
rect 16716 23326 16718 23378
rect 16770 23326 16772 23378
rect 16716 22820 16772 23326
rect 16716 22754 16772 22764
rect 16828 22372 16884 31612
rect 17052 30996 17108 32060
rect 17500 31778 17556 31790
rect 17500 31726 17502 31778
rect 17554 31726 17556 31778
rect 17500 31556 17556 31726
rect 17500 31490 17556 31500
rect 17052 30930 17108 30940
rect 17612 30996 17668 33518
rect 17724 33348 17780 33358
rect 17836 33348 17892 34078
rect 17724 33346 17892 33348
rect 17724 33294 17726 33346
rect 17778 33294 17892 33346
rect 17724 33292 17892 33294
rect 17724 33282 17780 33292
rect 17948 33124 18004 34188
rect 18060 34178 18116 34188
rect 19964 34242 20020 34300
rect 19964 34190 19966 34242
rect 20018 34190 20020 34242
rect 18172 34130 18228 34142
rect 18172 34078 18174 34130
rect 18226 34078 18228 34130
rect 18172 34020 18228 34078
rect 18620 34020 18676 34030
rect 18172 34018 18676 34020
rect 18172 33966 18622 34018
rect 18674 33966 18676 34018
rect 18172 33964 18676 33966
rect 18060 33460 18116 33470
rect 18060 33346 18116 33404
rect 18060 33294 18062 33346
rect 18114 33294 18116 33346
rect 18060 33282 18116 33294
rect 17724 33068 18004 33124
rect 17724 31220 17780 33068
rect 17836 32452 17892 32462
rect 18172 32452 18228 33964
rect 18620 33954 18676 33964
rect 19852 33906 19908 33918
rect 19852 33854 19854 33906
rect 19906 33854 19908 33906
rect 19404 33684 19460 33694
rect 18284 33234 18340 33246
rect 18284 33182 18286 33234
rect 18338 33182 18340 33234
rect 18284 32900 18340 33182
rect 18396 33234 18452 33246
rect 18396 33182 18398 33234
rect 18450 33182 18452 33234
rect 18396 33124 18452 33182
rect 19180 33236 19236 33246
rect 19180 33142 19236 33180
rect 18396 33058 18452 33068
rect 18844 33122 18900 33134
rect 18844 33070 18846 33122
rect 18898 33070 18900 33122
rect 18284 32834 18340 32844
rect 18844 32676 18900 33070
rect 18844 32610 18900 32620
rect 19404 32786 19460 33628
rect 19852 33346 19908 33854
rect 19964 33572 20020 34190
rect 21308 34020 21364 34030
rect 19964 33506 20020 33516
rect 20972 33572 21028 33582
rect 19852 33294 19854 33346
rect 19906 33294 19908 33346
rect 19852 33282 19908 33294
rect 20076 33234 20132 33246
rect 20076 33182 20078 33234
rect 20130 33182 20132 33234
rect 19404 32734 19406 32786
rect 19458 32734 19460 32786
rect 17836 32450 18228 32452
rect 17836 32398 17838 32450
rect 17890 32398 18228 32450
rect 17836 32396 18228 32398
rect 18956 32452 19012 32462
rect 17836 31332 17892 32396
rect 18956 32358 19012 32396
rect 19404 32340 19460 32734
rect 19516 33122 19572 33134
rect 20076 33124 20132 33182
rect 19516 33070 19518 33122
rect 19570 33070 19572 33122
rect 19516 32452 19572 33070
rect 19516 32386 19572 32396
rect 19628 33068 20132 33124
rect 20300 33234 20356 33246
rect 20300 33182 20302 33234
rect 20354 33182 20356 33234
rect 19628 32564 19684 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19404 32274 19460 32284
rect 18284 32004 18340 32014
rect 17948 31556 18004 31566
rect 18004 31500 18228 31556
rect 17948 31462 18004 31500
rect 17836 31276 18004 31332
rect 17724 31164 17892 31220
rect 17612 30930 17668 30940
rect 17388 30098 17444 30110
rect 17388 30046 17390 30098
rect 17442 30046 17444 30098
rect 17388 29092 17444 30046
rect 17836 29876 17892 31164
rect 17836 29810 17892 29820
rect 17388 29026 17444 29036
rect 17836 29428 17892 29438
rect 17836 28868 17892 29372
rect 17836 28802 17892 28812
rect 17500 28644 17556 28654
rect 17500 28550 17556 28588
rect 17164 28532 17220 28542
rect 17164 27300 17220 28476
rect 17164 27074 17220 27244
rect 17164 27022 17166 27074
rect 17218 27022 17220 27074
rect 17164 27010 17220 27022
rect 17276 28418 17332 28430
rect 17276 28366 17278 28418
rect 17330 28366 17332 28418
rect 17276 28196 17332 28366
rect 17836 28418 17892 28430
rect 17836 28366 17838 28418
rect 17890 28366 17892 28418
rect 17836 28196 17892 28366
rect 17276 28140 17892 28196
rect 17276 26628 17332 28140
rect 17612 27746 17668 27758
rect 17612 27694 17614 27746
rect 17666 27694 17668 27746
rect 17612 26740 17668 27694
rect 17948 26908 18004 31276
rect 18060 29426 18116 29438
rect 18060 29374 18062 29426
rect 18114 29374 18116 29426
rect 18060 29204 18116 29374
rect 18060 28082 18116 29148
rect 18060 28030 18062 28082
rect 18114 28030 18116 28082
rect 18060 28018 18116 28030
rect 17612 26674 17668 26684
rect 17724 26852 18004 26908
rect 17276 26562 17332 26572
rect 17388 26516 17444 26526
rect 17388 26422 17444 26460
rect 17724 26292 17780 26852
rect 17500 26236 17780 26292
rect 17500 25956 17556 26236
rect 17948 26180 18004 26190
rect 17948 26086 18004 26124
rect 17164 25900 17556 25956
rect 17612 26068 17668 26078
rect 17052 25508 17108 25518
rect 16828 22148 16884 22316
rect 16604 22092 16772 22148
rect 16716 21812 16772 22092
rect 16828 22082 16884 22092
rect 16940 23492 16996 23502
rect 16940 22370 16996 23436
rect 16940 22318 16942 22370
rect 16994 22318 16996 22370
rect 16940 22036 16996 22318
rect 16940 21970 16996 21980
rect 17052 22596 17108 25452
rect 17164 23492 17220 25900
rect 17388 25732 17444 25742
rect 17388 25638 17444 25676
rect 17276 25508 17332 25518
rect 17276 25506 17444 25508
rect 17276 25454 17278 25506
rect 17330 25454 17444 25506
rect 17276 25452 17444 25454
rect 17276 25442 17332 25452
rect 17276 25060 17332 25070
rect 17276 23938 17332 25004
rect 17276 23886 17278 23938
rect 17330 23886 17332 23938
rect 17276 23874 17332 23886
rect 17388 24722 17444 25452
rect 17500 25172 17556 25182
rect 17500 24946 17556 25116
rect 17500 24894 17502 24946
rect 17554 24894 17556 24946
rect 17500 24882 17556 24894
rect 17388 24670 17390 24722
rect 17442 24670 17444 24722
rect 17164 23426 17220 23436
rect 17388 23604 17444 24670
rect 17612 24722 17668 26012
rect 18060 25956 18116 25966
rect 17836 25506 17892 25518
rect 17836 25454 17838 25506
rect 17890 25454 17892 25506
rect 17724 25394 17780 25406
rect 17724 25342 17726 25394
rect 17778 25342 17780 25394
rect 17724 24836 17780 25342
rect 17836 25396 17892 25454
rect 17836 25330 17892 25340
rect 18060 25394 18116 25900
rect 18060 25342 18062 25394
rect 18114 25342 18116 25394
rect 18060 25330 18116 25342
rect 17724 24770 17780 24780
rect 18060 24836 18116 24846
rect 17612 24670 17614 24722
rect 17666 24670 17668 24722
rect 17500 24612 17556 24622
rect 17500 24388 17556 24556
rect 17612 24500 17668 24670
rect 18060 24722 18116 24780
rect 18060 24670 18062 24722
rect 18114 24670 18116 24722
rect 18060 24658 18116 24670
rect 17612 24444 17892 24500
rect 17500 24332 17668 24388
rect 17388 23266 17444 23548
rect 17388 23214 17390 23266
rect 17442 23214 17444 23266
rect 17388 23202 17444 23214
rect 17500 24052 17556 24062
rect 17500 22820 17556 23996
rect 17612 23940 17668 24332
rect 17724 23940 17780 23950
rect 17612 23938 17780 23940
rect 17612 23886 17726 23938
rect 17778 23886 17780 23938
rect 17612 23884 17780 23886
rect 17724 23874 17780 23884
rect 16716 21756 16996 21812
rect 16828 21474 16884 21486
rect 16828 21422 16830 21474
rect 16882 21422 16884 21474
rect 16828 21364 16884 21422
rect 16828 21298 16884 21308
rect 16940 20804 16996 21756
rect 16828 20802 16996 20804
rect 16828 20750 16942 20802
rect 16994 20750 16996 20802
rect 16828 20748 16996 20750
rect 16604 20580 16660 20590
rect 16604 20242 16660 20524
rect 16828 20356 16884 20748
rect 16940 20738 16996 20748
rect 16828 20290 16884 20300
rect 16940 20580 16996 20590
rect 16604 20190 16606 20242
rect 16658 20190 16660 20242
rect 16604 20178 16660 20190
rect 16828 20020 16884 20030
rect 16828 19926 16884 19964
rect 16716 19906 16772 19918
rect 16716 19854 16718 19906
rect 16770 19854 16772 19906
rect 16716 19572 16772 19854
rect 16716 19516 16884 19572
rect 16380 18396 16548 18452
rect 16716 19348 16772 19358
rect 16156 17574 16212 17612
rect 16268 18226 16324 18238
rect 16268 18174 16270 18226
rect 16322 18174 16324 18226
rect 15820 16994 15876 17052
rect 15820 16942 15822 16994
rect 15874 16942 15876 16994
rect 15820 16212 15876 16942
rect 15820 16146 15876 16156
rect 16044 17556 16100 17566
rect 15708 16046 15710 16098
rect 15762 16046 15764 16098
rect 15708 16034 15764 16046
rect 15932 16100 15988 16110
rect 16044 16100 16100 17500
rect 16156 16882 16212 16894
rect 16156 16830 16158 16882
rect 16210 16830 16212 16882
rect 16156 16660 16212 16830
rect 16156 16594 16212 16604
rect 16268 16658 16324 18174
rect 16380 17666 16436 18396
rect 16492 18226 16548 18238
rect 16492 18174 16494 18226
rect 16546 18174 16548 18226
rect 16492 17892 16548 18174
rect 16716 18116 16772 19292
rect 16716 18050 16772 18060
rect 16492 17826 16548 17836
rect 16716 17780 16772 17790
rect 16716 17686 16772 17724
rect 16380 17614 16382 17666
rect 16434 17614 16436 17666
rect 16380 17556 16436 17614
rect 16604 17668 16660 17678
rect 16604 17574 16660 17612
rect 16380 17490 16436 17500
rect 16716 17556 16772 17566
rect 16716 17462 16772 17500
rect 16380 16996 16436 17006
rect 16380 16902 16436 16940
rect 16828 16994 16884 19516
rect 16940 18674 16996 20524
rect 17052 20020 17108 22540
rect 17388 22764 17556 22820
rect 17612 23154 17668 23166
rect 17612 23102 17614 23154
rect 17666 23102 17668 23154
rect 17164 22372 17220 22382
rect 17164 22278 17220 22316
rect 17388 21812 17444 22764
rect 17500 22596 17556 22606
rect 17612 22596 17668 23102
rect 17836 23154 17892 24444
rect 17836 23102 17838 23154
rect 17890 23102 17892 23154
rect 17556 22540 17668 22596
rect 17724 23042 17780 23054
rect 17724 22990 17726 23042
rect 17778 22990 17780 23042
rect 17500 22530 17556 22540
rect 17724 22484 17780 22990
rect 17836 22932 17892 23102
rect 18060 23492 18116 23502
rect 18060 23154 18116 23436
rect 18060 23102 18062 23154
rect 18114 23102 18116 23154
rect 18060 23090 18116 23102
rect 17836 22866 17892 22876
rect 17948 23044 18004 23054
rect 17612 22428 17780 22484
rect 17500 22372 17556 22382
rect 17500 22278 17556 22316
rect 17612 21924 17668 22428
rect 17724 22260 17780 22270
rect 17724 22166 17780 22204
rect 17612 21858 17668 21868
rect 17052 19954 17108 19964
rect 17276 21756 17444 21812
rect 16940 18622 16942 18674
rect 16994 18622 16996 18674
rect 16940 18610 16996 18622
rect 17276 18340 17332 21756
rect 17500 21698 17556 21710
rect 17500 21646 17502 21698
rect 17554 21646 17556 21698
rect 17388 21588 17444 21598
rect 17388 21494 17444 21532
rect 17388 21364 17444 21374
rect 17500 21364 17556 21646
rect 17836 21588 17892 21598
rect 17444 21308 17668 21364
rect 17388 21298 17444 21308
rect 17612 20242 17668 21308
rect 17612 20190 17614 20242
rect 17666 20190 17668 20242
rect 17612 20178 17668 20190
rect 17836 20468 17892 21532
rect 17948 21364 18004 22988
rect 18172 22484 18228 31500
rect 18284 29650 18340 31948
rect 18620 30996 18676 31006
rect 18396 30884 18452 30922
rect 18620 30902 18676 30940
rect 18396 30818 18452 30828
rect 18956 30770 19012 30782
rect 18956 30718 18958 30770
rect 19010 30718 19012 30770
rect 18396 30660 18452 30670
rect 18396 30212 18452 30604
rect 18508 30212 18564 30222
rect 18396 30210 18564 30212
rect 18396 30158 18510 30210
rect 18562 30158 18564 30210
rect 18396 30156 18564 30158
rect 18508 30146 18564 30156
rect 18844 29988 18900 29998
rect 18844 29894 18900 29932
rect 18284 29598 18286 29650
rect 18338 29598 18340 29650
rect 18284 29428 18340 29598
rect 18508 29764 18564 29774
rect 18508 29650 18564 29708
rect 18508 29598 18510 29650
rect 18562 29598 18564 29650
rect 18508 29586 18564 29598
rect 18620 29652 18676 29662
rect 18284 29362 18340 29372
rect 18508 29314 18564 29326
rect 18508 29262 18510 29314
rect 18562 29262 18564 29314
rect 18396 28868 18452 28878
rect 18284 28418 18340 28430
rect 18284 28366 18286 28418
rect 18338 28366 18340 28418
rect 18284 28196 18340 28366
rect 18396 28308 18452 28812
rect 18508 28532 18564 29262
rect 18620 28642 18676 29596
rect 18956 29204 19012 30718
rect 19628 30212 19684 32508
rect 19852 32788 19908 32798
rect 20300 32788 20356 33182
rect 19908 32732 20356 32788
rect 20636 33122 20692 33134
rect 20636 33070 20638 33122
rect 20690 33070 20692 33122
rect 19852 32562 19908 32732
rect 19852 32510 19854 32562
rect 19906 32510 19908 32562
rect 19852 32498 19908 32510
rect 20076 32450 20132 32462
rect 20076 32398 20078 32450
rect 20130 32398 20132 32450
rect 19740 32338 19796 32350
rect 19740 32286 19742 32338
rect 19794 32286 19796 32338
rect 19740 32004 19796 32286
rect 19740 31938 19796 31948
rect 20076 31892 20132 32398
rect 20524 32452 20580 32462
rect 20524 32358 20580 32396
rect 20300 32340 20356 32350
rect 20300 32246 20356 32284
rect 20076 31826 20132 31836
rect 20636 31668 20692 33070
rect 20972 32562 21028 33516
rect 21308 32674 21364 33964
rect 23100 32676 23156 32686
rect 21308 32622 21310 32674
rect 21362 32622 21364 32674
rect 21308 32610 21364 32622
rect 22876 32674 23156 32676
rect 22876 32622 23102 32674
rect 23154 32622 23156 32674
rect 22876 32620 23156 32622
rect 20972 32510 20974 32562
rect 21026 32510 21028 32562
rect 20972 32498 21028 32510
rect 21196 32564 21252 32574
rect 21196 32470 21252 32508
rect 22204 32450 22260 32462
rect 22204 32398 22206 32450
rect 22258 32398 22260 32450
rect 20636 31602 20692 31612
rect 20748 32340 20804 32350
rect 21756 32340 21812 32350
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20524 30882 20580 30894
rect 20524 30830 20526 30882
rect 20578 30830 20580 30882
rect 20524 30772 20580 30830
rect 20524 30706 20580 30716
rect 19852 30212 19908 30222
rect 19628 30210 19908 30212
rect 19628 30158 19854 30210
rect 19906 30158 19908 30210
rect 19628 30156 19908 30158
rect 19404 30098 19460 30110
rect 19404 30046 19406 30098
rect 19458 30046 19460 30098
rect 19404 29876 19460 30046
rect 19852 30100 19908 30156
rect 19852 30034 19908 30044
rect 19404 29810 19460 29820
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20636 29652 20692 29662
rect 19068 29540 19124 29550
rect 19068 29538 19236 29540
rect 19068 29486 19070 29538
rect 19122 29486 19236 29538
rect 19068 29484 19236 29486
rect 19068 29474 19124 29484
rect 18956 29138 19012 29148
rect 18620 28590 18622 28642
rect 18674 28590 18676 28642
rect 18620 28578 18676 28590
rect 18732 28868 18788 28878
rect 18508 28466 18564 28476
rect 18396 28252 18676 28308
rect 18284 26292 18340 28140
rect 18620 28082 18676 28252
rect 18620 28030 18622 28082
rect 18674 28030 18676 28082
rect 18620 28018 18676 28030
rect 18396 27858 18452 27870
rect 18396 27806 18398 27858
rect 18450 27806 18452 27858
rect 18396 27412 18452 27806
rect 18732 27860 18788 28812
rect 18844 28756 18900 28766
rect 18844 28084 18900 28700
rect 19068 28642 19124 28654
rect 19068 28590 19070 28642
rect 19122 28590 19124 28642
rect 19068 28532 19124 28590
rect 19068 28466 19124 28476
rect 18844 28028 19012 28084
rect 18844 27860 18900 27870
rect 18732 27858 18900 27860
rect 18732 27806 18846 27858
rect 18898 27806 18900 27858
rect 18732 27804 18900 27806
rect 18844 27748 18900 27804
rect 18844 27682 18900 27692
rect 18956 27634 19012 28028
rect 19068 27860 19124 27870
rect 19068 27766 19124 27804
rect 18956 27582 18958 27634
rect 19010 27582 19012 27634
rect 18956 27570 19012 27582
rect 18396 27346 18452 27356
rect 18508 27300 18564 27310
rect 18284 26226 18340 26236
rect 18396 27188 18452 27198
rect 18396 26290 18452 27132
rect 18508 27074 18564 27244
rect 18508 27022 18510 27074
rect 18562 27022 18564 27074
rect 18508 27010 18564 27022
rect 19180 27076 19236 29484
rect 19404 29428 19460 29438
rect 19404 29334 19460 29372
rect 19292 28868 19348 28878
rect 19348 28812 19460 28868
rect 19292 28802 19348 28812
rect 19404 28642 19460 28812
rect 19404 28590 19406 28642
rect 19458 28590 19460 28642
rect 19404 28578 19460 28590
rect 20300 28644 20356 28654
rect 19292 28530 19348 28542
rect 19292 28478 19294 28530
rect 19346 28478 19348 28530
rect 19292 28420 19348 28478
rect 20188 28532 20244 28542
rect 19292 28354 19348 28364
rect 19852 28420 19908 28458
rect 20188 28438 20244 28476
rect 20300 28530 20356 28588
rect 20300 28478 20302 28530
rect 20354 28478 20356 28530
rect 20300 28466 20356 28478
rect 20524 28420 20580 28430
rect 19852 28354 19908 28364
rect 20412 28418 20580 28420
rect 20412 28366 20526 28418
rect 20578 28366 20580 28418
rect 20412 28364 20580 28366
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20188 28084 20244 28094
rect 19852 27972 19908 27982
rect 19852 27858 19908 27916
rect 19852 27806 19854 27858
rect 19906 27806 19908 27858
rect 19852 27794 19908 27806
rect 19740 27412 19796 27422
rect 19740 27298 19796 27356
rect 19740 27246 19742 27298
rect 19794 27246 19796 27298
rect 19740 27234 19796 27246
rect 20188 27188 20244 28028
rect 20300 27748 20356 27758
rect 20300 27654 20356 27692
rect 20300 27188 20356 27198
rect 20188 27132 20300 27188
rect 20300 27094 20356 27132
rect 19180 27020 19460 27076
rect 18732 26850 18788 26862
rect 18732 26798 18734 26850
rect 18786 26798 18788 26850
rect 18732 26404 18788 26798
rect 18396 26238 18398 26290
rect 18450 26238 18452 26290
rect 18284 25956 18340 25966
rect 18284 25060 18340 25900
rect 18284 24994 18340 25004
rect 18284 24724 18340 24734
rect 18284 24630 18340 24668
rect 18396 24612 18452 26238
rect 18508 26348 18788 26404
rect 19292 26850 19348 26862
rect 19292 26798 19294 26850
rect 19346 26798 19348 26850
rect 19292 26404 19348 26798
rect 18508 25508 18564 26348
rect 19292 26310 19348 26348
rect 19180 26290 19236 26302
rect 19180 26238 19182 26290
rect 19234 26238 19236 26290
rect 18508 25442 18564 25452
rect 18620 26180 18676 26190
rect 18620 25396 18676 26124
rect 18732 26178 18788 26190
rect 18732 26126 18734 26178
rect 18786 26126 18788 26178
rect 18732 26068 18788 26126
rect 18732 26002 18788 26012
rect 18620 25394 19012 25396
rect 18620 25342 18622 25394
rect 18674 25342 19012 25394
rect 18620 25340 19012 25342
rect 18620 25330 18676 25340
rect 18508 25060 18564 25070
rect 18508 24724 18564 25004
rect 18508 24658 18564 24668
rect 18620 24834 18676 24846
rect 18620 24782 18622 24834
rect 18674 24782 18676 24834
rect 18396 24546 18452 24556
rect 18620 24500 18676 24782
rect 18620 24434 18676 24444
rect 18956 24834 19012 25340
rect 19180 25172 19236 26238
rect 19404 26068 19460 27020
rect 19628 26962 19684 26974
rect 19628 26910 19630 26962
rect 19682 26910 19684 26962
rect 19516 26290 19572 26302
rect 19516 26238 19518 26290
rect 19570 26238 19572 26290
rect 19516 26180 19572 26238
rect 19516 26114 19572 26124
rect 19404 25506 19460 26012
rect 19404 25454 19406 25506
rect 19458 25454 19460 25506
rect 19404 25442 19460 25454
rect 19516 25620 19572 25630
rect 19516 25394 19572 25564
rect 19628 25618 19684 26910
rect 19740 26852 19796 26862
rect 20412 26852 20468 28364
rect 20524 28354 20580 28364
rect 20636 28196 20692 29596
rect 19740 26850 20244 26852
rect 19740 26798 19742 26850
rect 19794 26798 20244 26850
rect 19740 26796 20244 26798
rect 19740 26786 19796 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 25566 19630 25618
rect 19682 25566 19684 25618
rect 19628 25554 19684 25566
rect 19852 26516 19908 26526
rect 19516 25342 19518 25394
rect 19570 25342 19572 25394
rect 19516 25330 19572 25342
rect 19740 25396 19796 25406
rect 19852 25396 19908 26460
rect 20188 26404 20244 26796
rect 20076 26348 20244 26404
rect 19964 26178 20020 26190
rect 19964 26126 19966 26178
rect 20018 26126 20020 26178
rect 19964 25620 20020 26126
rect 19964 25554 20020 25564
rect 19964 25396 20020 25406
rect 19852 25340 19964 25396
rect 20076 25396 20132 26348
rect 20412 26292 20468 26796
rect 20188 26236 20468 26292
rect 20524 28140 20692 28196
rect 20188 26178 20244 26236
rect 20188 26126 20190 26178
rect 20242 26126 20244 26178
rect 20188 26114 20244 26126
rect 20412 26066 20468 26078
rect 20412 26014 20414 26066
rect 20466 26014 20468 26066
rect 20412 25956 20468 26014
rect 20412 25890 20468 25900
rect 20524 25508 20580 28140
rect 20748 28082 20804 32284
rect 21420 32338 21812 32340
rect 21420 32286 21758 32338
rect 21810 32286 21812 32338
rect 21420 32284 21812 32286
rect 21308 31892 21364 31902
rect 21308 31798 21364 31836
rect 21420 31332 21476 32284
rect 21756 32274 21812 32284
rect 21532 31780 21588 31790
rect 21532 31686 21588 31724
rect 21308 31276 21476 31332
rect 21868 31554 21924 31566
rect 21868 31502 21870 31554
rect 21922 31502 21924 31554
rect 20972 31220 21028 31230
rect 20972 31126 21028 31164
rect 21308 31108 21364 31276
rect 21308 31014 21364 31052
rect 21420 31108 21476 31118
rect 21420 31106 21588 31108
rect 21420 31054 21422 31106
rect 21474 31054 21588 31106
rect 21420 31052 21588 31054
rect 21420 31042 21476 31052
rect 21084 30884 21140 30894
rect 20972 29428 21028 29438
rect 20972 29314 21028 29372
rect 20972 29262 20974 29314
rect 21026 29262 21028 29314
rect 20972 29250 21028 29262
rect 21084 29204 21140 30828
rect 21420 30772 21476 30782
rect 21196 30770 21476 30772
rect 21196 30718 21422 30770
rect 21474 30718 21476 30770
rect 21196 30716 21476 30718
rect 21196 29426 21252 30716
rect 21420 30706 21476 30716
rect 21532 30436 21588 31052
rect 21532 30370 21588 30380
rect 21868 29764 21924 31502
rect 21980 31556 22036 31566
rect 22204 31556 22260 32398
rect 22764 32450 22820 32462
rect 22764 32398 22766 32450
rect 22818 32398 22820 32450
rect 22540 31892 22596 31902
rect 22540 31798 22596 31836
rect 22764 31892 22820 32398
rect 22316 31778 22372 31790
rect 22316 31726 22318 31778
rect 22370 31726 22372 31778
rect 22316 31668 22372 31726
rect 22316 31602 22372 31612
rect 22036 31500 22260 31556
rect 22652 31556 22708 31566
rect 21980 30994 22036 31500
rect 22652 31462 22708 31500
rect 21980 30942 21982 30994
rect 22034 30942 22036 30994
rect 21980 30772 22036 30942
rect 22204 31220 22260 31230
rect 22204 30994 22260 31164
rect 22540 31218 22596 31230
rect 22540 31166 22542 31218
rect 22594 31166 22596 31218
rect 22204 30942 22206 30994
rect 22258 30942 22260 30994
rect 22204 30930 22260 30942
rect 22428 31108 22484 31118
rect 21980 30706 22036 30716
rect 22428 30324 22484 31052
rect 22428 30258 22484 30268
rect 21868 29698 21924 29708
rect 21420 29540 21476 29550
rect 21420 29446 21476 29484
rect 21868 29538 21924 29550
rect 21868 29486 21870 29538
rect 21922 29486 21924 29538
rect 21196 29374 21198 29426
rect 21250 29374 21252 29426
rect 21196 29362 21252 29374
rect 21868 29316 21924 29486
rect 22540 29540 22596 31166
rect 22652 31220 22708 31230
rect 22764 31220 22820 31836
rect 22708 31164 22820 31220
rect 22876 31554 22932 32620
rect 23100 32610 23156 32620
rect 23100 31778 23156 31790
rect 23100 31726 23102 31778
rect 23154 31726 23156 31778
rect 23100 31668 23156 31726
rect 22876 31502 22878 31554
rect 22930 31502 22932 31554
rect 22876 31220 22932 31502
rect 22652 31154 22708 31164
rect 22876 31154 22932 31164
rect 22988 31612 23100 31668
rect 22988 30660 23044 31612
rect 23100 31602 23156 31612
rect 23100 31108 23156 31118
rect 23100 30994 23156 31052
rect 23100 30942 23102 30994
rect 23154 30942 23156 30994
rect 23100 30930 23156 30942
rect 22988 30594 23044 30604
rect 22988 30100 23044 30110
rect 22988 30006 23044 30044
rect 23100 29986 23156 29998
rect 23100 29934 23102 29986
rect 23154 29934 23156 29986
rect 23100 29540 23156 29934
rect 22540 29484 23156 29540
rect 21868 29250 21924 29260
rect 21084 29148 21364 29204
rect 21308 28754 21364 29148
rect 21308 28702 21310 28754
rect 21362 28702 21364 28754
rect 21308 28690 21364 28702
rect 21756 28756 21812 28766
rect 21756 28662 21812 28700
rect 21532 28644 21588 28654
rect 20748 28030 20750 28082
rect 20802 28030 20804 28082
rect 20748 27972 20804 28030
rect 20748 27906 20804 27916
rect 21420 28642 21588 28644
rect 21420 28590 21534 28642
rect 21586 28590 21588 28642
rect 21420 28588 21588 28590
rect 21420 27412 21476 28588
rect 21532 28578 21588 28588
rect 21980 28642 22036 28654
rect 21980 28590 21982 28642
rect 22034 28590 22036 28642
rect 21420 27298 21476 27356
rect 21420 27246 21422 27298
rect 21474 27246 21476 27298
rect 21420 27234 21476 27246
rect 21980 27300 22036 28590
rect 22428 28644 22484 28654
rect 22428 28550 22484 28588
rect 22540 27746 22596 27758
rect 22540 27694 22542 27746
rect 22594 27694 22596 27746
rect 22540 27524 22596 27694
rect 22540 27458 22596 27468
rect 21980 27234 22036 27244
rect 22316 27300 22372 27310
rect 22372 27244 22484 27300
rect 22316 27206 22372 27244
rect 20636 27188 20692 27198
rect 20636 26290 20692 27132
rect 22204 27076 22260 27086
rect 21756 27074 22260 27076
rect 21756 27022 22206 27074
rect 22258 27022 22260 27074
rect 21756 27020 22260 27022
rect 21532 26850 21588 26862
rect 21532 26798 21534 26850
rect 21586 26798 21588 26850
rect 21532 26516 21588 26798
rect 21644 26852 21700 26862
rect 21644 26758 21700 26796
rect 21532 26450 21588 26460
rect 21644 26516 21700 26526
rect 21756 26516 21812 27020
rect 22204 27010 22260 27020
rect 22316 26964 22372 26974
rect 22316 26870 22372 26908
rect 21644 26514 21812 26516
rect 21644 26462 21646 26514
rect 21698 26462 21812 26514
rect 21644 26460 21812 26462
rect 21980 26852 22036 26862
rect 21644 26450 21700 26460
rect 21420 26402 21476 26414
rect 21420 26350 21422 26402
rect 21474 26350 21476 26402
rect 20636 26238 20638 26290
rect 20690 26238 20692 26290
rect 20636 26226 20692 26238
rect 21084 26292 21140 26302
rect 21084 26198 21140 26236
rect 21308 26290 21364 26302
rect 21308 26238 21310 26290
rect 21362 26238 21364 26290
rect 21308 25956 21364 26238
rect 21308 25890 21364 25900
rect 20524 25414 20580 25452
rect 20636 25620 20692 25630
rect 21420 25620 21476 26350
rect 21644 25956 21700 25966
rect 20412 25396 20468 25406
rect 20076 25340 20356 25396
rect 19740 25302 19796 25340
rect 19964 25302 20020 25340
rect 19404 25284 19460 25294
rect 19404 25172 19460 25228
rect 19404 25116 19684 25172
rect 19180 25106 19236 25116
rect 19628 24948 19684 25116
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20076 24948 20132 24958
rect 20300 24948 20356 25340
rect 19628 24892 19796 24948
rect 18956 24782 18958 24834
rect 19010 24782 19012 24834
rect 18956 24164 19012 24782
rect 19180 24836 19236 24846
rect 19180 24742 19236 24780
rect 19404 24722 19460 24734
rect 19404 24670 19406 24722
rect 19458 24670 19460 24722
rect 19404 24500 19460 24670
rect 19628 24724 19684 24734
rect 19740 24724 19796 24892
rect 20076 24946 20356 24948
rect 20076 24894 20078 24946
rect 20130 24894 20356 24946
rect 20076 24892 20356 24894
rect 20076 24882 20132 24892
rect 20412 24836 20468 25340
rect 20188 24780 20468 24836
rect 19628 24722 19796 24724
rect 19628 24670 19630 24722
rect 19682 24670 19796 24722
rect 19628 24668 19796 24670
rect 19964 24722 20020 24734
rect 19964 24670 19966 24722
rect 20018 24670 20020 24722
rect 19628 24658 19684 24668
rect 19404 24434 19460 24444
rect 19516 24610 19572 24622
rect 19516 24558 19518 24610
rect 19570 24558 19572 24610
rect 19404 24164 19460 24174
rect 18956 24162 19460 24164
rect 18956 24110 19406 24162
rect 19458 24110 19460 24162
rect 18956 24108 19460 24110
rect 18956 23938 19012 24108
rect 19404 24098 19460 24108
rect 18956 23886 18958 23938
rect 19010 23886 19012 23938
rect 18956 23874 19012 23886
rect 18620 23772 18788 23828
rect 18508 23604 18564 23614
rect 18396 23268 18452 23278
rect 17948 21298 18004 21308
rect 18060 22428 18172 22484
rect 18060 20916 18116 22428
rect 18172 22418 18228 22428
rect 18284 22932 18340 22942
rect 18172 22148 18228 22158
rect 18284 22148 18340 22876
rect 18172 22146 18340 22148
rect 18172 22094 18174 22146
rect 18226 22094 18340 22146
rect 18172 22092 18340 22094
rect 18172 22082 18228 22092
rect 17724 20020 17780 20030
rect 17724 19926 17780 19964
rect 17836 19234 17892 20412
rect 17836 19182 17838 19234
rect 17890 19182 17892 19234
rect 17836 19170 17892 19182
rect 17948 20914 18116 20916
rect 17948 20862 18062 20914
rect 18114 20862 18116 20914
rect 17948 20860 18116 20862
rect 17948 18676 18004 20860
rect 18060 20850 18116 20860
rect 18172 20018 18228 20030
rect 18172 19966 18174 20018
rect 18226 19966 18228 20018
rect 18172 19908 18228 19966
rect 17836 18620 18004 18676
rect 18060 19852 18172 19908
rect 17276 17780 17332 18284
rect 17724 18564 17780 18574
rect 17388 17780 17444 17790
rect 17276 17778 17444 17780
rect 17276 17726 17390 17778
rect 17442 17726 17444 17778
rect 17276 17724 17444 17726
rect 17388 17714 17444 17724
rect 17500 17668 17556 17678
rect 17500 17106 17556 17612
rect 17500 17054 17502 17106
rect 17554 17054 17556 17106
rect 17500 17042 17556 17054
rect 17612 17108 17668 17118
rect 17612 17014 17668 17052
rect 17724 17106 17780 18508
rect 17836 17780 17892 18620
rect 17948 18452 18004 18462
rect 17948 18358 18004 18396
rect 18060 18340 18116 19852
rect 18172 19842 18228 19852
rect 18284 19124 18340 22092
rect 18396 20018 18452 23212
rect 18508 22820 18564 23548
rect 18620 23266 18676 23772
rect 18732 23716 18788 23772
rect 18732 23650 18788 23660
rect 18956 23604 19012 23614
rect 19180 23604 19236 23614
rect 19516 23604 19572 24558
rect 19964 24612 20020 24670
rect 20188 24722 20244 24780
rect 20524 24724 20580 24734
rect 20188 24670 20190 24722
rect 20242 24670 20244 24722
rect 20188 24658 20244 24670
rect 20412 24722 20580 24724
rect 20412 24670 20526 24722
rect 20578 24670 20580 24722
rect 20412 24668 20580 24670
rect 19964 24546 20020 24556
rect 20412 24500 20468 24668
rect 20524 24658 20580 24668
rect 20412 24434 20468 24444
rect 19852 24050 19908 24062
rect 19852 23998 19854 24050
rect 19906 23998 19908 24050
rect 19740 23940 19796 23950
rect 19628 23938 19796 23940
rect 19628 23886 19742 23938
rect 19794 23886 19796 23938
rect 19628 23884 19796 23886
rect 19628 23828 19684 23884
rect 19740 23874 19796 23884
rect 19852 23938 19908 23998
rect 19852 23886 19854 23938
rect 19906 23886 19908 23938
rect 19852 23874 19908 23886
rect 20300 23940 20356 23950
rect 20300 23846 20356 23884
rect 20524 23940 20580 23950
rect 20636 23940 20692 25564
rect 21308 25564 21588 25620
rect 20972 25508 21028 25518
rect 21028 25452 21140 25508
rect 20972 25442 21028 25452
rect 20748 25284 20804 25294
rect 20748 25190 20804 25228
rect 20524 23938 20692 23940
rect 20524 23886 20526 23938
rect 20578 23886 20692 23938
rect 20524 23884 20692 23886
rect 20524 23874 20580 23884
rect 19628 23762 19684 23772
rect 20412 23716 20468 23726
rect 20412 23622 20468 23660
rect 19516 23548 19684 23604
rect 18956 23492 19124 23548
rect 19068 23380 19124 23492
rect 19068 23314 19124 23324
rect 18620 23214 18622 23266
rect 18674 23214 18676 23266
rect 18620 23202 18676 23214
rect 18732 23266 18788 23278
rect 18732 23214 18734 23266
rect 18786 23214 18788 23266
rect 18732 23044 18788 23214
rect 18732 22978 18788 22988
rect 18956 23154 19012 23166
rect 18956 23102 18958 23154
rect 19010 23102 19012 23154
rect 18956 22932 19012 23102
rect 18956 22866 19012 22876
rect 18508 22764 18900 22820
rect 18732 22596 18788 22606
rect 18508 22484 18564 22494
rect 18508 22390 18564 22428
rect 18732 22482 18788 22540
rect 18732 22430 18734 22482
rect 18786 22430 18788 22482
rect 18732 22418 18788 22430
rect 18844 22370 18900 22764
rect 18844 22318 18846 22370
rect 18898 22318 18900 22370
rect 18508 22148 18564 22158
rect 18508 21026 18564 22092
rect 18844 21812 18900 22318
rect 19180 22370 19236 23548
rect 19516 23268 19572 23278
rect 19516 23154 19572 23212
rect 19516 23102 19518 23154
rect 19570 23102 19572 23154
rect 19516 23090 19572 23102
rect 19404 23044 19460 23054
rect 19180 22318 19182 22370
rect 19234 22318 19236 22370
rect 19180 22306 19236 22318
rect 19292 22370 19348 22382
rect 19292 22318 19294 22370
rect 19346 22318 19348 22370
rect 19292 22148 19348 22318
rect 19292 22082 19348 22092
rect 19404 21812 19460 22988
rect 19628 22932 19684 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 18844 21746 18900 21756
rect 19292 21756 19460 21812
rect 19516 22876 19684 22932
rect 18956 21700 19012 21710
rect 18508 20974 18510 21026
rect 18562 20974 18564 21026
rect 18508 20914 18564 20974
rect 18508 20862 18510 20914
rect 18562 20862 18564 20914
rect 18508 20850 18564 20862
rect 18844 21026 18900 21038
rect 18844 20974 18846 21026
rect 18898 20974 18900 21026
rect 18396 19966 18398 20018
rect 18450 19966 18452 20018
rect 18396 19954 18452 19966
rect 18844 20580 18900 20974
rect 18956 20804 19012 21644
rect 19292 21028 19348 21756
rect 19404 21588 19460 21598
rect 19404 21494 19460 21532
rect 19404 21028 19460 21038
rect 19292 21026 19460 21028
rect 19292 20974 19406 21026
rect 19458 20974 19460 21026
rect 19292 20972 19460 20974
rect 19404 20962 19460 20972
rect 19292 20804 19348 20814
rect 18956 20748 19124 20804
rect 18956 20580 19012 20590
rect 18844 20578 19012 20580
rect 18844 20526 18958 20578
rect 19010 20526 19012 20578
rect 18844 20524 19012 20526
rect 18732 19906 18788 19918
rect 18732 19854 18734 19906
rect 18786 19854 18788 19906
rect 18508 19348 18564 19358
rect 18284 19058 18340 19068
rect 18396 19236 18452 19246
rect 18284 18676 18340 18686
rect 18396 18676 18452 19180
rect 18340 18620 18452 18676
rect 18508 19234 18564 19292
rect 18508 19182 18510 19234
rect 18562 19182 18564 19234
rect 18284 18582 18340 18620
rect 18172 18564 18228 18574
rect 18172 18470 18228 18508
rect 18508 18564 18564 19182
rect 18508 18498 18564 18508
rect 18396 18340 18452 18350
rect 18060 18284 18340 18340
rect 18284 18226 18340 18284
rect 18284 18174 18286 18226
rect 18338 18174 18340 18226
rect 18284 18162 18340 18174
rect 18396 18004 18452 18284
rect 17836 17724 18340 17780
rect 18060 17444 18116 17454
rect 18060 17350 18116 17388
rect 17724 17054 17726 17106
rect 17778 17054 17780 17106
rect 17724 17042 17780 17054
rect 17948 17332 18004 17342
rect 16828 16942 16830 16994
rect 16882 16942 16884 16994
rect 16828 16930 16884 16942
rect 16604 16884 16660 16894
rect 16604 16790 16660 16828
rect 17836 16884 17892 16894
rect 17836 16790 17892 16828
rect 17948 16882 18004 17276
rect 17948 16830 17950 16882
rect 18002 16830 18004 16882
rect 17948 16818 18004 16830
rect 18060 17108 18116 17118
rect 16268 16606 16270 16658
rect 16322 16606 16324 16658
rect 16268 16594 16324 16606
rect 16380 16772 16436 16782
rect 15932 16098 16100 16100
rect 15932 16046 15934 16098
rect 15986 16046 16100 16098
rect 15932 16044 16100 16046
rect 16380 16100 16436 16716
rect 17612 16324 17668 16334
rect 15932 15988 15988 16044
rect 16380 16006 16436 16044
rect 17052 16098 17108 16110
rect 17052 16046 17054 16098
rect 17106 16046 17108 16098
rect 15932 15922 15988 15932
rect 16156 15988 16212 15998
rect 16156 15894 16212 15932
rect 15372 15262 15374 15314
rect 15426 15262 15428 15314
rect 15372 15250 15428 15262
rect 15820 15876 15876 15886
rect 15820 15540 15876 15820
rect 16044 15876 16100 15886
rect 16044 15782 16100 15820
rect 17052 15764 17108 16046
rect 17500 16100 17556 16110
rect 16380 15652 16436 15662
rect 16044 15540 16100 15550
rect 15820 15538 16100 15540
rect 15820 15486 16046 15538
rect 16098 15486 16100 15538
rect 15820 15484 16100 15486
rect 15372 14756 15428 14766
rect 15260 14700 15372 14756
rect 15372 14690 15428 14700
rect 14700 14590 14702 14642
rect 14754 14590 14756 14642
rect 14700 14578 14756 14590
rect 15372 14532 15428 14542
rect 15148 14476 15372 14532
rect 14812 13972 14868 13982
rect 14588 13970 14868 13972
rect 14588 13918 14814 13970
rect 14866 13918 14868 13970
rect 14588 13916 14868 13918
rect 14028 13906 14084 13916
rect 14812 13906 14868 13916
rect 15148 13970 15204 14476
rect 15372 14438 15428 14476
rect 15148 13918 15150 13970
rect 15202 13918 15204 13970
rect 15148 13906 15204 13918
rect 15708 13972 15764 13982
rect 15820 13972 15876 15484
rect 16044 15474 16100 15484
rect 16380 15538 16436 15596
rect 16380 15486 16382 15538
rect 16434 15486 16436 15538
rect 16380 15428 16436 15486
rect 15932 15314 15988 15326
rect 15932 15262 15934 15314
rect 15986 15262 15988 15314
rect 15932 14644 15988 15262
rect 16156 15316 16212 15326
rect 16156 15222 16212 15260
rect 16268 15314 16324 15326
rect 16268 15262 16270 15314
rect 16322 15262 16324 15314
rect 16268 14756 16324 15262
rect 16268 14690 16324 14700
rect 16156 14644 16212 14654
rect 15932 14588 16156 14644
rect 16380 14644 16436 15372
rect 17052 15148 17108 15708
rect 17164 15876 17220 15886
rect 17164 15316 17220 15820
rect 17276 15874 17332 15886
rect 17276 15822 17278 15874
rect 17330 15822 17332 15874
rect 17276 15540 17332 15822
rect 17388 15874 17444 15886
rect 17388 15822 17390 15874
rect 17442 15822 17444 15874
rect 17388 15652 17444 15822
rect 17500 15764 17556 16044
rect 17612 16098 17668 16268
rect 17612 16046 17614 16098
rect 17666 16046 17668 16098
rect 17612 16034 17668 16046
rect 18060 16098 18116 17052
rect 18060 16046 18062 16098
rect 18114 16046 18116 16098
rect 18060 16034 18116 16046
rect 18172 16884 18228 16894
rect 17500 15708 17668 15764
rect 17388 15596 17556 15652
rect 17276 15474 17332 15484
rect 17388 15426 17444 15438
rect 17388 15374 17390 15426
rect 17442 15374 17444 15426
rect 17388 15316 17444 15374
rect 17164 15260 17444 15316
rect 17500 15314 17556 15596
rect 17500 15262 17502 15314
rect 17554 15262 17556 15314
rect 17500 15250 17556 15262
rect 17052 15092 17220 15148
rect 16492 14644 16548 14654
rect 16380 14642 16548 14644
rect 16380 14590 16494 14642
rect 16546 14590 16548 14642
rect 16380 14588 16548 14590
rect 16156 14550 16212 14588
rect 16492 14578 16548 14588
rect 16940 14530 16996 14542
rect 16940 14478 16942 14530
rect 16994 14478 16996 14530
rect 15708 13970 15876 13972
rect 15708 13918 15710 13970
rect 15762 13918 15876 13970
rect 15708 13916 15876 13918
rect 16268 13972 16324 13982
rect 15708 13906 15764 13916
rect 16268 13878 16324 13916
rect 16940 13972 16996 14478
rect 17164 14420 17220 15092
rect 17612 14532 17668 15708
rect 18172 15314 18228 16828
rect 18172 15262 18174 15314
rect 18226 15262 18228 15314
rect 18172 14642 18228 15262
rect 18284 15986 18340 17724
rect 18396 16996 18452 17948
rect 18620 17892 18676 17902
rect 18620 17778 18676 17836
rect 18620 17726 18622 17778
rect 18674 17726 18676 17778
rect 18620 17714 18676 17726
rect 18508 17556 18564 17566
rect 18508 17220 18564 17500
rect 18508 17164 18676 17220
rect 18508 16996 18564 17006
rect 18396 16994 18564 16996
rect 18396 16942 18510 16994
rect 18562 16942 18564 16994
rect 18396 16940 18564 16942
rect 18284 15934 18286 15986
rect 18338 15934 18340 15986
rect 18284 15148 18340 15934
rect 18508 15988 18564 16940
rect 18620 16210 18676 17164
rect 18620 16158 18622 16210
rect 18674 16158 18676 16210
rect 18620 16146 18676 16158
rect 18508 15922 18564 15932
rect 18732 15538 18788 19854
rect 18844 19348 18900 20524
rect 18956 20514 19012 20524
rect 19068 19796 19124 20748
rect 19292 20710 19348 20748
rect 19404 20578 19460 20590
rect 19404 20526 19406 20578
rect 19458 20526 19460 20578
rect 19404 20468 19460 20526
rect 19404 20402 19460 20412
rect 19404 20020 19460 20030
rect 19068 19740 19348 19796
rect 18844 18452 18900 19292
rect 19180 19124 19236 19134
rect 19180 19030 19236 19068
rect 18844 18228 18900 18396
rect 18844 18162 18900 18172
rect 19180 18452 19236 18462
rect 19180 18116 19236 18396
rect 18956 18004 19012 18014
rect 18956 17890 19012 17948
rect 18956 17838 18958 17890
rect 19010 17838 19012 17890
rect 18956 17826 19012 17838
rect 18844 17668 18900 17678
rect 18844 17574 18900 17612
rect 18956 17444 19012 17454
rect 18956 17350 19012 17388
rect 18844 17332 18900 17342
rect 18844 17108 18900 17276
rect 19180 17108 19236 18060
rect 19292 17892 19348 19740
rect 19404 19346 19460 19964
rect 19404 19294 19406 19346
rect 19458 19294 19460 19346
rect 19404 19282 19460 19294
rect 19516 18564 19572 22876
rect 20636 22708 20692 23884
rect 20860 24834 20916 24846
rect 20860 24782 20862 24834
rect 20914 24782 20916 24834
rect 20860 23380 20916 24782
rect 21084 24722 21140 25452
rect 21308 25284 21364 25564
rect 21308 25218 21364 25228
rect 21420 25396 21476 25406
rect 21084 24670 21086 24722
rect 21138 24670 21140 24722
rect 21084 24658 21140 24670
rect 21420 24162 21476 25340
rect 21420 24110 21422 24162
rect 21474 24110 21476 24162
rect 21420 24098 21476 24110
rect 21308 23938 21364 23950
rect 21308 23886 21310 23938
rect 21362 23886 21364 23938
rect 21196 23828 21252 23838
rect 21308 23828 21364 23886
rect 21252 23772 21364 23828
rect 21532 23828 21588 25564
rect 21644 24948 21700 25900
rect 21644 24946 21924 24948
rect 21644 24894 21646 24946
rect 21698 24894 21924 24946
rect 21644 24892 21924 24894
rect 21644 24882 21700 24892
rect 21868 24052 21924 24892
rect 21532 23772 21700 23828
rect 21196 23762 21252 23772
rect 21420 23716 21476 23726
rect 21420 23548 21476 23660
rect 21420 23492 21588 23548
rect 20860 23324 21140 23380
rect 20860 23156 20916 23324
rect 20860 23090 20916 23100
rect 20972 23154 21028 23166
rect 20972 23102 20974 23154
rect 21026 23102 21028 23154
rect 20636 22652 20916 22708
rect 20076 22596 20132 22606
rect 20132 22540 20244 22596
rect 20076 22530 20132 22540
rect 19628 22484 19684 22494
rect 19628 22370 19684 22428
rect 19628 22318 19630 22370
rect 19682 22318 19684 22370
rect 19628 22306 19684 22318
rect 19852 22370 19908 22382
rect 19852 22318 19854 22370
rect 19906 22318 19908 22370
rect 19852 22148 19908 22318
rect 19852 22082 19908 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21028 20244 22540
rect 20636 22484 20692 22494
rect 20636 22390 20692 22428
rect 20748 22260 20804 22270
rect 20636 22258 20804 22260
rect 20636 22206 20750 22258
rect 20802 22206 20804 22258
rect 20636 22204 20804 22206
rect 20300 22148 20356 22158
rect 20300 22146 20468 22148
rect 20300 22094 20302 22146
rect 20354 22094 20468 22146
rect 20300 22092 20468 22094
rect 20300 22082 20356 22092
rect 20412 21140 20468 22092
rect 20300 21028 20356 21038
rect 20188 21026 20356 21028
rect 20188 20974 20302 21026
rect 20354 20974 20356 21026
rect 20188 20972 20356 20974
rect 20300 20962 20356 20972
rect 20076 20804 20132 20814
rect 20076 20802 20244 20804
rect 20076 20750 20078 20802
rect 20130 20750 20244 20802
rect 20076 20748 20244 20750
rect 20076 20738 20132 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20132 20244 20748
rect 20300 20244 20356 20254
rect 20412 20244 20468 21084
rect 20524 22146 20580 22158
rect 20524 22094 20526 22146
rect 20578 22094 20580 22146
rect 20524 20916 20580 22094
rect 20636 21028 20692 22204
rect 20748 22194 20804 22204
rect 20748 22036 20804 22046
rect 20748 21252 20804 21980
rect 20860 21924 20916 22652
rect 20860 21858 20916 21868
rect 20860 21700 20916 21710
rect 20860 21586 20916 21644
rect 20860 21534 20862 21586
rect 20914 21534 20916 21586
rect 20860 21522 20916 21534
rect 20748 21196 20916 21252
rect 20748 21028 20804 21038
rect 20636 21026 20748 21028
rect 20636 20974 20638 21026
rect 20690 20974 20748 21026
rect 20636 20972 20748 20974
rect 20636 20962 20692 20972
rect 20748 20962 20804 20972
rect 20524 20850 20580 20860
rect 20860 20804 20916 21196
rect 20300 20242 20468 20244
rect 20300 20190 20302 20242
rect 20354 20190 20468 20242
rect 20300 20188 20468 20190
rect 20636 20748 20916 20804
rect 20300 20178 20356 20188
rect 20076 20076 20244 20132
rect 20076 19684 20132 20076
rect 20188 19908 20244 19918
rect 20188 19814 20244 19852
rect 20076 19628 20244 19684
rect 19964 19572 20020 19582
rect 20020 19516 20132 19572
rect 19964 19506 20020 19516
rect 20076 19234 20132 19516
rect 20188 19346 20244 19628
rect 20188 19294 20190 19346
rect 20242 19294 20244 19346
rect 20188 19282 20244 19294
rect 20636 19236 20692 20748
rect 20972 20692 21028 23102
rect 21084 22036 21140 23324
rect 21084 21970 21140 21980
rect 21308 21810 21364 21822
rect 21308 21758 21310 21810
rect 21362 21758 21364 21810
rect 21308 21700 21364 21758
rect 21308 21634 21364 21644
rect 21420 21812 21476 21822
rect 21420 21698 21476 21756
rect 21420 21646 21422 21698
rect 21474 21646 21476 21698
rect 21308 21252 21364 21262
rect 21420 21252 21476 21646
rect 21364 21196 21476 21252
rect 21308 21186 21364 21196
rect 21084 21140 21140 21150
rect 21140 21084 21252 21140
rect 21084 21074 21140 21084
rect 21196 20916 21252 21084
rect 21308 20916 21364 20926
rect 21196 20914 21364 20916
rect 21196 20862 21310 20914
rect 21362 20862 21364 20914
rect 21196 20860 21364 20862
rect 21308 20850 21364 20860
rect 21420 20916 21476 20926
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 20076 19170 20132 19182
rect 20412 19234 20692 19236
rect 20412 19182 20638 19234
rect 20690 19182 20692 19234
rect 20412 19180 20692 19182
rect 19628 19012 19684 19022
rect 19628 18676 19684 18956
rect 20300 19012 20356 19022
rect 20300 18918 20356 18956
rect 20188 18900 20244 18910
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19852 18676 19908 18686
rect 19628 18674 19908 18676
rect 19628 18622 19854 18674
rect 19906 18622 19908 18674
rect 19628 18620 19908 18622
rect 19852 18610 19908 18620
rect 19964 18676 20020 18686
rect 19516 18508 19796 18564
rect 19404 18450 19460 18462
rect 19404 18398 19406 18450
rect 19458 18398 19460 18450
rect 19404 18228 19460 18398
rect 19404 18162 19460 18172
rect 19628 18004 19684 18014
rect 19292 17836 19572 17892
rect 19404 17668 19460 17678
rect 18844 17106 19012 17108
rect 18844 17054 18846 17106
rect 18898 17054 19012 17106
rect 18844 17052 19012 17054
rect 18844 17042 18900 17052
rect 18732 15486 18734 15538
rect 18786 15486 18788 15538
rect 18732 15474 18788 15486
rect 18844 16212 18900 16222
rect 18620 15316 18676 15326
rect 18620 15222 18676 15260
rect 18844 15148 18900 16156
rect 18956 15876 19012 17052
rect 19180 17042 19236 17052
rect 19292 17666 19460 17668
rect 19292 17614 19406 17666
rect 19458 17614 19460 17666
rect 19292 17612 19460 17614
rect 19180 16882 19236 16894
rect 19180 16830 19182 16882
rect 19234 16830 19236 16882
rect 19068 16324 19124 16334
rect 19180 16324 19236 16830
rect 19124 16268 19236 16324
rect 19068 16098 19124 16268
rect 19292 16212 19348 17612
rect 19404 17602 19460 17612
rect 19404 17108 19460 17118
rect 19516 17108 19572 17836
rect 19628 17554 19684 17948
rect 19628 17502 19630 17554
rect 19682 17502 19684 17554
rect 19628 17490 19684 17502
rect 19740 17444 19796 18508
rect 19964 18450 20020 18620
rect 19964 18398 19966 18450
rect 20018 18398 20020 18450
rect 19964 18386 20020 18398
rect 20076 18450 20132 18462
rect 20076 18398 20078 18450
rect 20130 18398 20132 18450
rect 20076 18004 20132 18398
rect 20076 17938 20132 17948
rect 20076 17556 20132 17566
rect 20076 17462 20132 17500
rect 19740 17378 19796 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19404 17106 19572 17108
rect 19404 17054 19406 17106
rect 19458 17054 19572 17106
rect 19404 17052 19572 17054
rect 19628 17108 19684 17118
rect 20188 17108 20244 18844
rect 20412 18674 20468 19180
rect 20636 19170 20692 19180
rect 20748 20636 21028 20692
rect 21420 20690 21476 20860
rect 21420 20638 21422 20690
rect 21474 20638 21476 20690
rect 20412 18622 20414 18674
rect 20466 18622 20468 18674
rect 19404 17042 19460 17052
rect 19628 17014 19684 17052
rect 20076 17052 20244 17108
rect 20300 18228 20356 18238
rect 19852 16996 19908 17006
rect 19852 16882 19908 16940
rect 19852 16830 19854 16882
rect 19906 16830 19908 16882
rect 19852 16818 19908 16830
rect 19516 16772 19572 16782
rect 19516 16678 19572 16716
rect 19404 16212 19460 16222
rect 19292 16210 19460 16212
rect 19292 16158 19406 16210
rect 19458 16158 19460 16210
rect 19292 16156 19460 16158
rect 19404 16146 19460 16156
rect 19068 16046 19070 16098
rect 19122 16046 19124 16098
rect 19068 16034 19124 16046
rect 19740 16100 19796 16110
rect 19740 16006 19796 16044
rect 19404 15988 19460 15998
rect 19292 15876 19348 15886
rect 18956 15874 19348 15876
rect 18956 15822 19294 15874
rect 19346 15822 19348 15874
rect 18956 15820 19348 15822
rect 19292 15810 19348 15820
rect 19404 15538 19460 15932
rect 19404 15486 19406 15538
rect 19458 15486 19460 15538
rect 19404 15474 19460 15486
rect 19516 15874 19572 15886
rect 19516 15822 19518 15874
rect 19570 15822 19572 15874
rect 19516 15540 19572 15822
rect 19516 15474 19572 15484
rect 19628 15876 19684 15886
rect 20076 15876 20132 17052
rect 20188 16772 20244 16782
rect 20188 16678 20244 16716
rect 20188 15876 20244 15886
rect 20076 15874 20244 15876
rect 20076 15822 20190 15874
rect 20242 15822 20244 15874
rect 20076 15820 20244 15822
rect 19628 15428 19684 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19740 15428 19796 15438
rect 19628 15426 19796 15428
rect 19628 15374 19742 15426
rect 19794 15374 19796 15426
rect 19628 15372 19796 15374
rect 19740 15204 19796 15372
rect 18284 15092 18564 15148
rect 18844 15092 19012 15148
rect 19740 15138 19796 15148
rect 18172 14590 18174 14642
rect 18226 14590 18228 14642
rect 18172 14578 18228 14590
rect 18508 14644 18564 15092
rect 17612 14530 18116 14532
rect 17612 14478 17614 14530
rect 17666 14478 18116 14530
rect 17612 14476 18116 14478
rect 17612 14466 17668 14476
rect 17500 14420 17556 14430
rect 17164 14418 17556 14420
rect 17164 14366 17502 14418
rect 17554 14366 17556 14418
rect 17164 14364 17556 14366
rect 17500 14354 17556 14364
rect 16940 13906 16996 13916
rect 18060 13972 18116 14476
rect 18060 13878 18116 13916
rect 18508 13970 18564 14588
rect 18620 15036 19012 15092
rect 18620 14642 18676 15036
rect 18620 14590 18622 14642
rect 18674 14590 18676 14642
rect 18620 14578 18676 14590
rect 18508 13918 18510 13970
rect 18562 13918 18564 13970
rect 18508 13906 18564 13918
rect 18956 14532 19012 14542
rect 19516 14532 19572 14542
rect 18956 14530 19572 14532
rect 18956 14478 18958 14530
rect 19010 14478 19518 14530
rect 19570 14478 19572 14530
rect 18956 14476 19572 14478
rect 18956 13972 19012 14476
rect 19516 14466 19572 14476
rect 20076 14532 20132 14542
rect 20188 14532 20244 15820
rect 20300 15876 20356 18172
rect 20412 17668 20468 18622
rect 20636 18562 20692 18574
rect 20636 18510 20638 18562
rect 20690 18510 20692 18562
rect 20412 17602 20468 17612
rect 20524 18338 20580 18350
rect 20524 18286 20526 18338
rect 20578 18286 20580 18338
rect 20524 16994 20580 18286
rect 20636 18228 20692 18510
rect 20636 18162 20692 18172
rect 20636 17780 20692 17790
rect 20748 17780 20804 20636
rect 21420 20626 21476 20638
rect 20860 20468 20916 20478
rect 21532 20468 21588 23492
rect 21644 21140 21700 23772
rect 21868 23826 21924 23996
rect 21868 23774 21870 23826
rect 21922 23774 21924 23826
rect 21868 23762 21924 23774
rect 21868 22708 21924 22718
rect 21868 22258 21924 22652
rect 21868 22206 21870 22258
rect 21922 22206 21924 22258
rect 21868 22194 21924 22206
rect 21756 21812 21812 21822
rect 21756 21718 21812 21756
rect 21644 21084 21812 21140
rect 21644 20916 21700 20926
rect 21644 20802 21700 20860
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21644 20738 21700 20750
rect 20860 19684 20916 20412
rect 21420 20412 21588 20468
rect 21308 20018 21364 20030
rect 21308 19966 21310 20018
rect 21362 19966 21364 20018
rect 21084 19908 21140 19918
rect 21308 19908 21364 19966
rect 21420 20020 21476 20412
rect 21756 20244 21812 21084
rect 21644 20188 21812 20244
rect 21868 20692 21924 20702
rect 21532 20132 21588 20142
rect 21532 20038 21588 20076
rect 21420 19954 21476 19964
rect 21140 19852 21364 19908
rect 21084 19814 21140 19852
rect 20860 18674 20916 19628
rect 21420 19348 21476 19358
rect 21420 19234 21476 19292
rect 21420 19182 21422 19234
rect 21474 19182 21476 19234
rect 21420 19170 21476 19182
rect 21532 19124 21588 19134
rect 21532 19030 21588 19068
rect 21644 18900 21700 20188
rect 20860 18622 20862 18674
rect 20914 18622 20916 18674
rect 20860 18452 20916 18622
rect 21084 18844 21700 18900
rect 21756 20018 21812 20030
rect 21756 19966 21758 20018
rect 21810 19966 21812 20018
rect 20916 18396 21028 18452
rect 20860 18386 20916 18396
rect 20636 17778 20804 17780
rect 20636 17726 20638 17778
rect 20690 17726 20804 17778
rect 20636 17724 20804 17726
rect 20636 17714 20692 17724
rect 20972 17668 21028 18396
rect 20972 17602 21028 17612
rect 20524 16942 20526 16994
rect 20578 16942 20580 16994
rect 20524 16930 20580 16942
rect 20748 17444 20804 17454
rect 20412 16882 20468 16894
rect 20412 16830 20414 16882
rect 20466 16830 20468 16882
rect 20412 16210 20468 16830
rect 20748 16882 20804 17388
rect 20748 16830 20750 16882
rect 20802 16830 20804 16882
rect 20748 16818 20804 16830
rect 21084 16660 21140 18844
rect 21756 18676 21812 19966
rect 21868 19348 21924 20636
rect 21980 20130 22036 26796
rect 22204 26628 22260 26638
rect 22428 26628 22484 27244
rect 22876 26908 22932 29484
rect 22988 28980 23044 28990
rect 22988 28754 23044 28924
rect 23212 28866 23268 37212
rect 23324 37202 23380 37212
rect 25676 37268 25732 37278
rect 25900 37268 25956 37326
rect 26236 37268 26292 37278
rect 25676 37266 25844 37268
rect 25676 37214 25678 37266
rect 25730 37214 25844 37266
rect 25676 37212 25844 37214
rect 25900 37266 26292 37268
rect 25900 37214 26238 37266
rect 26290 37214 26292 37266
rect 25900 37212 26292 37214
rect 25676 37202 25732 37212
rect 23436 33122 23492 33134
rect 23436 33070 23438 33122
rect 23490 33070 23492 33122
rect 23436 32788 23492 33070
rect 23436 32732 23940 32788
rect 23436 32562 23492 32574
rect 23436 32510 23438 32562
rect 23490 32510 23492 32562
rect 23436 31892 23492 32510
rect 23884 32452 23940 32732
rect 24332 32452 24388 32462
rect 23884 32450 24388 32452
rect 23884 32398 23886 32450
rect 23938 32398 24334 32450
rect 24386 32398 24388 32450
rect 23884 32396 24388 32398
rect 23884 32386 23940 32396
rect 23436 31826 23492 31836
rect 23772 32338 23828 32350
rect 23772 32286 23774 32338
rect 23826 32286 23828 32338
rect 23772 31780 23828 32286
rect 23548 31724 23828 31780
rect 23884 31778 23940 31790
rect 23884 31726 23886 31778
rect 23938 31726 23940 31778
rect 23436 31556 23492 31566
rect 23548 31556 23604 31724
rect 23436 31554 23604 31556
rect 23436 31502 23438 31554
rect 23490 31502 23604 31554
rect 23436 31500 23604 31502
rect 23660 31556 23716 31566
rect 23436 31108 23492 31500
rect 23660 31462 23716 31500
rect 23772 31554 23828 31566
rect 23772 31502 23774 31554
rect 23826 31502 23828 31554
rect 23436 31014 23492 31052
rect 23436 30660 23492 30670
rect 23436 30548 23492 30604
rect 23436 30492 23604 30548
rect 23324 30436 23380 30446
rect 23380 30380 23492 30436
rect 23324 30370 23380 30380
rect 23324 29988 23380 29998
rect 23324 29894 23380 29932
rect 23436 29764 23492 30380
rect 23324 29708 23492 29764
rect 23324 29538 23380 29708
rect 23548 29652 23604 30492
rect 23324 29486 23326 29538
rect 23378 29486 23380 29538
rect 23324 29474 23380 29486
rect 23436 29596 23604 29652
rect 23436 29538 23492 29596
rect 23436 29486 23438 29538
rect 23490 29486 23492 29538
rect 23212 28814 23214 28866
rect 23266 28814 23268 28866
rect 23212 28802 23268 28814
rect 22988 28702 22990 28754
rect 23042 28702 23044 28754
rect 22988 28690 23044 28702
rect 23324 27860 23380 27870
rect 22988 27746 23044 27758
rect 22988 27694 22990 27746
rect 23042 27694 23044 27746
rect 22988 27636 23044 27694
rect 22988 27570 23044 27580
rect 23100 27634 23156 27646
rect 23100 27582 23102 27634
rect 23154 27582 23156 27634
rect 23100 27412 23156 27582
rect 23100 27356 23268 27412
rect 23100 27188 23156 27198
rect 23100 27094 23156 27132
rect 22876 26852 23044 26908
rect 22260 26572 22372 26628
rect 22204 26562 22260 26572
rect 22316 26514 22372 26572
rect 22428 26562 22484 26572
rect 22316 26462 22318 26514
rect 22370 26462 22372 26514
rect 22316 26450 22372 26462
rect 22876 26516 22932 26526
rect 22876 26422 22932 26460
rect 22652 26402 22708 26414
rect 22652 26350 22654 26402
rect 22706 26350 22708 26402
rect 22540 26066 22596 26078
rect 22540 26014 22542 26066
rect 22594 26014 22596 26066
rect 22092 25172 22148 25182
rect 22092 24946 22148 25116
rect 22092 24894 22094 24946
rect 22146 24894 22148 24946
rect 22092 24882 22148 24894
rect 22204 23268 22260 23278
rect 22204 22146 22260 23212
rect 22428 23268 22484 23278
rect 22428 23174 22484 23212
rect 22316 23156 22372 23166
rect 22316 23062 22372 23100
rect 22428 22260 22484 22270
rect 22204 22094 22206 22146
rect 22258 22094 22260 22146
rect 22204 22082 22260 22094
rect 22316 22258 22484 22260
rect 22316 22206 22430 22258
rect 22482 22206 22484 22258
rect 22316 22204 22484 22206
rect 22204 21362 22260 21374
rect 22204 21310 22206 21362
rect 22258 21310 22260 21362
rect 22092 20916 22148 20926
rect 22092 20802 22148 20860
rect 22092 20750 22094 20802
rect 22146 20750 22148 20802
rect 22092 20738 22148 20750
rect 22204 20580 22260 21310
rect 22316 21026 22372 22204
rect 22428 22194 22484 22204
rect 22428 21588 22484 21598
rect 22540 21588 22596 26014
rect 22652 24724 22708 26350
rect 22764 24948 22820 24958
rect 22764 24854 22820 24892
rect 22652 24658 22708 24668
rect 22652 23714 22708 23726
rect 22652 23662 22654 23714
rect 22706 23662 22708 23714
rect 22652 22370 22708 23662
rect 22988 23156 23044 26852
rect 23212 26290 23268 27356
rect 23324 27076 23380 27804
rect 23324 27010 23380 27020
rect 23212 26238 23214 26290
rect 23266 26238 23268 26290
rect 23212 26226 23268 26238
rect 23324 26740 23380 26750
rect 23324 26290 23380 26684
rect 23324 26238 23326 26290
rect 23378 26238 23380 26290
rect 23324 26226 23380 26238
rect 23212 24724 23268 24734
rect 22988 23090 23044 23100
rect 23100 24164 23156 24174
rect 22652 22318 22654 22370
rect 22706 22318 22708 22370
rect 22652 22306 22708 22318
rect 22764 23042 22820 23054
rect 22764 22990 22766 23042
rect 22818 22990 22820 23042
rect 22428 21586 22596 21588
rect 22428 21534 22430 21586
rect 22482 21534 22596 21586
rect 22428 21532 22596 21534
rect 22652 21812 22708 21822
rect 22652 21586 22708 21756
rect 22652 21534 22654 21586
rect 22706 21534 22708 21586
rect 22428 21522 22484 21532
rect 22316 20974 22318 21026
rect 22370 20974 22372 21026
rect 22316 20962 22372 20974
rect 22428 21364 22484 21374
rect 22204 20514 22260 20524
rect 22428 20132 22484 21308
rect 22540 20804 22596 20814
rect 22652 20804 22708 21534
rect 22764 21140 22820 22990
rect 22876 22484 22932 22494
rect 22876 21698 22932 22428
rect 23100 22036 23156 24108
rect 23100 21970 23156 21980
rect 22876 21646 22878 21698
rect 22930 21646 22932 21698
rect 22876 21634 22932 21646
rect 22764 21084 23044 21140
rect 22540 20802 22708 20804
rect 22540 20750 22542 20802
rect 22594 20750 22708 20802
rect 22540 20748 22708 20750
rect 22764 20916 22820 20926
rect 22540 20738 22596 20748
rect 22764 20690 22820 20860
rect 22764 20638 22766 20690
rect 22818 20638 22820 20690
rect 22764 20626 22820 20638
rect 22876 20690 22932 20702
rect 22876 20638 22878 20690
rect 22930 20638 22932 20690
rect 22876 20580 22932 20638
rect 22876 20514 22932 20524
rect 21980 20078 21982 20130
rect 22034 20078 22036 20130
rect 21980 20066 22036 20078
rect 22204 20076 22484 20132
rect 22652 20468 22708 20478
rect 22092 19908 22148 19918
rect 22092 19814 22148 19852
rect 21868 19282 21924 19292
rect 21980 19122 22036 19134
rect 21980 19070 21982 19122
rect 22034 19070 22036 19122
rect 21980 19012 22036 19070
rect 21980 18946 22036 18956
rect 21196 18620 21812 18676
rect 21196 17106 21252 18620
rect 22092 18562 22148 18574
rect 22092 18510 22094 18562
rect 22146 18510 22148 18562
rect 21644 18452 21700 18462
rect 21308 18450 21700 18452
rect 21308 18398 21646 18450
rect 21698 18398 21700 18450
rect 21308 18396 21700 18398
rect 21308 18340 21364 18396
rect 21644 18386 21700 18396
rect 21980 18450 22036 18462
rect 21980 18398 21982 18450
rect 22034 18398 22036 18450
rect 21308 18274 21364 18284
rect 21420 18116 21476 18126
rect 21196 17054 21198 17106
rect 21250 17054 21252 17106
rect 21196 17042 21252 17054
rect 21308 17892 21364 17902
rect 21308 17108 21364 17836
rect 21308 16772 21364 17052
rect 20748 16604 21140 16660
rect 21196 16716 21364 16772
rect 20412 16158 20414 16210
rect 20466 16158 20468 16210
rect 20412 16146 20468 16158
rect 20524 16436 20580 16446
rect 20300 15782 20356 15820
rect 20524 16098 20580 16380
rect 20524 16046 20526 16098
rect 20578 16046 20580 16098
rect 20524 15652 20580 16046
rect 20748 16100 20804 16604
rect 20748 16006 20804 16044
rect 20300 15596 20580 15652
rect 20300 15314 20356 15596
rect 20300 15262 20302 15314
rect 20354 15262 20356 15314
rect 20300 15250 20356 15262
rect 20524 15428 20580 15438
rect 20524 15314 20580 15372
rect 20524 15262 20526 15314
rect 20578 15262 20580 15314
rect 20524 15250 20580 15262
rect 21196 15314 21252 16716
rect 21196 15262 21198 15314
rect 21250 15262 21252 15314
rect 21196 15250 21252 15262
rect 21308 16098 21364 16110
rect 21308 16046 21310 16098
rect 21362 16046 21364 16098
rect 21308 15148 21364 16046
rect 21420 15538 21476 18060
rect 21644 18004 21700 18014
rect 21644 17668 21700 17948
rect 21980 17780 22036 18398
rect 21980 17714 22036 17724
rect 21644 17666 21812 17668
rect 21644 17614 21646 17666
rect 21698 17614 21812 17666
rect 21644 17612 21812 17614
rect 21644 17602 21700 17612
rect 21644 17220 21700 17230
rect 21532 16436 21588 16446
rect 21532 16098 21588 16380
rect 21644 16210 21700 17164
rect 21644 16158 21646 16210
rect 21698 16158 21700 16210
rect 21644 16146 21700 16158
rect 21532 16046 21534 16098
rect 21586 16046 21588 16098
rect 21532 16034 21588 16046
rect 21756 16098 21812 17612
rect 22092 17220 22148 18510
rect 22204 17892 22260 20076
rect 22428 19906 22484 19918
rect 22428 19854 22430 19906
rect 22482 19854 22484 19906
rect 22428 19684 22484 19854
rect 22428 19618 22484 19628
rect 22428 19460 22484 19470
rect 22428 19346 22484 19404
rect 22428 19294 22430 19346
rect 22482 19294 22484 19346
rect 22428 19282 22484 19294
rect 22316 18676 22372 18686
rect 22652 18676 22708 20412
rect 22316 18674 22708 18676
rect 22316 18622 22318 18674
rect 22370 18622 22708 18674
rect 22316 18620 22708 18622
rect 22316 18610 22372 18620
rect 22764 18450 22820 18462
rect 22764 18398 22766 18450
rect 22818 18398 22820 18450
rect 22540 18340 22596 18350
rect 22204 17826 22260 17836
rect 22428 18338 22596 18340
rect 22428 18286 22542 18338
rect 22594 18286 22596 18338
rect 22428 18284 22596 18286
rect 22092 17154 22148 17164
rect 22204 17666 22260 17678
rect 22204 17614 22206 17666
rect 22258 17614 22260 17666
rect 21980 16994 22036 17006
rect 21980 16942 21982 16994
rect 22034 16942 22036 16994
rect 21980 16884 22036 16942
rect 22092 16996 22148 17006
rect 22204 16996 22260 17614
rect 22428 17108 22484 18284
rect 22540 18274 22596 18284
rect 22652 18340 22708 18350
rect 22764 18340 22820 18398
rect 22708 18284 22820 18340
rect 22876 18452 22932 18462
rect 22652 18274 22708 18284
rect 22540 17892 22596 17902
rect 22540 17332 22596 17836
rect 22764 17668 22820 17678
rect 22764 17574 22820 17612
rect 22876 17554 22932 18396
rect 22988 17780 23044 21084
rect 23212 20356 23268 24668
rect 23324 24612 23380 24622
rect 23324 21476 23380 24556
rect 23436 23268 23492 29486
rect 23660 29428 23716 29438
rect 23660 29334 23716 29372
rect 23660 28980 23716 28990
rect 23660 28866 23716 28924
rect 23660 28814 23662 28866
rect 23714 28814 23716 28866
rect 23660 28802 23716 28814
rect 23772 27970 23828 31502
rect 23884 30996 23940 31726
rect 23996 31444 24052 32396
rect 24332 32386 24388 32396
rect 23996 31378 24052 31388
rect 24108 31890 24164 31902
rect 24108 31838 24110 31890
rect 24162 31838 24164 31890
rect 23996 31220 24052 31230
rect 23996 31106 24052 31164
rect 23996 31054 23998 31106
rect 24050 31054 24052 31106
rect 23996 31042 24052 31054
rect 23884 30930 23940 30940
rect 24108 30436 24164 31838
rect 24220 31554 24276 31566
rect 24220 31502 24222 31554
rect 24274 31502 24276 31554
rect 24220 31444 24276 31502
rect 24220 31378 24276 31388
rect 24444 31554 24500 31566
rect 24444 31502 24446 31554
rect 24498 31502 24500 31554
rect 24444 31220 24500 31502
rect 24892 31556 24948 31566
rect 24892 31462 24948 31500
rect 24444 31154 24500 31164
rect 25452 31220 25508 31230
rect 25452 31126 25508 31164
rect 25228 31108 25284 31118
rect 25228 31014 25284 31052
rect 24332 30882 24388 30894
rect 24332 30830 24334 30882
rect 24386 30830 24388 30882
rect 24220 30436 24276 30446
rect 24108 30434 24276 30436
rect 24108 30382 24222 30434
rect 24274 30382 24276 30434
rect 24108 30380 24276 30382
rect 24220 30370 24276 30380
rect 23996 30210 24052 30222
rect 23996 30158 23998 30210
rect 24050 30158 24052 30210
rect 23996 29316 24052 30158
rect 23996 29250 24052 29260
rect 24332 28868 24388 30830
rect 25340 30882 25396 30894
rect 25340 30830 25342 30882
rect 25394 30830 25396 30882
rect 25340 30436 25396 30830
rect 25340 30370 25396 30380
rect 24332 28802 24388 28812
rect 24556 29986 24612 29998
rect 24556 29934 24558 29986
rect 24610 29934 24612 29986
rect 24556 28756 24612 29934
rect 25340 29764 25396 29774
rect 24668 29428 24724 29438
rect 24724 29372 24948 29428
rect 24668 29362 24724 29372
rect 24556 28690 24612 28700
rect 24780 28866 24836 28878
rect 24780 28814 24782 28866
rect 24834 28814 24836 28866
rect 23884 28644 23940 28654
rect 23884 28550 23940 28588
rect 24108 28644 24164 28654
rect 24108 28550 24164 28588
rect 24780 28644 24836 28814
rect 24780 28578 24836 28588
rect 24892 28642 24948 29372
rect 24892 28590 24894 28642
rect 24946 28590 24948 28642
rect 24892 28578 24948 28590
rect 25340 28980 25396 29708
rect 25340 28924 25732 28980
rect 25340 28642 25396 28924
rect 25340 28590 25342 28642
rect 25394 28590 25396 28642
rect 25340 28578 25396 28590
rect 25452 28756 25508 28766
rect 24332 28532 24388 28542
rect 24220 28530 24388 28532
rect 24220 28478 24334 28530
rect 24386 28478 24388 28530
rect 24220 28476 24388 28478
rect 23772 27918 23774 27970
rect 23826 27918 23828 27970
rect 23772 27906 23828 27918
rect 23884 28420 23940 28430
rect 23548 27748 23604 27758
rect 23548 27300 23604 27692
rect 23548 27074 23604 27244
rect 23548 27022 23550 27074
rect 23602 27022 23604 27074
rect 23548 27010 23604 27022
rect 23660 27412 23716 27422
rect 23660 27076 23716 27356
rect 23660 26740 23716 27020
rect 23660 26674 23716 26684
rect 23772 27188 23828 27198
rect 23772 26514 23828 27132
rect 23884 26964 23940 28364
rect 23996 27970 24052 27982
rect 23996 27918 23998 27970
rect 24050 27918 24052 27970
rect 23996 27412 24052 27918
rect 24108 27972 24164 27982
rect 24108 27858 24164 27916
rect 24108 27806 24110 27858
rect 24162 27806 24164 27858
rect 24108 27794 24164 27806
rect 23996 27346 24052 27356
rect 24108 27300 24164 27310
rect 24108 27188 24164 27244
rect 23884 26898 23940 26908
rect 23996 27132 24164 27188
rect 23772 26462 23774 26514
rect 23826 26462 23828 26514
rect 23772 26450 23828 26462
rect 23996 26514 24052 27132
rect 23996 26462 23998 26514
rect 24050 26462 24052 26514
rect 23996 26450 24052 26462
rect 24108 26908 24164 26918
rect 23884 26178 23940 26190
rect 23884 26126 23886 26178
rect 23938 26126 23940 26178
rect 23772 25844 23828 25854
rect 23548 25732 23604 25742
rect 23548 23492 23604 25676
rect 23772 25394 23828 25788
rect 23772 25342 23774 25394
rect 23826 25342 23828 25394
rect 23772 25330 23828 25342
rect 23772 24948 23828 24958
rect 23772 24722 23828 24892
rect 23772 24670 23774 24722
rect 23826 24670 23828 24722
rect 23772 24658 23828 24670
rect 23548 23426 23604 23436
rect 23660 23938 23716 23950
rect 23660 23886 23662 23938
rect 23714 23886 23716 23938
rect 23660 23378 23716 23886
rect 23884 23828 23940 26126
rect 23996 24836 24052 24846
rect 23996 24742 24052 24780
rect 24108 24722 24164 26852
rect 24108 24670 24110 24722
rect 24162 24670 24164 24722
rect 23884 23762 23940 23772
rect 23996 23938 24052 23950
rect 23996 23886 23998 23938
rect 24050 23886 24052 23938
rect 23660 23326 23662 23378
rect 23714 23326 23716 23378
rect 23660 23314 23716 23326
rect 23436 23202 23492 23212
rect 23772 23266 23828 23278
rect 23772 23214 23774 23266
rect 23826 23214 23828 23266
rect 23548 22372 23604 22382
rect 23548 22278 23604 22316
rect 23772 22260 23828 23214
rect 23996 23156 24052 23886
rect 23884 22484 23940 22494
rect 23884 22370 23940 22428
rect 23884 22318 23886 22370
rect 23938 22318 23940 22370
rect 23884 22306 23940 22318
rect 23996 22372 24052 23100
rect 24108 22820 24164 24670
rect 24108 22754 24164 22764
rect 24220 22482 24276 28476
rect 24332 28466 24388 28476
rect 24668 28530 24724 28542
rect 24668 28478 24670 28530
rect 24722 28478 24724 28530
rect 24332 27972 24388 27982
rect 24332 26514 24388 27916
rect 24668 26908 24724 28478
rect 25116 28418 25172 28430
rect 25116 28366 25118 28418
rect 25170 28366 25172 28418
rect 25116 27972 25172 28366
rect 25116 27906 25172 27916
rect 25228 27860 25284 27870
rect 25228 27766 25284 27804
rect 25340 27524 25396 27534
rect 24780 27188 24836 27198
rect 24780 27074 24836 27132
rect 24780 27022 24782 27074
rect 24834 27022 24836 27074
rect 24780 27010 24836 27022
rect 24332 26462 24334 26514
rect 24386 26462 24388 26514
rect 24332 26450 24388 26462
rect 24556 26852 24724 26908
rect 24332 24722 24388 24734
rect 24332 24670 24334 24722
rect 24386 24670 24388 24722
rect 24332 24612 24388 24670
rect 24332 24546 24388 24556
rect 24556 24052 24612 26852
rect 24668 26402 24724 26414
rect 24668 26350 24670 26402
rect 24722 26350 24724 26402
rect 24668 25284 24724 26350
rect 25228 26402 25284 26414
rect 25228 26350 25230 26402
rect 25282 26350 25284 26402
rect 25228 26180 25284 26350
rect 25228 26114 25284 26124
rect 25340 25732 25396 27468
rect 25228 25676 25396 25732
rect 24892 25508 24948 25518
rect 24892 25414 24948 25452
rect 24668 25218 24724 25228
rect 25116 25284 25172 25294
rect 24780 24500 24836 24510
rect 24780 24406 24836 24444
rect 24556 23996 24724 24052
rect 24556 23828 24612 23838
rect 24556 23734 24612 23772
rect 24332 23492 24388 23502
rect 24332 23268 24388 23436
rect 24332 23174 24388 23212
rect 24556 23154 24612 23166
rect 24556 23102 24558 23154
rect 24610 23102 24612 23154
rect 24556 22594 24612 23102
rect 24556 22542 24558 22594
rect 24610 22542 24612 22594
rect 24556 22530 24612 22542
rect 24220 22430 24222 22482
rect 24274 22430 24276 22482
rect 24220 22418 24276 22430
rect 24108 22372 24164 22382
rect 23996 22316 24108 22372
rect 24108 22306 24164 22316
rect 23660 22204 23828 22260
rect 24332 22260 24388 22270
rect 23660 22148 23716 22204
rect 23548 21700 23604 21710
rect 23660 21700 23716 22092
rect 24108 22146 24164 22158
rect 24108 22094 24110 22146
rect 24162 22094 24164 22146
rect 24108 21812 24164 22094
rect 23604 21644 23716 21700
rect 23772 21756 24164 21812
rect 23548 21634 23604 21644
rect 23324 21420 23492 21476
rect 23100 20300 23268 20356
rect 23324 20580 23380 20590
rect 23100 18788 23156 20300
rect 23212 19348 23268 19358
rect 23212 19254 23268 19292
rect 23100 18732 23268 18788
rect 23100 18228 23156 18238
rect 23100 18134 23156 18172
rect 22988 17724 23156 17780
rect 22876 17502 22878 17554
rect 22930 17502 22932 17554
rect 22540 17276 22820 17332
rect 22428 17052 22708 17108
rect 22148 16940 22260 16996
rect 22092 16930 22148 16940
rect 21980 16818 22036 16828
rect 22092 16548 22148 16558
rect 21756 16046 21758 16098
rect 21810 16046 21812 16098
rect 21420 15486 21422 15538
rect 21474 15486 21476 15538
rect 21420 15474 21476 15486
rect 21644 15876 21700 15886
rect 21644 15426 21700 15820
rect 21644 15374 21646 15426
rect 21698 15374 21700 15426
rect 21644 15362 21700 15374
rect 21756 15148 21812 16046
rect 21868 16100 21924 16110
rect 21868 16006 21924 16044
rect 22092 15988 22148 16492
rect 22204 16100 22260 16940
rect 22428 16882 22484 16894
rect 22428 16830 22430 16882
rect 22482 16830 22484 16882
rect 22428 16322 22484 16830
rect 22428 16270 22430 16322
rect 22482 16270 22484 16322
rect 22428 16258 22484 16270
rect 22540 16100 22596 16110
rect 22204 16044 22540 16100
rect 22540 16006 22596 16044
rect 22092 15932 22484 15988
rect 22428 15876 22484 15932
rect 22428 15782 22484 15820
rect 22092 15540 22148 15550
rect 22092 15446 22148 15484
rect 20132 14476 20244 14532
rect 20860 15092 21364 15148
rect 21420 15092 21812 15148
rect 22316 15316 22372 15326
rect 20860 14642 20916 15092
rect 20860 14590 20862 14642
rect 20914 14590 20916 14642
rect 20076 14466 20132 14476
rect 19852 14308 19908 14318
rect 19628 14252 19852 14308
rect 19628 14196 19684 14252
rect 19852 14242 19908 14252
rect 20860 14308 20916 14590
rect 21420 14642 21476 15092
rect 21756 15036 22148 15092
rect 21980 14868 22036 14878
rect 21980 14756 22036 14812
rect 21420 14590 21422 14642
rect 21474 14590 21476 14642
rect 21420 14578 21476 14590
rect 21868 14754 22036 14756
rect 21868 14702 21982 14754
rect 22034 14702 22036 14754
rect 21868 14700 22036 14702
rect 20860 14242 20916 14252
rect 21868 14308 21924 14700
rect 21980 14690 22036 14700
rect 22092 14644 22148 15036
rect 22204 14644 22260 14654
rect 22092 14588 22204 14644
rect 22092 14530 22148 14588
rect 22204 14578 22260 14588
rect 22092 14478 22094 14530
rect 22146 14478 22148 14530
rect 22092 14466 22148 14478
rect 21980 14420 22036 14430
rect 21980 14326 22036 14364
rect 21868 14242 21924 14252
rect 19628 14130 19684 14140
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 18956 13878 19012 13916
rect 13692 13860 13748 13870
rect 13580 13804 13692 13860
rect 13244 13766 13300 13804
rect 13692 13766 13748 13804
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 8876 11442 8932 11452
rect 22316 11396 22372 15260
rect 22540 14644 22596 14654
rect 22540 14550 22596 14588
rect 22652 14420 22708 17052
rect 22764 15538 22820 17276
rect 22876 17108 22932 17502
rect 22876 17042 22932 17052
rect 22988 17556 23044 17566
rect 22988 16994 23044 17500
rect 22988 16942 22990 16994
rect 23042 16942 23044 16994
rect 22988 16930 23044 16942
rect 23100 16772 23156 17724
rect 23212 17778 23268 18732
rect 23212 17726 23214 17778
rect 23266 17726 23268 17778
rect 23212 17714 23268 17726
rect 22764 15486 22766 15538
rect 22818 15486 22820 15538
rect 22764 15428 22820 15486
rect 22764 15362 22820 15372
rect 22876 16716 23156 16772
rect 22652 14354 22708 14364
rect 22876 11620 22932 16716
rect 23100 16100 23156 16138
rect 23100 16034 23156 16044
rect 23212 15986 23268 15998
rect 23212 15934 23214 15986
rect 23266 15934 23268 15986
rect 23100 15876 23156 15886
rect 23212 15876 23268 15934
rect 23156 15820 23268 15876
rect 23100 15810 23156 15820
rect 23324 15652 23380 20524
rect 23100 15596 23380 15652
rect 23100 14868 23156 15596
rect 23212 15428 23268 15438
rect 23212 15334 23268 15372
rect 23324 15316 23380 15326
rect 23436 15316 23492 21420
rect 23772 21474 23828 21756
rect 24220 21700 24276 21710
rect 24220 21606 24276 21644
rect 23996 21588 24052 21598
rect 23996 21494 24052 21532
rect 24332 21586 24388 22204
rect 24556 22146 24612 22158
rect 24556 22094 24558 22146
rect 24610 22094 24612 22146
rect 24556 22036 24612 22094
rect 24556 21970 24612 21980
rect 24332 21534 24334 21586
rect 24386 21534 24388 21586
rect 24332 21522 24388 21534
rect 23772 21422 23774 21474
rect 23826 21422 23828 21474
rect 23548 20018 23604 20030
rect 23548 19966 23550 20018
rect 23602 19966 23604 20018
rect 23548 18676 23604 19966
rect 23548 18610 23604 18620
rect 23660 19348 23716 19358
rect 23548 18452 23604 18462
rect 23660 18452 23716 19292
rect 23772 18900 23828 21422
rect 24668 20916 24724 23996
rect 25116 23044 25172 25228
rect 25228 24948 25284 25676
rect 25228 24882 25284 24892
rect 25340 25506 25396 25518
rect 25340 25454 25342 25506
rect 25394 25454 25396 25506
rect 25228 24724 25284 24734
rect 25228 24630 25284 24668
rect 25340 24610 25396 25454
rect 25340 24558 25342 24610
rect 25394 24558 25396 24610
rect 25340 24546 25396 24558
rect 25452 23044 25508 28700
rect 25676 28642 25732 28924
rect 25676 28590 25678 28642
rect 25730 28590 25732 28642
rect 25676 28578 25732 28590
rect 25788 28644 25844 37212
rect 26236 37202 26292 37212
rect 26908 32676 26964 32686
rect 26124 28868 26180 28878
rect 25788 28588 25956 28644
rect 25564 27970 25620 27982
rect 25564 27918 25566 27970
rect 25618 27918 25620 27970
rect 25564 27860 25620 27918
rect 25564 27794 25620 27804
rect 25788 27858 25844 27870
rect 25788 27806 25790 27858
rect 25842 27806 25844 27858
rect 25788 26290 25844 27806
rect 25788 26238 25790 26290
rect 25842 26238 25844 26290
rect 25788 26226 25844 26238
rect 25788 25396 25844 25406
rect 25788 25302 25844 25340
rect 25564 23380 25620 23390
rect 25900 23380 25956 28588
rect 26124 28084 26180 28812
rect 26236 28642 26292 28654
rect 26236 28590 26238 28642
rect 26290 28590 26292 28642
rect 26236 28308 26292 28590
rect 26236 28242 26292 28252
rect 26124 28028 26292 28084
rect 26012 27970 26068 27982
rect 26012 27918 26014 27970
rect 26066 27918 26068 27970
rect 26012 27524 26068 27918
rect 26124 27860 26180 27870
rect 26124 27766 26180 27804
rect 26236 27524 26292 28028
rect 26572 27746 26628 27758
rect 26572 27694 26574 27746
rect 26626 27694 26628 27746
rect 26012 27458 26068 27468
rect 26124 27468 26292 27524
rect 26348 27524 26404 27534
rect 26572 27524 26628 27694
rect 26404 27468 26628 27524
rect 25564 23378 25956 23380
rect 25564 23326 25566 23378
rect 25618 23326 25956 23378
rect 25564 23324 25956 23326
rect 26012 27298 26068 27310
rect 26012 27246 26014 27298
rect 26066 27246 26068 27298
rect 25564 23314 25620 23324
rect 26012 23156 26068 27246
rect 26124 24834 26180 27468
rect 26348 27458 26404 27468
rect 26236 27076 26292 27086
rect 26236 26982 26292 27020
rect 26348 26964 26404 26974
rect 26908 26964 26964 32620
rect 28140 28308 28196 28318
rect 26348 26962 26964 26964
rect 26348 26910 26350 26962
rect 26402 26910 26964 26962
rect 26348 26908 26964 26910
rect 27356 27860 27412 27870
rect 26348 26898 26404 26908
rect 26684 26516 26740 26526
rect 26684 26422 26740 26460
rect 26796 26404 26852 26414
rect 26796 26310 26852 26348
rect 26236 26292 26292 26302
rect 27244 26292 27300 26302
rect 26236 26198 26292 26236
rect 27020 26290 27300 26292
rect 27020 26238 27246 26290
rect 27298 26238 27300 26290
rect 27020 26236 27300 26238
rect 26796 25284 26852 25294
rect 27020 25284 27076 26236
rect 27244 26226 27300 26236
rect 27356 26068 27412 27804
rect 27580 26516 27636 26526
rect 27580 26402 27636 26460
rect 27580 26350 27582 26402
rect 27634 26350 27636 26402
rect 27580 26338 27636 26350
rect 28140 26404 28196 28252
rect 28364 27076 28420 27086
rect 28140 26402 28308 26404
rect 28140 26350 28142 26402
rect 28194 26350 28308 26402
rect 28140 26348 28308 26350
rect 28140 26338 28196 26348
rect 26796 25282 27076 25284
rect 26796 25230 26798 25282
rect 26850 25230 27076 25282
rect 26796 25228 27076 25230
rect 27244 26012 27412 26068
rect 27468 26292 27524 26302
rect 27244 25394 27300 26012
rect 27244 25342 27246 25394
rect 27298 25342 27300 25394
rect 26796 25218 26852 25228
rect 26124 24782 26126 24834
rect 26178 24782 26180 24834
rect 26124 24770 26180 24782
rect 27020 24834 27076 24846
rect 27020 24782 27022 24834
rect 27074 24782 27076 24834
rect 26908 24276 26964 24286
rect 26908 23938 26964 24220
rect 26908 23886 26910 23938
rect 26962 23886 26964 23938
rect 26908 23874 26964 23886
rect 26908 23268 26964 23278
rect 25116 22594 25172 22988
rect 25116 22542 25118 22594
rect 25170 22542 25172 22594
rect 25004 22146 25060 22158
rect 25004 22094 25006 22146
rect 25058 22094 25060 22146
rect 25004 22036 25060 22094
rect 25004 21970 25060 21980
rect 24780 21364 24836 21374
rect 24780 21362 25060 21364
rect 24780 21310 24782 21362
rect 24834 21310 25060 21362
rect 24780 21308 25060 21310
rect 24780 21298 24836 21308
rect 24332 20860 24724 20916
rect 23884 20132 23940 20142
rect 23884 20038 23940 20076
rect 24332 20130 24388 20860
rect 24780 20802 24836 20814
rect 24780 20750 24782 20802
rect 24834 20750 24836 20802
rect 24444 20580 24500 20590
rect 24780 20580 24836 20750
rect 24444 20578 24836 20580
rect 24444 20526 24446 20578
rect 24498 20526 24836 20578
rect 24444 20524 24836 20526
rect 24892 20690 24948 20702
rect 24892 20638 24894 20690
rect 24946 20638 24948 20690
rect 24444 20244 24500 20524
rect 24892 20356 24948 20638
rect 24444 20178 24500 20188
rect 24780 20300 24948 20356
rect 24332 20078 24334 20130
rect 24386 20078 24388 20130
rect 24108 19460 24164 19470
rect 24108 19366 24164 19404
rect 23996 19124 24052 19134
rect 23996 19030 24052 19068
rect 24108 19010 24164 19022
rect 24108 18958 24110 19010
rect 24162 18958 24164 19010
rect 24108 18900 24164 18958
rect 23772 18844 24164 18900
rect 23772 18676 23828 18686
rect 23772 18674 23940 18676
rect 23772 18622 23774 18674
rect 23826 18622 23940 18674
rect 23772 18620 23940 18622
rect 23772 18610 23828 18620
rect 23548 18450 23716 18452
rect 23548 18398 23550 18450
rect 23602 18398 23716 18450
rect 23548 18396 23716 18398
rect 23772 18450 23828 18462
rect 23772 18398 23774 18450
rect 23826 18398 23828 18450
rect 23548 18386 23604 18396
rect 23772 15876 23828 18398
rect 23884 18452 23940 18620
rect 23884 18386 23940 18396
rect 23772 15810 23828 15820
rect 23380 15260 23492 15316
rect 23324 15250 23380 15260
rect 23884 15092 23940 15102
rect 23996 15092 24052 18844
rect 24108 18450 24164 18462
rect 24108 18398 24110 18450
rect 24162 18398 24164 18450
rect 24108 18228 24164 18398
rect 24108 17668 24164 18172
rect 24108 17602 24164 17612
rect 24332 16210 24388 20078
rect 24780 20130 24836 20300
rect 24780 20078 24782 20130
rect 24834 20078 24836 20130
rect 24780 20066 24836 20078
rect 25004 20020 25060 21308
rect 25004 19954 25060 19964
rect 25116 19796 25172 22542
rect 24892 19740 25172 19796
rect 25228 22988 25508 23044
rect 25788 23100 26068 23156
rect 26460 23266 26964 23268
rect 26460 23214 26910 23266
rect 26962 23214 26964 23266
rect 26460 23212 26964 23214
rect 26460 23154 26516 23212
rect 26908 23202 26964 23212
rect 27020 23268 27076 24782
rect 27244 24836 27300 25342
rect 27356 25284 27412 25294
rect 27356 25190 27412 25228
rect 27244 24770 27300 24780
rect 27244 24500 27300 24510
rect 27244 23826 27300 24444
rect 27244 23774 27246 23826
rect 27298 23774 27300 23826
rect 27244 23762 27300 23774
rect 27020 23202 27076 23212
rect 26460 23102 26462 23154
rect 26514 23102 26516 23154
rect 24668 19236 24724 19246
rect 24668 19142 24724 19180
rect 24892 19234 24948 19740
rect 24892 19182 24894 19234
rect 24946 19182 24948 19234
rect 24892 19170 24948 19182
rect 25228 19234 25284 22988
rect 25340 22820 25396 22830
rect 25340 22370 25396 22764
rect 25340 22318 25342 22370
rect 25394 22318 25396 22370
rect 25340 22306 25396 22318
rect 25452 22148 25508 22158
rect 25452 22054 25508 22092
rect 25676 22146 25732 22158
rect 25676 22094 25678 22146
rect 25730 22094 25732 22146
rect 25564 22036 25620 22046
rect 25564 21698 25620 21980
rect 25564 21646 25566 21698
rect 25618 21646 25620 21698
rect 25564 21634 25620 21646
rect 25676 20804 25732 22094
rect 25788 21588 25844 23100
rect 26460 23090 26516 23102
rect 27356 23156 27412 23166
rect 27468 23156 27524 26236
rect 27580 25284 27636 25294
rect 27580 25282 27748 25284
rect 27580 25230 27582 25282
rect 27634 25230 27748 25282
rect 27580 25228 27748 25230
rect 27580 25218 27636 25228
rect 27356 23154 27524 23156
rect 27356 23102 27358 23154
rect 27410 23102 27524 23154
rect 27356 23100 27524 23102
rect 27580 23156 27636 23166
rect 27692 23156 27748 25228
rect 28140 24052 28196 24062
rect 28140 23958 28196 23996
rect 27804 23828 27860 23838
rect 27804 23826 27972 23828
rect 27804 23774 27806 23826
rect 27858 23774 27972 23826
rect 27804 23772 27972 23774
rect 27804 23762 27860 23772
rect 27580 23154 27748 23156
rect 27580 23102 27582 23154
rect 27634 23102 27748 23154
rect 27580 23100 27748 23102
rect 27804 23156 27860 23166
rect 27356 23090 27412 23100
rect 27580 23090 27636 23100
rect 27804 23062 27860 23100
rect 26684 23044 26740 23054
rect 26684 23042 26852 23044
rect 26684 22990 26686 23042
rect 26738 22990 26852 23042
rect 26684 22988 26852 22990
rect 26684 22978 26740 22988
rect 26012 22930 26068 22942
rect 26012 22878 26014 22930
rect 26066 22878 26068 22930
rect 26012 22820 26068 22878
rect 26012 22754 26068 22764
rect 26124 22932 26180 22942
rect 25788 21522 25844 21532
rect 25900 22370 25956 22382
rect 25900 22318 25902 22370
rect 25954 22318 25956 22370
rect 25676 20738 25732 20748
rect 25788 21364 25844 21374
rect 25900 21364 25956 22318
rect 25788 21362 25956 21364
rect 25788 21310 25790 21362
rect 25842 21310 25956 21362
rect 25788 21308 25956 21310
rect 26012 21364 26068 21374
rect 26124 21364 26180 22876
rect 26236 22932 26292 22942
rect 26460 22932 26516 22942
rect 26236 22930 26404 22932
rect 26236 22878 26238 22930
rect 26290 22878 26404 22930
rect 26236 22876 26404 22878
rect 26236 22866 26292 22876
rect 26236 21588 26292 21598
rect 26236 21494 26292 21532
rect 26012 21362 26180 21364
rect 26012 21310 26014 21362
rect 26066 21310 26180 21362
rect 26012 21308 26180 21310
rect 25788 20468 25844 21308
rect 26012 21298 26068 21308
rect 25788 20402 25844 20412
rect 26124 20020 26180 20030
rect 25676 20018 26180 20020
rect 25676 19966 26126 20018
rect 26178 19966 26180 20018
rect 25676 19964 26180 19966
rect 25676 19458 25732 19964
rect 26124 19954 26180 19964
rect 26236 19908 26292 19918
rect 26348 19908 26404 22876
rect 26460 22258 26516 22876
rect 26572 22820 26628 22830
rect 26628 22764 26740 22820
rect 26572 22754 26628 22764
rect 26460 22206 26462 22258
rect 26514 22206 26516 22258
rect 26460 22194 26516 22206
rect 26684 21810 26740 22764
rect 26684 21758 26686 21810
rect 26738 21758 26740 21810
rect 26684 21746 26740 21758
rect 26796 21812 26852 22988
rect 27916 22932 27972 23772
rect 28140 23268 28196 23278
rect 28140 23154 28196 23212
rect 28140 23102 28142 23154
rect 28194 23102 28196 23154
rect 28140 23090 28196 23102
rect 28140 22932 28196 22942
rect 27916 22876 28140 22932
rect 27692 22370 27748 22382
rect 27692 22318 27694 22370
rect 27746 22318 27748 22370
rect 27692 22036 27748 22318
rect 27692 21970 27748 21980
rect 26796 21746 26852 21756
rect 27468 21698 27524 21710
rect 27468 21646 27470 21698
rect 27522 21646 27524 21698
rect 27356 21588 27412 21598
rect 26796 20804 26852 20814
rect 26796 20710 26852 20748
rect 27356 20690 27412 21532
rect 27468 20914 27524 21646
rect 28140 21586 28196 22876
rect 28252 22820 28308 26348
rect 28364 24722 28420 27020
rect 28476 26404 28532 26414
rect 28476 26310 28532 26348
rect 28364 24670 28366 24722
rect 28418 24670 28420 24722
rect 28364 24658 28420 24670
rect 28700 23380 28756 37996
rect 29036 38050 29092 38062
rect 29036 37998 29038 38050
rect 29090 37998 29092 38050
rect 29036 31948 29092 37998
rect 28700 23314 28756 23324
rect 28812 31892 29092 31948
rect 32844 38050 32900 38062
rect 32844 37998 32846 38050
rect 32898 37998 32900 38050
rect 28364 23154 28420 23166
rect 28364 23102 28366 23154
rect 28418 23102 28420 23154
rect 28364 23044 28420 23102
rect 28364 22978 28420 22988
rect 28476 23154 28532 23166
rect 28476 23102 28478 23154
rect 28530 23102 28532 23154
rect 28252 22764 28420 22820
rect 28140 21534 28142 21586
rect 28194 21534 28196 21586
rect 28140 21522 28196 21534
rect 28252 22146 28308 22158
rect 28252 22094 28254 22146
rect 28306 22094 28308 22146
rect 28252 21924 28308 22094
rect 28364 22036 28420 22764
rect 28476 22484 28532 23102
rect 28476 22418 28532 22428
rect 28364 21980 28756 22036
rect 28252 21868 28644 21924
rect 27468 20862 27470 20914
rect 27522 20862 27524 20914
rect 27468 20850 27524 20862
rect 27356 20638 27358 20690
rect 27410 20638 27412 20690
rect 27356 20626 27412 20638
rect 28252 20188 28308 21868
rect 28588 21586 28644 21868
rect 28588 21534 28590 21586
rect 28642 21534 28644 21586
rect 28588 21522 28644 21534
rect 28700 21698 28756 21980
rect 28700 21646 28702 21698
rect 28754 21646 28756 21698
rect 28700 20916 28756 21646
rect 28812 21474 28868 31892
rect 30380 29876 30436 29886
rect 30268 25508 30324 25518
rect 28924 22932 28980 22942
rect 28924 22838 28980 22876
rect 28812 21422 28814 21474
rect 28866 21422 28868 21474
rect 28812 21410 28868 21422
rect 28700 20850 28756 20860
rect 26292 19852 26404 19908
rect 26684 20130 26740 20142
rect 26684 20078 26686 20130
rect 26738 20078 26740 20130
rect 26236 19842 26292 19852
rect 26684 19796 26740 20078
rect 27916 20132 28308 20188
rect 27916 20130 27972 20132
rect 27916 20078 27918 20130
rect 27970 20078 27972 20130
rect 27916 20066 27972 20078
rect 27692 20020 27748 20030
rect 27692 19926 27748 19964
rect 29484 19908 29540 19918
rect 29484 19814 29540 19852
rect 26684 19730 26740 19740
rect 25676 19406 25678 19458
rect 25730 19406 25732 19458
rect 25676 19394 25732 19406
rect 25228 19182 25230 19234
rect 25282 19182 25284 19234
rect 25228 19170 25284 19182
rect 25004 19122 25060 19134
rect 25004 19070 25006 19122
rect 25058 19070 25060 19122
rect 24556 18564 24612 18574
rect 24444 17892 24500 17902
rect 24444 17666 24500 17836
rect 24444 17614 24446 17666
rect 24498 17614 24500 17666
rect 24444 17602 24500 17614
rect 24556 16882 24612 18508
rect 25004 18452 25060 19070
rect 25004 18386 25060 18396
rect 25676 17668 25732 17678
rect 25676 17574 25732 17612
rect 24556 16830 24558 16882
rect 24610 16830 24612 16882
rect 24556 16818 24612 16830
rect 24780 16772 24836 16782
rect 24780 16678 24836 16716
rect 30268 16772 30324 25452
rect 30380 20132 30436 29820
rect 32844 26404 32900 37998
rect 36428 38050 36484 38062
rect 36428 37998 36430 38050
rect 36482 37998 36484 38050
rect 32844 26338 32900 26348
rect 34412 37156 34468 37166
rect 34412 24052 34468 37100
rect 35980 37156 36036 37166
rect 35980 37062 36036 37100
rect 36428 37156 36484 37998
rect 39452 37378 39508 41200
rect 39452 37326 39454 37378
rect 39506 37326 39508 37378
rect 39452 37314 39508 37326
rect 37660 37266 37716 37278
rect 37660 37214 37662 37266
rect 37714 37214 37716 37266
rect 36428 37090 36484 37100
rect 37436 37156 37492 37166
rect 37660 37156 37716 37214
rect 37436 37154 37716 37156
rect 37436 37102 37438 37154
rect 37490 37102 37716 37154
rect 37436 37100 37716 37102
rect 37436 37090 37492 37100
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34412 23986 34468 23996
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 30380 20066 30436 20076
rect 37660 19908 37716 37100
rect 37660 19842 37716 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 30268 16706 30324 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 24332 16158 24334 16210
rect 24386 16158 24388 16210
rect 24332 16146 24388 16158
rect 23940 15036 24052 15092
rect 24668 16098 24724 16110
rect 24668 16046 24670 16098
rect 24722 16046 24724 16098
rect 24668 15092 24724 16046
rect 26012 16098 26068 16110
rect 26012 16046 26014 16098
rect 26066 16046 26068 16098
rect 26012 15428 26068 16046
rect 26012 15362 26068 15372
rect 23884 15026 23940 15036
rect 24668 15026 24724 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 23100 14802 23156 14812
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 22876 11554 22932 11564
rect 22316 11330 22372 11340
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 6300 9202 6356 9212
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4844 7634 4900 7644
rect 4060 7410 4116 7420
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 3724 6290 3780 6300
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 2044 6066 2100 6076
rect 2492 6066 2548 6076
rect 1932 5852 2100 5908
rect 1708 5236 1764 5740
rect 1708 5170 1764 5180
rect 1260 4722 1316 4732
rect 1708 5010 1764 5022
rect 1708 4958 1710 5010
rect 1762 4958 1764 5010
rect 1708 4900 1764 4958
rect 2044 5010 2100 5852
rect 2492 5796 2548 5806
rect 2492 5702 2548 5740
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 2044 4958 2046 5010
rect 2098 4958 2100 5010
rect 2044 4946 2100 4958
rect 2492 5122 2548 5134
rect 2492 5070 2494 5122
rect 2546 5070 2548 5122
rect 1708 4340 1764 4844
rect 2492 4900 2548 5070
rect 2492 4834 2548 4844
rect 1708 4274 1764 4284
rect 2044 4788 2100 4798
rect 1708 3444 1764 3482
rect 1708 3378 1764 3388
rect 2044 3442 2100 4732
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 2044 3390 2046 3442
rect 2098 3390 2100 3442
rect 2044 3378 2100 3390
rect 2492 3444 2548 3482
rect 2492 3378 2548 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
<< via2 >>
rect 1148 35980 1204 36036
rect 2380 37938 2436 37940
rect 2380 37886 2382 37938
rect 2382 37886 2434 37938
rect 2434 37886 2436 37938
rect 2380 37884 2436 37886
rect 2268 37772 2324 37828
rect 2380 37436 2436 37492
rect 2716 37324 2772 37380
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4284 38108 4340 38164
rect 5964 38050 6020 38052
rect 5964 37998 5966 38050
rect 5966 37998 6018 38050
rect 6018 37998 6020 38050
rect 5964 37996 6020 37998
rect 3948 37826 4004 37828
rect 3948 37774 3950 37826
rect 3950 37774 4002 37826
rect 4002 37774 4004 37826
rect 3948 37772 4004 37774
rect 3388 37324 3444 37380
rect 2044 36876 2100 36932
rect 1596 35868 1652 35924
rect 1596 33852 1652 33908
rect 1820 35756 1876 35812
rect 3164 37212 3220 37268
rect 2716 37154 2772 37156
rect 2716 37102 2718 37154
rect 2718 37102 2770 37154
rect 2770 37102 2772 37154
rect 2716 37100 2772 37102
rect 2940 36876 2996 36932
rect 2604 36482 2660 36484
rect 2604 36430 2606 36482
rect 2606 36430 2658 36482
rect 2658 36430 2660 36482
rect 2604 36428 2660 36430
rect 3836 36876 3892 36932
rect 3500 36652 3556 36708
rect 4060 36594 4116 36596
rect 4060 36542 4062 36594
rect 4062 36542 4114 36594
rect 4114 36542 4116 36594
rect 4060 36540 4116 36542
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4284 36428 4340 36484
rect 2156 36092 2212 36148
rect 4844 36652 4900 36708
rect 5404 37266 5460 37268
rect 5404 37214 5406 37266
rect 5406 37214 5458 37266
rect 5458 37214 5460 37266
rect 5404 37212 5460 37214
rect 5852 37212 5908 37268
rect 5292 36428 5348 36484
rect 4956 36316 5012 36372
rect 1932 34412 1988 34468
rect 4396 35810 4452 35812
rect 4396 35758 4398 35810
rect 4398 35758 4450 35810
rect 4450 35758 4452 35810
rect 4396 35756 4452 35758
rect 4956 35756 5012 35812
rect 3948 35644 4004 35700
rect 2604 35532 2660 35588
rect 3612 35586 3668 35588
rect 3612 35534 3614 35586
rect 3614 35534 3666 35586
rect 3666 35534 3668 35586
rect 3612 35532 3668 35534
rect 2380 34860 2436 34916
rect 2828 34748 2884 34804
rect 2044 34130 2100 34132
rect 2044 34078 2046 34130
rect 2046 34078 2098 34130
rect 2098 34078 2100 34130
rect 2044 34076 2100 34078
rect 2604 34690 2660 34692
rect 2604 34638 2606 34690
rect 2606 34638 2658 34690
rect 2658 34638 2660 34690
rect 2604 34636 2660 34638
rect 1708 30994 1764 30996
rect 1708 30942 1710 30994
rect 1710 30942 1762 30994
rect 1762 30942 1764 30994
rect 1708 30940 1764 30942
rect 1708 29820 1764 29876
rect 2268 34412 2324 34468
rect 2156 33292 2212 33348
rect 2268 34242 2324 34244
rect 2268 34190 2270 34242
rect 2270 34190 2322 34242
rect 2322 34190 2324 34242
rect 2268 34188 2324 34190
rect 2268 33068 2324 33124
rect 2492 33234 2548 33236
rect 2492 33182 2494 33234
rect 2494 33182 2546 33234
rect 2546 33182 2548 33234
rect 2492 33180 2548 33182
rect 2492 32674 2548 32676
rect 2492 32622 2494 32674
rect 2494 32622 2546 32674
rect 2546 32622 2548 32674
rect 2492 32620 2548 32622
rect 2940 34412 2996 34468
rect 3836 34690 3892 34692
rect 3836 34638 3838 34690
rect 3838 34638 3890 34690
rect 3890 34638 3892 34690
rect 3836 34636 3892 34638
rect 3388 34188 3444 34244
rect 2828 33964 2884 34020
rect 3052 34076 3108 34132
rect 2828 33068 2884 33124
rect 3164 33964 3220 34020
rect 2268 32002 2324 32004
rect 2268 31950 2270 32002
rect 2270 31950 2322 32002
rect 2322 31950 2324 32002
rect 2268 31948 2324 31950
rect 2604 31554 2660 31556
rect 2604 31502 2606 31554
rect 2606 31502 2658 31554
rect 2658 31502 2660 31554
rect 2604 31500 2660 31502
rect 2492 31164 2548 31220
rect 2044 31106 2100 31108
rect 2044 31054 2046 31106
rect 2046 31054 2098 31106
rect 2098 31054 2100 31106
rect 2044 31052 2100 31054
rect 1932 30940 1988 30996
rect 1932 30268 1988 30324
rect 2044 30380 2100 30436
rect 2604 29820 2660 29876
rect 1372 29484 1428 29540
rect 1148 13804 1204 13860
rect 1260 20748 1316 20804
rect 2044 29538 2100 29540
rect 2044 29486 2046 29538
rect 2046 29486 2098 29538
rect 2098 29486 2100 29538
rect 2044 29484 2100 29486
rect 2380 29426 2436 29428
rect 2380 29374 2382 29426
rect 2382 29374 2434 29426
rect 2434 29374 2436 29426
rect 2380 29372 2436 29374
rect 1820 28476 1876 28532
rect 1708 26796 1764 26852
rect 2268 26460 2324 26516
rect 2156 25564 2212 25620
rect 2380 25788 2436 25844
rect 2044 25282 2100 25284
rect 2044 25230 2046 25282
rect 2046 25230 2098 25282
rect 2098 25230 2100 25282
rect 2044 25228 2100 25230
rect 1820 24892 1876 24948
rect 1708 23996 1764 24052
rect 1596 21308 1652 21364
rect 1932 23154 1988 23156
rect 1932 23102 1934 23154
rect 1934 23102 1986 23154
rect 1986 23102 1988 23154
rect 1932 23100 1988 23102
rect 2604 27916 2660 27972
rect 3500 33458 3556 33460
rect 3500 33406 3502 33458
rect 3502 33406 3554 33458
rect 3554 33406 3556 33458
rect 3500 33404 3556 33406
rect 3612 32620 3668 32676
rect 3276 31948 3332 32004
rect 3500 31890 3556 31892
rect 3500 31838 3502 31890
rect 3502 31838 3554 31890
rect 3554 31838 3556 31890
rect 3500 31836 3556 31838
rect 3388 31724 3444 31780
rect 3724 31948 3780 32004
rect 5740 36482 5796 36484
rect 5740 36430 5742 36482
rect 5742 36430 5794 36482
rect 5794 36430 5796 36482
rect 5740 36428 5796 36430
rect 5964 36540 6020 36596
rect 6076 35586 6132 35588
rect 6076 35534 6078 35586
rect 6078 35534 6130 35586
rect 6130 35534 6132 35586
rect 6076 35532 6132 35534
rect 5068 35420 5124 35476
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 6412 37548 6468 37604
rect 7756 38162 7812 38164
rect 7756 38110 7758 38162
rect 7758 38110 7810 38162
rect 7810 38110 7812 38162
rect 7756 38108 7812 38110
rect 7308 38050 7364 38052
rect 7308 37998 7310 38050
rect 7310 37998 7362 38050
rect 7362 37998 7364 38050
rect 7308 37996 7364 37998
rect 6524 37436 6580 37492
rect 6300 37100 6356 37156
rect 6748 37378 6804 37380
rect 6748 37326 6750 37378
rect 6750 37326 6802 37378
rect 6802 37326 6804 37378
rect 6748 37324 6804 37326
rect 6860 37154 6916 37156
rect 6860 37102 6862 37154
rect 6862 37102 6914 37154
rect 6914 37102 6916 37154
rect 6860 37100 6916 37102
rect 6524 36988 6580 37044
rect 6412 36540 6468 36596
rect 8204 37938 8260 37940
rect 8204 37886 8206 37938
rect 8206 37886 8258 37938
rect 8258 37886 8260 37938
rect 8204 37884 8260 37886
rect 9548 37884 9604 37940
rect 9548 37548 9604 37604
rect 8652 37436 8708 37492
rect 7308 36540 7364 36596
rect 7756 36988 7812 37044
rect 6972 36482 7028 36484
rect 6972 36430 6974 36482
rect 6974 36430 7026 36482
rect 7026 36430 7028 36482
rect 6972 36428 7028 36430
rect 6412 36258 6468 36260
rect 6412 36206 6414 36258
rect 6414 36206 6466 36258
rect 6466 36206 6468 36258
rect 6412 36204 6468 36206
rect 6860 35922 6916 35924
rect 6860 35870 6862 35922
rect 6862 35870 6914 35922
rect 6914 35870 6916 35922
rect 6860 35868 6916 35870
rect 7308 35810 7364 35812
rect 7308 35758 7310 35810
rect 7310 35758 7362 35810
rect 7362 35758 7364 35810
rect 7308 35756 7364 35758
rect 6412 35420 6468 35476
rect 7644 35308 7700 35364
rect 4844 34802 4900 34804
rect 4844 34750 4846 34802
rect 4846 34750 4898 34802
rect 4898 34750 4900 34802
rect 4844 34748 4900 34750
rect 4732 34636 4788 34692
rect 4284 33852 4340 33908
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4284 32956 4340 33012
rect 4396 32732 4452 32788
rect 6188 34412 6244 34468
rect 5628 33964 5684 34020
rect 6300 34076 6356 34132
rect 5852 33516 5908 33572
rect 4956 33292 5012 33348
rect 5628 33346 5684 33348
rect 5628 33294 5630 33346
rect 5630 33294 5682 33346
rect 5682 33294 5684 33346
rect 5628 33292 5684 33294
rect 6300 33180 6356 33236
rect 5180 33122 5236 33124
rect 5180 33070 5182 33122
rect 5182 33070 5234 33122
rect 5234 33070 5236 33122
rect 5180 33068 5236 33070
rect 3948 32060 4004 32116
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4732 31948 4788 32004
rect 3836 31612 3892 31668
rect 3052 30322 3108 30324
rect 3052 30270 3054 30322
rect 3054 30270 3106 30322
rect 3106 30270 3108 30322
rect 3052 30268 3108 30270
rect 2828 29986 2884 29988
rect 2828 29934 2830 29986
rect 2830 29934 2882 29986
rect 2882 29934 2884 29986
rect 2828 29932 2884 29934
rect 3052 29820 3108 29876
rect 2828 28476 2884 28532
rect 4844 31724 4900 31780
rect 3612 31052 3668 31108
rect 3612 29932 3668 29988
rect 3500 29260 3556 29316
rect 3612 29372 3668 29428
rect 3500 29036 3556 29092
rect 3276 27916 3332 27972
rect 3164 27074 3220 27076
rect 3164 27022 3166 27074
rect 3166 27022 3218 27074
rect 3218 27022 3220 27074
rect 3164 27020 3220 27022
rect 2604 26460 2660 26516
rect 2604 26290 2660 26292
rect 2604 26238 2606 26290
rect 2606 26238 2658 26290
rect 2658 26238 2660 26290
rect 2604 26236 2660 26238
rect 2940 24050 2996 24052
rect 2940 23998 2942 24050
rect 2942 23998 2994 24050
rect 2994 23998 2996 24050
rect 2940 23996 2996 23998
rect 2716 23324 2772 23380
rect 1820 22370 1876 22372
rect 1820 22318 1822 22370
rect 1822 22318 1874 22370
rect 1874 22318 1876 22370
rect 1820 22316 1876 22318
rect 2380 22316 2436 22372
rect 2044 22146 2100 22148
rect 2044 22094 2046 22146
rect 2046 22094 2098 22146
rect 2098 22094 2100 22146
rect 2044 22092 2100 22094
rect 2044 21698 2100 21700
rect 2044 21646 2046 21698
rect 2046 21646 2098 21698
rect 2098 21646 2100 21698
rect 2044 21644 2100 21646
rect 2268 21420 2324 21476
rect 1708 20690 1764 20692
rect 1708 20638 1710 20690
rect 1710 20638 1762 20690
rect 1762 20638 1764 20690
rect 1708 20636 1764 20638
rect 1708 20412 1764 20468
rect 1708 19740 1764 19796
rect 1708 19122 1764 19124
rect 1708 19070 1710 19122
rect 1710 19070 1762 19122
rect 1762 19070 1764 19122
rect 1708 19068 1764 19070
rect 1708 18620 1764 18676
rect 1708 17724 1764 17780
rect 2940 22370 2996 22372
rect 2940 22318 2942 22370
rect 2942 22318 2994 22370
rect 2994 22318 2996 22370
rect 2940 22316 2996 22318
rect 3276 26460 3332 26516
rect 3388 26124 3444 26180
rect 3388 25228 3444 25284
rect 3164 25004 3220 25060
rect 2828 21532 2884 21588
rect 2716 21420 2772 21476
rect 3612 24444 3668 24500
rect 3948 30380 4004 30436
rect 4732 30828 4788 30884
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4284 30380 4340 30436
rect 4508 30268 4564 30324
rect 3836 29596 3892 29652
rect 3948 29372 4004 29428
rect 3836 28588 3892 28644
rect 3836 27020 3892 27076
rect 3388 22540 3444 22596
rect 3500 24108 3556 24164
rect 2380 20860 2436 20916
rect 3164 21532 3220 21588
rect 2380 20018 2436 20020
rect 2380 19966 2382 20018
rect 2382 19966 2434 20018
rect 2434 19966 2436 20018
rect 2380 19964 2436 19966
rect 2940 20860 2996 20916
rect 3052 20802 3108 20804
rect 3052 20750 3054 20802
rect 3054 20750 3106 20802
rect 3106 20750 3108 20802
rect 3052 20748 3108 20750
rect 3388 21586 3444 21588
rect 3388 21534 3390 21586
rect 3390 21534 3442 21586
rect 3442 21534 3444 21586
rect 3388 21532 3444 21534
rect 3276 20860 3332 20916
rect 4844 29932 4900 29988
rect 4172 29260 4228 29316
rect 4396 29426 4452 29428
rect 4396 29374 4398 29426
rect 4398 29374 4450 29426
rect 4450 29374 4452 29426
rect 4396 29372 4452 29374
rect 4284 29036 4340 29092
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4284 28588 4340 28644
rect 4844 27916 4900 27972
rect 5292 32060 5348 32116
rect 5180 31948 5236 32004
rect 5628 31500 5684 31556
rect 5964 31388 6020 31444
rect 6188 31612 6244 31668
rect 4956 29538 5012 29540
rect 4956 29486 4958 29538
rect 4958 29486 5010 29538
rect 5010 29486 5012 29538
rect 4956 29484 5012 29486
rect 6076 30268 6132 30324
rect 5180 30156 5236 30212
rect 8204 36428 8260 36484
rect 8092 36258 8148 36260
rect 8092 36206 8094 36258
rect 8094 36206 8146 36258
rect 8146 36206 8148 36258
rect 8092 36204 8148 36206
rect 8204 35420 8260 35476
rect 6524 34802 6580 34804
rect 6524 34750 6526 34802
rect 6526 34750 6578 34802
rect 6578 34750 6580 34802
rect 6524 34748 6580 34750
rect 8204 34412 8260 34468
rect 7868 34354 7924 34356
rect 7868 34302 7870 34354
rect 7870 34302 7922 34354
rect 7922 34302 7924 34354
rect 7868 34300 7924 34302
rect 6412 32172 6468 32228
rect 6748 33516 6804 33572
rect 7868 33852 7924 33908
rect 6860 32956 6916 33012
rect 6524 31836 6580 31892
rect 6636 31724 6692 31780
rect 7084 33458 7140 33460
rect 7084 33406 7086 33458
rect 7086 33406 7138 33458
rect 7138 33406 7140 33458
rect 7084 33404 7140 33406
rect 6524 30828 6580 30884
rect 6412 30322 6468 30324
rect 6412 30270 6414 30322
rect 6414 30270 6466 30322
rect 6466 30270 6468 30322
rect 6412 30268 6468 30270
rect 6636 30210 6692 30212
rect 6636 30158 6638 30210
rect 6638 30158 6690 30210
rect 6690 30158 6692 30210
rect 6636 30156 6692 30158
rect 5068 28754 5124 28756
rect 5068 28702 5070 28754
rect 5070 28702 5122 28754
rect 5122 28702 5124 28754
rect 5068 28700 5124 28702
rect 5180 29484 5236 29540
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4956 27186 5012 27188
rect 4956 27134 4958 27186
rect 4958 27134 5010 27186
rect 5010 27134 5012 27186
rect 4956 27132 5012 27134
rect 5068 27074 5124 27076
rect 5068 27022 5070 27074
rect 5070 27022 5122 27074
rect 5122 27022 5124 27074
rect 5068 27020 5124 27022
rect 4060 26178 4116 26180
rect 4060 26126 4062 26178
rect 4062 26126 4114 26178
rect 4114 26126 4116 26178
rect 4060 26124 4116 26126
rect 4060 24946 4116 24948
rect 4060 24894 4062 24946
rect 4062 24894 4114 24946
rect 4114 24894 4116 24946
rect 4060 24892 4116 24894
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4508 25564 4564 25620
rect 4620 25452 4676 25508
rect 4172 24722 4228 24724
rect 4172 24670 4174 24722
rect 4174 24670 4226 24722
rect 4226 24670 4228 24722
rect 4172 24668 4228 24670
rect 4508 25394 4564 25396
rect 4508 25342 4510 25394
rect 4510 25342 4562 25394
rect 4562 25342 4564 25394
rect 4508 25340 4564 25342
rect 3948 24108 4004 24164
rect 4060 24498 4116 24500
rect 4060 24446 4062 24498
rect 4062 24446 4114 24498
rect 4114 24446 4116 24498
rect 4060 24444 4116 24446
rect 3948 23938 4004 23940
rect 3948 23886 3950 23938
rect 3950 23886 4002 23938
rect 4002 23886 4004 23938
rect 3948 23884 4004 23886
rect 5068 25564 5124 25620
rect 4956 24892 5012 24948
rect 4620 24444 4676 24500
rect 5068 24780 5124 24836
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4172 23826 4228 23828
rect 4172 23774 4174 23826
rect 4174 23774 4226 23826
rect 4226 23774 4228 23826
rect 4172 23772 4228 23774
rect 4620 23826 4676 23828
rect 4620 23774 4622 23826
rect 4622 23774 4674 23826
rect 4674 23774 4676 23826
rect 4620 23772 4676 23774
rect 4732 23660 4788 23716
rect 4844 23548 4900 23604
rect 4956 23100 5012 23156
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4172 22482 4228 22484
rect 4172 22430 4174 22482
rect 4174 22430 4226 22482
rect 4226 22430 4228 22482
rect 4172 22428 4228 22430
rect 5068 22764 5124 22820
rect 4284 22370 4340 22372
rect 4284 22318 4286 22370
rect 4286 22318 4338 22370
rect 4338 22318 4340 22370
rect 4284 22316 4340 22318
rect 3724 22258 3780 22260
rect 3724 22206 3726 22258
rect 3726 22206 3778 22258
rect 3778 22206 3780 22258
rect 3724 22204 3780 22206
rect 4172 22146 4228 22148
rect 4172 22094 4174 22146
rect 4174 22094 4226 22146
rect 4226 22094 4228 22146
rect 4172 22092 4228 22094
rect 3948 21980 4004 22036
rect 3836 21810 3892 21812
rect 3836 21758 3838 21810
rect 3838 21758 3890 21810
rect 3890 21758 3892 21810
rect 3836 21756 3892 21758
rect 4844 22146 4900 22148
rect 4844 22094 4846 22146
rect 4846 22094 4898 22146
rect 4898 22094 4900 22146
rect 4844 22092 4900 22094
rect 4732 21756 4788 21812
rect 4284 21532 4340 21588
rect 3836 20972 3892 21028
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3164 20524 3220 20580
rect 2828 20076 2884 20132
rect 3052 19852 3108 19908
rect 2380 19516 2436 19572
rect 2716 19180 2772 19236
rect 2268 18732 2324 18788
rect 2716 18844 2772 18900
rect 2380 18620 2436 18676
rect 2380 17948 2436 18004
rect 1932 17666 1988 17668
rect 1932 17614 1934 17666
rect 1934 17614 1986 17666
rect 1986 17614 1988 17666
rect 1932 17612 1988 17614
rect 1932 17164 1988 17220
rect 1372 16044 1428 16100
rect 1708 16828 1764 16884
rect 1484 15932 1540 15988
rect 1708 15708 1764 15764
rect 1484 14364 1540 14420
rect 2268 16716 2324 16772
rect 2492 16716 2548 16772
rect 2492 15708 2548 15764
rect 2380 15314 2436 15316
rect 2380 15262 2382 15314
rect 2382 15262 2434 15314
rect 2434 15262 2436 15314
rect 2380 15260 2436 15262
rect 2492 14364 2548 14420
rect 1708 14140 1764 14196
rect 1708 13580 1764 13636
rect 1708 13244 1764 13300
rect 1708 12348 1764 12404
rect 1708 12012 1764 12068
rect 1708 11452 1764 11508
rect 1708 11116 1764 11172
rect 1708 10556 1764 10612
rect 2044 13970 2100 13972
rect 2044 13918 2046 13970
rect 2046 13918 2098 13970
rect 2098 13918 2100 13970
rect 2044 13916 2100 13918
rect 3724 20524 3780 20580
rect 3612 19964 3668 20020
rect 3052 18620 3108 18676
rect 2940 18562 2996 18564
rect 2940 18510 2942 18562
rect 2942 18510 2994 18562
rect 2994 18510 2996 18562
rect 2940 18508 2996 18510
rect 3276 17666 3332 17668
rect 3276 17614 3278 17666
rect 3278 17614 3330 17666
rect 3330 17614 3332 17666
rect 3276 17612 3332 17614
rect 3164 16716 3220 16772
rect 3276 16268 3332 16324
rect 3164 15932 3220 15988
rect 5628 28642 5684 28644
rect 5628 28590 5630 28642
rect 5630 28590 5682 28642
rect 5682 28590 5684 28642
rect 5628 28588 5684 28590
rect 5740 28530 5796 28532
rect 5740 28478 5742 28530
rect 5742 28478 5794 28530
rect 5794 28478 5796 28530
rect 5740 28476 5796 28478
rect 5740 27020 5796 27076
rect 6188 29596 6244 29652
rect 5292 25228 5348 25284
rect 6860 30994 6916 30996
rect 6860 30942 6862 30994
rect 6862 30942 6914 30994
rect 6914 30942 6916 30994
rect 6860 30940 6916 30942
rect 6972 30380 7028 30436
rect 7084 31666 7140 31668
rect 7084 31614 7086 31666
rect 7086 31614 7138 31666
rect 7138 31614 7140 31666
rect 7084 31612 7140 31614
rect 6972 29596 7028 29652
rect 6412 28476 6468 28532
rect 6748 28700 6804 28756
rect 6524 27970 6580 27972
rect 6524 27918 6526 27970
rect 6526 27918 6578 27970
rect 6578 27918 6580 27970
rect 6524 27916 6580 27918
rect 5516 25340 5572 25396
rect 5852 25618 5908 25620
rect 5852 25566 5854 25618
rect 5854 25566 5906 25618
rect 5906 25566 5908 25618
rect 5852 25564 5908 25566
rect 5628 24892 5684 24948
rect 5964 26124 6020 26180
rect 5852 24668 5908 24724
rect 5628 23772 5684 23828
rect 6636 26572 6692 26628
rect 6188 25506 6244 25508
rect 6188 25454 6190 25506
rect 6190 25454 6242 25506
rect 6242 25454 6244 25506
rect 6188 25452 6244 25454
rect 6524 25340 6580 25396
rect 6636 25228 6692 25284
rect 6076 24780 6132 24836
rect 6412 24834 6468 24836
rect 6412 24782 6414 24834
rect 6414 24782 6466 24834
rect 6466 24782 6468 24834
rect 6412 24780 6468 24782
rect 6636 23714 6692 23716
rect 6636 23662 6638 23714
rect 6638 23662 6690 23714
rect 6690 23662 6692 23714
rect 6636 23660 6692 23662
rect 6972 23660 7028 23716
rect 5964 23436 6020 23492
rect 6860 23378 6916 23380
rect 6860 23326 6862 23378
rect 6862 23326 6914 23378
rect 6914 23326 6916 23378
rect 6860 23324 6916 23326
rect 6412 23212 6468 23268
rect 6076 22764 6132 22820
rect 5740 22316 5796 22372
rect 6412 22316 6468 22372
rect 5740 22092 5796 22148
rect 5180 21084 5236 21140
rect 5516 21980 5572 22036
rect 5180 20690 5236 20692
rect 5180 20638 5182 20690
rect 5182 20638 5234 20690
rect 5234 20638 5236 20690
rect 5180 20636 5236 20638
rect 5852 21644 5908 21700
rect 6188 21756 6244 21812
rect 5852 20636 5908 20692
rect 3836 18956 3892 19012
rect 4396 19906 4452 19908
rect 4396 19854 4398 19906
rect 4398 19854 4450 19906
rect 4450 19854 4452 19906
rect 4396 19852 4452 19854
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 5404 20130 5460 20132
rect 5404 20078 5406 20130
rect 5406 20078 5458 20130
rect 5458 20078 5460 20130
rect 5404 20076 5460 20078
rect 4956 20018 5012 20020
rect 4956 19966 4958 20018
rect 4958 19966 5010 20018
rect 5010 19966 5012 20018
rect 4956 19964 5012 19966
rect 4172 18620 4228 18676
rect 3948 18508 4004 18564
rect 3836 17612 3892 17668
rect 3836 17106 3892 17108
rect 3836 17054 3838 17106
rect 3838 17054 3890 17106
rect 3890 17054 3892 17106
rect 3836 17052 3892 17054
rect 4060 17106 4116 17108
rect 4060 17054 4062 17106
rect 4062 17054 4114 17106
rect 4114 17054 4116 17106
rect 4060 17052 4116 17054
rect 3948 16940 4004 16996
rect 3724 16156 3780 16212
rect 3836 16828 3892 16884
rect 3612 16098 3668 16100
rect 3612 16046 3614 16098
rect 3614 16046 3666 16098
rect 3666 16046 3668 16098
rect 3612 16044 3668 16046
rect 3612 15708 3668 15764
rect 4844 19010 4900 19012
rect 4844 18958 4846 19010
rect 4846 18958 4898 19010
rect 4898 18958 4900 19010
rect 4844 18956 4900 18958
rect 4508 18562 4564 18564
rect 4508 18510 4510 18562
rect 4510 18510 4562 18562
rect 4562 18510 4564 18562
rect 4508 18508 4564 18510
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4620 17778 4676 17780
rect 4620 17726 4622 17778
rect 4622 17726 4674 17778
rect 4674 17726 4676 17778
rect 4620 17724 4676 17726
rect 4284 17052 4340 17108
rect 4732 17106 4788 17108
rect 4732 17054 4734 17106
rect 4734 17054 4786 17106
rect 4786 17054 4788 17106
rect 4732 17052 4788 17054
rect 5292 19180 5348 19236
rect 5068 18562 5124 18564
rect 5068 18510 5070 18562
rect 5070 18510 5122 18562
rect 5122 18510 5124 18562
rect 5068 18508 5124 18510
rect 6188 20188 6244 20244
rect 5628 20018 5684 20020
rect 5628 19966 5630 20018
rect 5630 19966 5682 20018
rect 5682 19966 5684 20018
rect 5628 19964 5684 19966
rect 5740 19122 5796 19124
rect 5740 19070 5742 19122
rect 5742 19070 5794 19122
rect 5794 19070 5796 19122
rect 5740 19068 5796 19070
rect 5852 18508 5908 18564
rect 5292 17836 5348 17892
rect 4508 16716 4564 16772
rect 4844 16770 4900 16772
rect 4844 16718 4846 16770
rect 4846 16718 4898 16770
rect 4898 16718 4900 16770
rect 4844 16716 4900 16718
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4172 15708 4228 15764
rect 4060 15596 4116 15652
rect 2828 14588 2884 14644
rect 2940 14924 2996 14980
rect 3052 14812 3108 14868
rect 2940 13634 2996 13636
rect 2940 13582 2942 13634
rect 2942 13582 2994 13634
rect 2994 13582 2996 13634
rect 2940 13580 2996 13582
rect 2044 13356 2100 13412
rect 3836 14754 3892 14756
rect 3836 14702 3838 14754
rect 3838 14702 3890 14754
rect 3890 14702 3892 14754
rect 3836 14700 3892 14702
rect 3388 14140 3444 14196
rect 3836 13916 3892 13972
rect 2492 12348 2548 12404
rect 2492 12066 2548 12068
rect 2492 12014 2494 12066
rect 2494 12014 2546 12066
rect 2546 12014 2548 12066
rect 2492 12012 2548 12014
rect 2492 11170 2548 11172
rect 2492 11118 2494 11170
rect 2494 11118 2546 11170
rect 2546 11118 2548 11170
rect 2492 11116 2548 11118
rect 1932 9660 1988 9716
rect 2492 9714 2548 9716
rect 2492 9662 2494 9714
rect 2494 9662 2546 9714
rect 2546 9662 2548 9714
rect 2492 9660 2548 9662
rect 1708 8764 1764 8820
rect 1708 7868 1764 7924
rect 1708 6972 1764 7028
rect 1708 6076 1764 6132
rect 2044 9266 2100 9268
rect 2044 9214 2046 9266
rect 2046 9214 2098 9266
rect 2098 9214 2100 9266
rect 2044 9212 2100 9214
rect 2492 8764 2548 8820
rect 4060 11340 4116 11396
rect 4620 15932 4676 15988
rect 4620 15260 4676 15316
rect 4844 16156 4900 16212
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 2044 8146 2100 8148
rect 2044 8094 2046 8146
rect 2046 8094 2098 8146
rect 2098 8094 2100 8146
rect 2044 8092 2100 8094
rect 2492 7868 2548 7924
rect 2044 7698 2100 7700
rect 2044 7646 2046 7698
rect 2046 7646 2098 7698
rect 2098 7646 2100 7698
rect 2044 7644 2100 7646
rect 2044 7420 2100 7476
rect 2492 6972 2548 7028
rect 2156 6300 2212 6356
rect 5068 16268 5124 16324
rect 5180 16044 5236 16100
rect 4956 15148 5012 15204
rect 5404 17276 5460 17332
rect 5628 16268 5684 16324
rect 5852 16098 5908 16100
rect 5852 16046 5854 16098
rect 5854 16046 5906 16098
rect 5906 16046 5908 16098
rect 5852 16044 5908 16046
rect 6076 15820 6132 15876
rect 6972 22428 7028 22484
rect 6412 20972 6468 21028
rect 6412 19906 6468 19908
rect 6412 19854 6414 19906
rect 6414 19854 6466 19906
rect 6466 19854 6468 19906
rect 6412 19852 6468 19854
rect 6636 21420 6692 21476
rect 6972 19292 7028 19348
rect 7756 32956 7812 33012
rect 7868 31836 7924 31892
rect 7420 31388 7476 31444
rect 7868 31500 7924 31556
rect 7532 30828 7588 30884
rect 7308 30268 7364 30324
rect 7196 27746 7252 27748
rect 7196 27694 7198 27746
rect 7198 27694 7250 27746
rect 7250 27694 7252 27746
rect 7196 27692 7252 27694
rect 8428 34130 8484 34132
rect 8428 34078 8430 34130
rect 8430 34078 8482 34130
rect 8482 34078 8484 34130
rect 8428 34076 8484 34078
rect 8652 35308 8708 35364
rect 8652 34972 8708 35028
rect 8764 34914 8820 34916
rect 8764 34862 8766 34914
rect 8766 34862 8818 34914
rect 8818 34862 8820 34914
rect 8764 34860 8820 34862
rect 8316 32284 8372 32340
rect 8204 30268 8260 30324
rect 8316 31388 8372 31444
rect 7868 30156 7924 30212
rect 7868 29708 7924 29764
rect 7644 29372 7700 29428
rect 7756 29314 7812 29316
rect 7756 29262 7758 29314
rect 7758 29262 7810 29314
rect 7810 29262 7812 29314
rect 7756 29260 7812 29262
rect 7756 28700 7812 28756
rect 8092 28754 8148 28756
rect 8092 28702 8094 28754
rect 8094 28702 8146 28754
rect 8146 28702 8148 28754
rect 8092 28700 8148 28702
rect 7196 26348 7252 26404
rect 7308 26572 7364 26628
rect 7308 25452 7364 25508
rect 7980 28476 8036 28532
rect 8092 27132 8148 27188
rect 8540 31500 8596 31556
rect 8428 30268 8484 30324
rect 8876 31778 8932 31780
rect 8876 31726 8878 31778
rect 8878 31726 8930 31778
rect 8930 31726 8932 31778
rect 8876 31724 8932 31726
rect 8652 30156 8708 30212
rect 8988 30434 9044 30436
rect 8988 30382 8990 30434
rect 8990 30382 9042 30434
rect 9042 30382 9044 30434
rect 8988 30380 9044 30382
rect 9100 30210 9156 30212
rect 9100 30158 9102 30210
rect 9102 30158 9154 30210
rect 9154 30158 9156 30210
rect 9100 30156 9156 30158
rect 8764 29650 8820 29652
rect 8764 29598 8766 29650
rect 8766 29598 8818 29650
rect 8818 29598 8820 29650
rect 8764 29596 8820 29598
rect 8316 29260 8372 29316
rect 8428 28364 8484 28420
rect 8652 29426 8708 29428
rect 8652 29374 8654 29426
rect 8654 29374 8706 29426
rect 8706 29374 8708 29426
rect 8652 29372 8708 29374
rect 8876 29260 8932 29316
rect 9548 33180 9604 33236
rect 11004 38162 11060 38164
rect 11004 38110 11006 38162
rect 11006 38110 11058 38162
rect 11058 38110 11060 38162
rect 11004 38108 11060 38110
rect 9996 37100 10052 37156
rect 10220 37212 10276 37268
rect 9772 34130 9828 34132
rect 9772 34078 9774 34130
rect 9774 34078 9826 34130
rect 9826 34078 9828 34130
rect 9772 34076 9828 34078
rect 11004 36988 11060 37044
rect 11004 35698 11060 35700
rect 11004 35646 11006 35698
rect 11006 35646 11058 35698
rect 11058 35646 11060 35698
rect 11004 35644 11060 35646
rect 10780 34972 10836 35028
rect 10108 33292 10164 33348
rect 10332 33234 10388 33236
rect 10332 33182 10334 33234
rect 10334 33182 10386 33234
rect 10386 33182 10388 33234
rect 10332 33180 10388 33182
rect 10780 33068 10836 33124
rect 10108 32284 10164 32340
rect 9996 32172 10052 32228
rect 9436 30044 9492 30100
rect 9548 31612 9604 31668
rect 9548 29986 9604 29988
rect 9548 29934 9550 29986
rect 9550 29934 9602 29986
rect 9602 29934 9604 29986
rect 9548 29932 9604 29934
rect 9996 31388 10052 31444
rect 10220 30994 10276 30996
rect 10220 30942 10222 30994
rect 10222 30942 10274 30994
rect 10274 30942 10276 30994
rect 10220 30940 10276 30942
rect 9884 30828 9940 30884
rect 10220 30716 10276 30772
rect 9996 30322 10052 30324
rect 9996 30270 9998 30322
rect 9998 30270 10050 30322
rect 10050 30270 10052 30322
rect 9996 30268 10052 30270
rect 9772 29484 9828 29540
rect 9884 30044 9940 30100
rect 8428 26572 8484 26628
rect 8092 26178 8148 26180
rect 8092 26126 8094 26178
rect 8094 26126 8146 26178
rect 8146 26126 8148 26178
rect 8092 26124 8148 26126
rect 7420 25228 7476 25284
rect 7756 25282 7812 25284
rect 7756 25230 7758 25282
rect 7758 25230 7810 25282
rect 7810 25230 7812 25282
rect 7756 25228 7812 25230
rect 7532 24668 7588 24724
rect 7420 24556 7476 24612
rect 7644 24444 7700 24500
rect 8092 24332 8148 24388
rect 7868 23996 7924 24052
rect 7756 23154 7812 23156
rect 7756 23102 7758 23154
rect 7758 23102 7810 23154
rect 7810 23102 7812 23154
rect 7756 23100 7812 23102
rect 7420 23042 7476 23044
rect 7420 22990 7422 23042
rect 7422 22990 7474 23042
rect 7474 22990 7476 23042
rect 7420 22988 7476 22990
rect 7532 22652 7588 22708
rect 7308 21868 7364 21924
rect 7196 21532 7252 21588
rect 7308 21084 7364 21140
rect 7756 20860 7812 20916
rect 7644 20188 7700 20244
rect 9548 29426 9604 29428
rect 9548 29374 9550 29426
rect 9550 29374 9602 29426
rect 9602 29374 9604 29426
rect 9548 29372 9604 29374
rect 9996 29426 10052 29428
rect 9996 29374 9998 29426
rect 9998 29374 10050 29426
rect 10050 29374 10052 29426
rect 9996 29372 10052 29374
rect 9772 28588 9828 28644
rect 9660 28364 9716 28420
rect 8988 26684 9044 26740
rect 8204 23324 8260 23380
rect 8316 24668 8372 24724
rect 8428 23938 8484 23940
rect 8428 23886 8430 23938
rect 8430 23886 8482 23938
rect 8482 23886 8484 23938
rect 8428 23884 8484 23886
rect 8092 22876 8148 22932
rect 8652 25004 8708 25060
rect 8876 24946 8932 24948
rect 8876 24894 8878 24946
rect 8878 24894 8930 24946
rect 8930 24894 8932 24946
rect 8876 24892 8932 24894
rect 8764 24610 8820 24612
rect 8764 24558 8766 24610
rect 8766 24558 8818 24610
rect 8818 24558 8820 24610
rect 8764 24556 8820 24558
rect 8876 22988 8932 23044
rect 8540 22764 8596 22820
rect 8876 22764 8932 22820
rect 8316 21756 8372 21812
rect 8652 21586 8708 21588
rect 8652 21534 8654 21586
rect 8654 21534 8706 21586
rect 8706 21534 8708 21586
rect 8652 21532 8708 21534
rect 8204 20802 8260 20804
rect 8204 20750 8206 20802
rect 8206 20750 8258 20802
rect 8258 20750 8260 20802
rect 8204 20748 8260 20750
rect 9436 26684 9492 26740
rect 9100 25228 9156 25284
rect 9212 24220 9268 24276
rect 9324 26460 9380 26516
rect 9100 23154 9156 23156
rect 9100 23102 9102 23154
rect 9102 23102 9154 23154
rect 9154 23102 9156 23154
rect 9100 23100 9156 23102
rect 8988 22316 9044 22372
rect 7196 17106 7252 17108
rect 7196 17054 7198 17106
rect 7198 17054 7250 17106
rect 7250 17054 7252 17106
rect 7196 17052 7252 17054
rect 6860 16828 6916 16884
rect 7532 18226 7588 18228
rect 7532 18174 7534 18226
rect 7534 18174 7586 18226
rect 7586 18174 7588 18226
rect 7532 18172 7588 18174
rect 8092 17724 8148 17780
rect 7868 16994 7924 16996
rect 7868 16942 7870 16994
rect 7870 16942 7922 16994
rect 7922 16942 7924 16994
rect 7868 16940 7924 16942
rect 8316 17276 8372 17332
rect 7756 16882 7812 16884
rect 7756 16830 7758 16882
rect 7758 16830 7810 16882
rect 7810 16830 7812 16882
rect 7756 16828 7812 16830
rect 7420 16716 7476 16772
rect 7868 16380 7924 16436
rect 8204 15986 8260 15988
rect 8204 15934 8206 15986
rect 8206 15934 8258 15986
rect 8258 15934 8260 15986
rect 8204 15932 8260 15934
rect 7980 15708 8036 15764
rect 5292 14700 5348 14756
rect 7196 15314 7252 15316
rect 7196 15262 7198 15314
rect 7198 15262 7250 15314
rect 7250 15262 7252 15314
rect 7196 15260 7252 15262
rect 6972 13692 7028 13748
rect 8876 19852 8932 19908
rect 9100 19852 9156 19908
rect 9548 26124 9604 26180
rect 9996 26402 10052 26404
rect 9996 26350 9998 26402
rect 9998 26350 10050 26402
rect 10050 26350 10052 26402
rect 9996 26348 10052 26350
rect 9996 25228 10052 25284
rect 9884 25004 9940 25060
rect 9436 23324 9492 23380
rect 10332 30492 10388 30548
rect 11228 33180 11284 33236
rect 11004 31948 11060 32004
rect 11116 31890 11172 31892
rect 11116 31838 11118 31890
rect 11118 31838 11170 31890
rect 11170 31838 11172 31890
rect 11116 31836 11172 31838
rect 10444 30156 10500 30212
rect 10556 30380 10612 30436
rect 10444 29372 10500 29428
rect 10332 29036 10388 29092
rect 10332 28252 10388 28308
rect 10668 28700 10724 28756
rect 10668 27244 10724 27300
rect 10668 27020 10724 27076
rect 11228 31612 11284 31668
rect 11452 33628 11508 33684
rect 11452 33234 11508 33236
rect 11452 33182 11454 33234
rect 11454 33182 11506 33234
rect 11506 33182 11508 33234
rect 11452 33180 11508 33182
rect 11452 32338 11508 32340
rect 11452 32286 11454 32338
rect 11454 32286 11506 32338
rect 11506 32286 11508 32338
rect 11452 32284 11508 32286
rect 15932 38220 15988 38276
rect 17164 38274 17220 38276
rect 17164 38222 17166 38274
rect 17166 38222 17218 38274
rect 17218 38222 17220 38274
rect 17164 38220 17220 38222
rect 12572 37996 12628 38052
rect 13132 38108 13188 38164
rect 13692 38108 13748 38164
rect 11788 35644 11844 35700
rect 12348 36764 12404 36820
rect 11900 36652 11956 36708
rect 11788 34748 11844 34804
rect 12012 36428 12068 36484
rect 13468 37938 13524 37940
rect 13468 37886 13470 37938
rect 13470 37886 13522 37938
rect 13522 37886 13524 37938
rect 13468 37884 13524 37886
rect 13468 37436 13524 37492
rect 14252 38050 14308 38052
rect 14252 37998 14254 38050
rect 14254 37998 14306 38050
rect 14306 37998 14308 38050
rect 14252 37996 14308 37998
rect 15036 38050 15092 38052
rect 15036 37998 15038 38050
rect 15038 37998 15090 38050
rect 15090 37998 15092 38050
rect 15036 37996 15092 37998
rect 13356 36988 13412 37044
rect 12796 36540 12852 36596
rect 12908 36482 12964 36484
rect 12908 36430 12910 36482
rect 12910 36430 12962 36482
rect 12962 36430 12964 36482
rect 12908 36428 12964 36430
rect 12572 35698 12628 35700
rect 12572 35646 12574 35698
rect 12574 35646 12626 35698
rect 12626 35646 12628 35698
rect 12572 35644 12628 35646
rect 12236 35420 12292 35476
rect 13692 36428 13748 36484
rect 13804 36316 13860 36372
rect 12908 34802 12964 34804
rect 12908 34750 12910 34802
rect 12910 34750 12962 34802
rect 12962 34750 12964 34802
rect 12908 34748 12964 34750
rect 12460 34018 12516 34020
rect 12460 33966 12462 34018
rect 12462 33966 12514 34018
rect 12514 33966 12516 34018
rect 12460 33964 12516 33966
rect 11788 33346 11844 33348
rect 11788 33294 11790 33346
rect 11790 33294 11842 33346
rect 11842 33294 11844 33346
rect 11788 33292 11844 33294
rect 12460 32844 12516 32900
rect 11676 31554 11732 31556
rect 11676 31502 11678 31554
rect 11678 31502 11730 31554
rect 11730 31502 11732 31554
rect 11676 31500 11732 31502
rect 11116 30716 11172 30772
rect 11004 30268 11060 30324
rect 11340 31106 11396 31108
rect 11340 31054 11342 31106
rect 11342 31054 11394 31106
rect 11394 31054 11396 31106
rect 11340 31052 11396 31054
rect 11340 30380 11396 30436
rect 11452 30940 11508 30996
rect 11228 29314 11284 29316
rect 11228 29262 11230 29314
rect 11230 29262 11282 29314
rect 11282 29262 11284 29314
rect 11228 29260 11284 29262
rect 11340 29148 11396 29204
rect 11004 28700 11060 28756
rect 11228 28252 11284 28308
rect 11452 28642 11508 28644
rect 11452 28590 11454 28642
rect 11454 28590 11506 28642
rect 11506 28590 11508 28642
rect 11452 28588 11508 28590
rect 11676 29148 11732 29204
rect 11564 28476 11620 28532
rect 11340 27244 11396 27300
rect 10780 26012 10836 26068
rect 9996 24220 10052 24276
rect 9884 23436 9940 23492
rect 9660 23100 9716 23156
rect 9772 22876 9828 22932
rect 10220 23548 10276 23604
rect 10220 23212 10276 23268
rect 10108 22092 10164 22148
rect 9660 21532 9716 21588
rect 9772 20578 9828 20580
rect 9772 20526 9774 20578
rect 9774 20526 9826 20578
rect 9826 20526 9828 20578
rect 9772 20524 9828 20526
rect 9548 19234 9604 19236
rect 9548 19182 9550 19234
rect 9550 19182 9602 19234
rect 9602 19182 9604 19234
rect 9548 19180 9604 19182
rect 9324 19010 9380 19012
rect 9324 18958 9326 19010
rect 9326 18958 9378 19010
rect 9378 18958 9380 19010
rect 9324 18956 9380 18958
rect 8764 18732 8820 18788
rect 8876 18620 8932 18676
rect 8764 17666 8820 17668
rect 8764 17614 8766 17666
rect 8766 17614 8818 17666
rect 8818 17614 8820 17666
rect 8764 17612 8820 17614
rect 8652 17106 8708 17108
rect 8652 17054 8654 17106
rect 8654 17054 8706 17106
rect 8706 17054 8708 17106
rect 8652 17052 8708 17054
rect 8540 15874 8596 15876
rect 8540 15822 8542 15874
rect 8542 15822 8594 15874
rect 8594 15822 8596 15874
rect 8540 15820 8596 15822
rect 8652 15708 8708 15764
rect 8092 11564 8148 11620
rect 8988 18450 9044 18452
rect 8988 18398 8990 18450
rect 8990 18398 9042 18450
rect 9042 18398 9044 18450
rect 8988 18396 9044 18398
rect 8988 17106 9044 17108
rect 8988 17054 8990 17106
rect 8990 17054 9042 17106
rect 9042 17054 9044 17106
rect 8988 17052 9044 17054
rect 8988 16828 9044 16884
rect 9548 18620 9604 18676
rect 9548 18450 9604 18452
rect 9548 18398 9550 18450
rect 9550 18398 9602 18450
rect 9602 18398 9604 18450
rect 9548 18396 9604 18398
rect 9772 20188 9828 20244
rect 9884 20076 9940 20132
rect 9772 18396 9828 18452
rect 9660 17052 9716 17108
rect 9436 16380 9492 16436
rect 9212 15986 9268 15988
rect 9212 15934 9214 15986
rect 9214 15934 9266 15986
rect 9266 15934 9268 15986
rect 9212 15932 9268 15934
rect 10220 20412 10276 20468
rect 10444 23436 10500 23492
rect 10668 24722 10724 24724
rect 10668 24670 10670 24722
rect 10670 24670 10722 24722
rect 10722 24670 10724 24722
rect 10668 24668 10724 24670
rect 10780 24108 10836 24164
rect 10668 21980 10724 22036
rect 10780 23324 10836 23380
rect 10444 20524 10500 20580
rect 10556 21532 10612 21588
rect 10108 18450 10164 18452
rect 10108 18398 10110 18450
rect 10110 18398 10162 18450
rect 10162 18398 10164 18450
rect 10108 18396 10164 18398
rect 10444 20300 10500 20356
rect 10332 18956 10388 19012
rect 9996 16770 10052 16772
rect 9996 16718 9998 16770
rect 9998 16718 10050 16770
rect 10050 16718 10052 16770
rect 9996 16716 10052 16718
rect 10108 16940 10164 16996
rect 10556 18674 10612 18676
rect 10556 18622 10558 18674
rect 10558 18622 10610 18674
rect 10610 18622 10612 18674
rect 10556 18620 10612 18622
rect 11004 26124 11060 26180
rect 11004 25676 11060 25732
rect 11228 27020 11284 27076
rect 11228 23884 11284 23940
rect 11564 26290 11620 26292
rect 11564 26238 11566 26290
rect 11566 26238 11618 26290
rect 11618 26238 11620 26290
rect 11564 26236 11620 26238
rect 12012 31554 12068 31556
rect 12012 31502 12014 31554
rect 12014 31502 12066 31554
rect 12066 31502 12068 31554
rect 12012 31500 12068 31502
rect 11900 30098 11956 30100
rect 11900 30046 11902 30098
rect 11902 30046 11954 30098
rect 11954 30046 11956 30098
rect 11900 30044 11956 30046
rect 12348 31836 12404 31892
rect 12348 30940 12404 30996
rect 13580 34018 13636 34020
rect 13580 33966 13582 34018
rect 13582 33966 13634 34018
rect 13634 33966 13636 34018
rect 13580 33964 13636 33966
rect 13580 33068 13636 33124
rect 14140 36652 14196 36708
rect 14252 36876 14308 36932
rect 14028 36482 14084 36484
rect 14028 36430 14030 36482
rect 14030 36430 14082 36482
rect 14082 36430 14084 36482
rect 14028 36428 14084 36430
rect 14252 36092 14308 36148
rect 13916 34076 13972 34132
rect 14252 35026 14308 35028
rect 14252 34974 14254 35026
rect 14254 34974 14306 35026
rect 14306 34974 14308 35026
rect 14252 34972 14308 34974
rect 14140 33906 14196 33908
rect 14140 33854 14142 33906
rect 14142 33854 14194 33906
rect 14194 33854 14196 33906
rect 14140 33852 14196 33854
rect 14028 33516 14084 33572
rect 13692 32732 13748 32788
rect 14700 37490 14756 37492
rect 14700 37438 14702 37490
rect 14702 37438 14754 37490
rect 14754 37438 14756 37490
rect 14700 37436 14756 37438
rect 22652 38220 22708 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 19516 38050 19572 38052
rect 19516 37998 19518 38050
rect 19518 37998 19570 38050
rect 19570 37998 19572 38050
rect 19516 37996 19572 37998
rect 19964 38050 20020 38052
rect 19964 37998 19966 38050
rect 19966 37998 20018 38050
rect 20018 37998 20020 38050
rect 19964 37996 20020 37998
rect 21308 37938 21364 37940
rect 21308 37886 21310 37938
rect 21310 37886 21362 37938
rect 21362 37886 21364 37938
rect 21308 37884 21364 37886
rect 20972 37826 21028 37828
rect 20972 37774 20974 37826
rect 20974 37774 21026 37826
rect 21026 37774 21028 37826
rect 20972 37772 21028 37774
rect 21644 37772 21700 37828
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 32732 38220 32788 38276
rect 33852 38274 33908 38276
rect 33852 38222 33854 38274
rect 33854 38222 33906 38274
rect 33906 38222 33908 38274
rect 33852 38220 33908 38222
rect 36092 38220 36148 38276
rect 37324 38274 37380 38276
rect 37324 38222 37326 38274
rect 37326 38222 37378 38274
rect 37378 38222 37380 38274
rect 37324 38220 37380 38222
rect 28700 37996 28756 38052
rect 26012 37436 26068 37492
rect 27244 37490 27300 37492
rect 27244 37438 27246 37490
rect 27246 37438 27298 37490
rect 27298 37438 27300 37490
rect 27244 37436 27300 37438
rect 14700 36428 14756 36484
rect 15148 36764 15204 36820
rect 15260 36652 15316 36708
rect 14588 36316 14644 36372
rect 15260 36370 15316 36372
rect 15260 36318 15262 36370
rect 15262 36318 15314 36370
rect 15314 36318 15316 36370
rect 15260 36316 15316 36318
rect 15596 36092 15652 36148
rect 16044 36092 16100 36148
rect 16380 34914 16436 34916
rect 16380 34862 16382 34914
rect 16382 34862 16434 34914
rect 16434 34862 16436 34914
rect 16380 34860 16436 34862
rect 16492 35308 16548 35364
rect 14700 34130 14756 34132
rect 14700 34078 14702 34130
rect 14702 34078 14754 34130
rect 14754 34078 14756 34130
rect 14700 34076 14756 34078
rect 16044 34130 16100 34132
rect 16044 34078 16046 34130
rect 16046 34078 16098 34130
rect 16098 34078 16100 34130
rect 16044 34076 16100 34078
rect 15148 33852 15204 33908
rect 14140 32562 14196 32564
rect 14140 32510 14142 32562
rect 14142 32510 14194 32562
rect 14194 32510 14196 32562
rect 14140 32508 14196 32510
rect 12796 31836 12852 31892
rect 13244 31836 13300 31892
rect 13020 31724 13076 31780
rect 14588 32396 14644 32452
rect 13356 31500 13412 31556
rect 12908 30828 12964 30884
rect 12460 30156 12516 30212
rect 12236 29932 12292 29988
rect 12124 29708 12180 29764
rect 11900 29426 11956 29428
rect 11900 29374 11902 29426
rect 11902 29374 11954 29426
rect 11954 29374 11956 29426
rect 11900 29372 11956 29374
rect 12572 29820 12628 29876
rect 13244 29708 13300 29764
rect 12796 29484 12852 29540
rect 12012 29314 12068 29316
rect 12012 29262 12014 29314
rect 12014 29262 12066 29314
rect 12066 29262 12068 29314
rect 12012 29260 12068 29262
rect 12460 29036 12516 29092
rect 11900 28754 11956 28756
rect 11900 28702 11902 28754
rect 11902 28702 11954 28754
rect 11954 28702 11956 28754
rect 11900 28700 11956 28702
rect 12460 28700 12516 28756
rect 12236 28364 12292 28420
rect 13244 29260 13300 29316
rect 11788 26908 11844 26964
rect 12124 26460 12180 26516
rect 11788 25506 11844 25508
rect 11788 25454 11790 25506
rect 11790 25454 11842 25506
rect 11842 25454 11844 25506
rect 11788 25452 11844 25454
rect 11676 24892 11732 24948
rect 12348 24332 12404 24388
rect 11116 23324 11172 23380
rect 11452 23436 11508 23492
rect 11116 23042 11172 23044
rect 11116 22990 11118 23042
rect 11118 22990 11170 23042
rect 11170 22990 11172 23042
rect 11116 22988 11172 22990
rect 11228 22876 11284 22932
rect 11340 23154 11396 23156
rect 11340 23102 11342 23154
rect 11342 23102 11394 23154
rect 11394 23102 11396 23154
rect 11340 23100 11396 23102
rect 11004 22428 11060 22484
rect 11004 22092 11060 22148
rect 11228 21308 11284 21364
rect 11228 20972 11284 21028
rect 10780 20578 10836 20580
rect 10780 20526 10782 20578
rect 10782 20526 10834 20578
rect 10834 20526 10836 20578
rect 10780 20524 10836 20526
rect 10780 20130 10836 20132
rect 10780 20078 10782 20130
rect 10782 20078 10834 20130
rect 10834 20078 10836 20130
rect 10780 20076 10836 20078
rect 10780 19122 10836 19124
rect 10780 19070 10782 19122
rect 10782 19070 10834 19122
rect 10834 19070 10836 19122
rect 10780 19068 10836 19070
rect 11564 22092 11620 22148
rect 11676 21810 11732 21812
rect 11676 21758 11678 21810
rect 11678 21758 11730 21810
rect 11730 21758 11732 21810
rect 11676 21756 11732 21758
rect 11564 21308 11620 21364
rect 11340 19404 11396 19460
rect 11228 19068 11284 19124
rect 11004 18956 11060 19012
rect 10780 18844 10836 18900
rect 10668 17052 10724 17108
rect 10444 16828 10500 16884
rect 10444 16098 10500 16100
rect 10444 16046 10446 16098
rect 10446 16046 10498 16098
rect 10498 16046 10500 16098
rect 10444 16044 10500 16046
rect 10220 15986 10276 15988
rect 10220 15934 10222 15986
rect 10222 15934 10274 15986
rect 10274 15934 10276 15986
rect 10220 15932 10276 15934
rect 10556 15708 10612 15764
rect 10668 16716 10724 16772
rect 10780 16044 10836 16100
rect 10780 15820 10836 15876
rect 9884 14306 9940 14308
rect 9884 14254 9886 14306
rect 9886 14254 9938 14306
rect 9938 14254 9940 14306
rect 9884 14252 9940 14254
rect 11004 17388 11060 17444
rect 10892 15538 10948 15540
rect 10892 15486 10894 15538
rect 10894 15486 10946 15538
rect 10946 15486 10948 15538
rect 10892 15484 10948 15486
rect 11004 15372 11060 15428
rect 10332 13970 10388 13972
rect 10332 13918 10334 13970
rect 10334 13918 10386 13970
rect 10386 13918 10388 13970
rect 10332 13916 10388 13918
rect 11340 17948 11396 18004
rect 11228 17666 11284 17668
rect 11228 17614 11230 17666
rect 11230 17614 11282 17666
rect 11282 17614 11284 17666
rect 11228 17612 11284 17614
rect 11228 16994 11284 16996
rect 11228 16942 11230 16994
rect 11230 16942 11282 16994
rect 11282 16942 11284 16994
rect 11228 16940 11284 16942
rect 14140 31052 14196 31108
rect 13692 30994 13748 30996
rect 13692 30942 13694 30994
rect 13694 30942 13746 30994
rect 13746 30942 13748 30994
rect 13692 30940 13748 30942
rect 13580 29708 13636 29764
rect 14252 30380 14308 30436
rect 13692 29484 13748 29540
rect 13916 29484 13972 29540
rect 13132 29036 13188 29092
rect 12908 27692 12964 27748
rect 12796 27020 12852 27076
rect 12796 26852 12852 26908
rect 12124 22876 12180 22932
rect 13020 26572 13076 26628
rect 13132 26236 13188 26292
rect 13580 29314 13636 29316
rect 13580 29262 13582 29314
rect 13582 29262 13634 29314
rect 13634 29262 13636 29314
rect 13580 29260 13636 29262
rect 13468 29036 13524 29092
rect 14028 29426 14084 29428
rect 14028 29374 14030 29426
rect 14030 29374 14082 29426
rect 14082 29374 14084 29426
rect 14028 29372 14084 29374
rect 14364 30268 14420 30324
rect 14700 30882 14756 30884
rect 14700 30830 14702 30882
rect 14702 30830 14754 30882
rect 14754 30830 14756 30882
rect 14700 30828 14756 30830
rect 14588 29708 14644 29764
rect 14700 30044 14756 30100
rect 14028 28476 14084 28532
rect 13244 26348 13300 26404
rect 13356 28418 13412 28420
rect 13356 28366 13358 28418
rect 13358 28366 13410 28418
rect 13410 28366 13412 28418
rect 13356 28364 13412 28366
rect 12908 25618 12964 25620
rect 12908 25566 12910 25618
rect 12910 25566 12962 25618
rect 12962 25566 12964 25618
rect 12908 25564 12964 25566
rect 12908 25116 12964 25172
rect 12684 24444 12740 24500
rect 12572 22764 12628 22820
rect 12684 23884 12740 23940
rect 12460 22258 12516 22260
rect 12460 22206 12462 22258
rect 12462 22206 12514 22258
rect 12514 22206 12516 22258
rect 12460 22204 12516 22206
rect 12124 21644 12180 21700
rect 12124 21474 12180 21476
rect 12124 21422 12126 21474
rect 12126 21422 12178 21474
rect 12178 21422 12180 21474
rect 12124 21420 12180 21422
rect 12460 21756 12516 21812
rect 12908 22764 12964 22820
rect 12908 21868 12964 21924
rect 13580 28140 13636 28196
rect 13692 27970 13748 27972
rect 13692 27918 13694 27970
rect 13694 27918 13746 27970
rect 13746 27918 13748 27970
rect 13692 27916 13748 27918
rect 14364 29036 14420 29092
rect 14140 28140 14196 28196
rect 14252 28364 14308 28420
rect 14028 27692 14084 27748
rect 13580 27356 13636 27412
rect 13580 26460 13636 26516
rect 14028 27132 14084 27188
rect 13468 26348 13524 26404
rect 13580 26124 13636 26180
rect 13580 25676 13636 25732
rect 13468 25282 13524 25284
rect 13468 25230 13470 25282
rect 13470 25230 13522 25282
rect 13522 25230 13524 25282
rect 13468 25228 13524 25230
rect 13356 25116 13412 25172
rect 13468 23772 13524 23828
rect 13244 23548 13300 23604
rect 13244 22876 13300 22932
rect 12572 21532 12628 21588
rect 13244 21868 13300 21924
rect 11564 17106 11620 17108
rect 11564 17054 11566 17106
rect 11566 17054 11618 17106
rect 11618 17054 11620 17106
rect 11564 17052 11620 17054
rect 11900 18956 11956 19012
rect 12012 17836 12068 17892
rect 12460 20130 12516 20132
rect 12460 20078 12462 20130
rect 12462 20078 12514 20130
rect 12514 20078 12516 20130
rect 12460 20076 12516 20078
rect 12348 19404 12404 19460
rect 12348 18732 12404 18788
rect 12012 17666 12068 17668
rect 12012 17614 12014 17666
rect 12014 17614 12066 17666
rect 12066 17614 12068 17666
rect 12012 17612 12068 17614
rect 11452 16940 11508 16996
rect 12572 16940 12628 16996
rect 12236 16268 12292 16324
rect 12460 16882 12516 16884
rect 12460 16830 12462 16882
rect 12462 16830 12514 16882
rect 12514 16830 12516 16882
rect 12460 16828 12516 16830
rect 12796 21196 12852 21252
rect 13580 22482 13636 22484
rect 13580 22430 13582 22482
rect 13582 22430 13634 22482
rect 13634 22430 13636 22482
rect 13580 22428 13636 22430
rect 13580 21644 13636 21700
rect 13580 20972 13636 21028
rect 13468 20636 13524 20692
rect 12908 19234 12964 19236
rect 12908 19182 12910 19234
rect 12910 19182 12962 19234
rect 12962 19182 12964 19234
rect 12908 19180 12964 19182
rect 12796 19068 12852 19124
rect 14588 29260 14644 29316
rect 15036 33068 15092 33124
rect 15708 34018 15764 34020
rect 15708 33966 15710 34018
rect 15710 33966 15762 34018
rect 15762 33966 15764 34018
rect 15708 33964 15764 33966
rect 15596 33458 15652 33460
rect 15596 33406 15598 33458
rect 15598 33406 15650 33458
rect 15650 33406 15652 33458
rect 15596 33404 15652 33406
rect 15260 33234 15316 33236
rect 15260 33182 15262 33234
rect 15262 33182 15314 33234
rect 15314 33182 15316 33234
rect 15260 33180 15316 33182
rect 15484 33122 15540 33124
rect 15484 33070 15486 33122
rect 15486 33070 15538 33122
rect 15538 33070 15540 33122
rect 15484 33068 15540 33070
rect 15036 32508 15092 32564
rect 15148 31666 15204 31668
rect 15148 31614 15150 31666
rect 15150 31614 15202 31666
rect 15202 31614 15204 31666
rect 15148 31612 15204 31614
rect 15036 31276 15092 31332
rect 15148 31106 15204 31108
rect 15148 31054 15150 31106
rect 15150 31054 15202 31106
rect 15202 31054 15204 31106
rect 15148 31052 15204 31054
rect 15148 30492 15204 30548
rect 15372 32732 15428 32788
rect 15484 32396 15540 32452
rect 15596 31948 15652 32004
rect 15372 31612 15428 31668
rect 15372 30156 15428 30212
rect 16268 33516 16324 33572
rect 16492 34130 16548 34132
rect 16492 34078 16494 34130
rect 16494 34078 16546 34130
rect 16546 34078 16548 34130
rect 16492 34076 16548 34078
rect 16380 33122 16436 33124
rect 16380 33070 16382 33122
rect 16382 33070 16434 33122
rect 16434 33070 16436 33122
rect 16380 33068 16436 33070
rect 16492 32620 16548 32676
rect 16268 32338 16324 32340
rect 16268 32286 16270 32338
rect 16270 32286 16322 32338
rect 16322 32286 16324 32338
rect 16268 32284 16324 32286
rect 16044 32172 16100 32228
rect 16044 31836 16100 31892
rect 16268 31948 16324 32004
rect 15596 31666 15652 31668
rect 15596 31614 15598 31666
rect 15598 31614 15650 31666
rect 15650 31614 15652 31666
rect 15596 31612 15652 31614
rect 16044 31500 16100 31556
rect 17388 35532 17444 35588
rect 16828 32732 16884 32788
rect 16380 31612 16436 31668
rect 14924 29484 14980 29540
rect 15148 29426 15204 29428
rect 15148 29374 15150 29426
rect 15150 29374 15202 29426
rect 15202 29374 15204 29426
rect 15148 29372 15204 29374
rect 15260 29148 15316 29204
rect 14700 29036 14756 29092
rect 15372 28700 15428 28756
rect 14364 27692 14420 27748
rect 14252 26460 14308 26516
rect 14476 26796 14532 26852
rect 14028 25452 14084 25508
rect 13804 22428 13860 22484
rect 14476 26012 14532 26068
rect 14252 24668 14308 24724
rect 14028 24610 14084 24612
rect 14028 24558 14030 24610
rect 14030 24558 14082 24610
rect 14082 24558 14084 24610
rect 14028 24556 14084 24558
rect 14140 23938 14196 23940
rect 14140 23886 14142 23938
rect 14142 23886 14194 23938
rect 14194 23886 14196 23938
rect 14140 23884 14196 23886
rect 14140 23548 14196 23604
rect 13804 21308 13860 21364
rect 13916 21868 13972 21924
rect 13804 20300 13860 20356
rect 14028 21698 14084 21700
rect 14028 21646 14030 21698
rect 14030 21646 14082 21698
rect 14082 21646 14084 21698
rect 14028 21644 14084 21646
rect 14028 21196 14084 21252
rect 14140 21532 14196 21588
rect 13692 19180 13748 19236
rect 14028 19516 14084 19572
rect 14028 19234 14084 19236
rect 14028 19182 14030 19234
rect 14030 19182 14082 19234
rect 14082 19182 14084 19234
rect 14028 19180 14084 19182
rect 13020 17612 13076 17668
rect 14028 18396 14084 18452
rect 13580 17778 13636 17780
rect 13580 17726 13582 17778
rect 13582 17726 13634 17778
rect 13634 17726 13636 17778
rect 13580 17724 13636 17726
rect 13468 17666 13524 17668
rect 13468 17614 13470 17666
rect 13470 17614 13522 17666
rect 13522 17614 13524 17666
rect 13468 17612 13524 17614
rect 13356 17276 13412 17332
rect 13468 17052 13524 17108
rect 11676 16156 11732 16212
rect 11228 15426 11284 15428
rect 11228 15374 11230 15426
rect 11230 15374 11282 15426
rect 11282 15374 11284 15426
rect 11228 15372 11284 15374
rect 11788 16098 11844 16100
rect 11788 16046 11790 16098
rect 11790 16046 11842 16098
rect 11842 16046 11844 16098
rect 11788 16044 11844 16046
rect 12460 16098 12516 16100
rect 12460 16046 12462 16098
rect 12462 16046 12514 16098
rect 12514 16046 12516 16098
rect 12460 16044 12516 16046
rect 12236 15932 12292 15988
rect 11900 15874 11956 15876
rect 11900 15822 11902 15874
rect 11902 15822 11954 15874
rect 11954 15822 11956 15874
rect 11900 15820 11956 15822
rect 12572 15820 12628 15876
rect 11676 15484 11732 15540
rect 12572 15314 12628 15316
rect 12572 15262 12574 15314
rect 12574 15262 12626 15314
rect 12626 15262 12628 15314
rect 12572 15260 12628 15262
rect 11676 15202 11732 15204
rect 11676 15150 11678 15202
rect 11678 15150 11730 15202
rect 11730 15150 11732 15202
rect 11676 15148 11732 15150
rect 13020 15484 13076 15540
rect 12908 15426 12964 15428
rect 12908 15374 12910 15426
rect 12910 15374 12962 15426
rect 12962 15374 12964 15426
rect 12908 15372 12964 15374
rect 12796 15036 12852 15092
rect 13244 16268 13300 16324
rect 14140 17724 14196 17780
rect 14140 17388 14196 17444
rect 14476 23100 14532 23156
rect 14588 24892 14644 24948
rect 14364 22428 14420 22484
rect 14364 20860 14420 20916
rect 14028 17052 14084 17108
rect 13580 16604 13636 16660
rect 13244 16044 13300 16100
rect 15708 29148 15764 29204
rect 14812 27132 14868 27188
rect 14924 27692 14980 27748
rect 15036 27132 15092 27188
rect 15148 27074 15204 27076
rect 15148 27022 15150 27074
rect 15150 27022 15202 27074
rect 15202 27022 15204 27074
rect 15148 27020 15204 27022
rect 15148 26796 15204 26852
rect 15484 28252 15540 28308
rect 15484 27580 15540 27636
rect 15484 27244 15540 27300
rect 15708 28530 15764 28532
rect 15708 28478 15710 28530
rect 15710 28478 15762 28530
rect 15762 28478 15764 28530
rect 15708 28476 15764 28478
rect 15932 30210 15988 30212
rect 15932 30158 15934 30210
rect 15934 30158 15986 30210
rect 15986 30158 15988 30210
rect 15932 30156 15988 30158
rect 19836 36090 19892 36092
rect 19628 35980 19684 36036
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 17836 35308 17892 35364
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 17052 33404 17108 33460
rect 17500 33122 17556 33124
rect 17500 33070 17502 33122
rect 17502 33070 17554 33122
rect 17554 33070 17556 33122
rect 17500 33068 17556 33070
rect 17276 32844 17332 32900
rect 17388 32674 17444 32676
rect 17388 32622 17390 32674
rect 17390 32622 17442 32674
rect 17442 32622 17444 32674
rect 17388 32620 17444 32622
rect 16940 31836 16996 31892
rect 16604 31276 16660 31332
rect 16380 30604 16436 30660
rect 16044 29820 16100 29876
rect 16380 30380 16436 30436
rect 16716 30828 16772 30884
rect 16492 30268 16548 30324
rect 16492 29820 16548 29876
rect 15708 27804 15764 27860
rect 15708 27244 15764 27300
rect 15484 26684 15540 26740
rect 14812 25506 14868 25508
rect 14812 25454 14814 25506
rect 14814 25454 14866 25506
rect 14866 25454 14868 25506
rect 14812 25452 14868 25454
rect 15372 25228 15428 25284
rect 15596 26236 15652 26292
rect 15372 24946 15428 24948
rect 15372 24894 15374 24946
rect 15374 24894 15426 24946
rect 15426 24894 15428 24946
rect 15372 24892 15428 24894
rect 14700 23938 14756 23940
rect 14700 23886 14702 23938
rect 14702 23886 14754 23938
rect 14754 23886 14756 23938
rect 14700 23884 14756 23886
rect 14924 23996 14980 24052
rect 14924 23100 14980 23156
rect 14812 22146 14868 22148
rect 14812 22094 14814 22146
rect 14814 22094 14866 22146
rect 14866 22094 14868 22146
rect 14812 22092 14868 22094
rect 14700 21084 14756 21140
rect 14700 20860 14756 20916
rect 15148 20802 15204 20804
rect 15148 20750 15150 20802
rect 15150 20750 15202 20802
rect 15202 20750 15204 20802
rect 15148 20748 15204 20750
rect 15148 20018 15204 20020
rect 15148 19966 15150 20018
rect 15150 19966 15202 20018
rect 15202 19966 15204 20018
rect 15148 19964 15204 19966
rect 14812 19234 14868 19236
rect 14812 19182 14814 19234
rect 14814 19182 14866 19234
rect 14866 19182 14868 19234
rect 14812 19180 14868 19182
rect 14588 18396 14644 18452
rect 14588 17442 14644 17444
rect 14588 17390 14590 17442
rect 14590 17390 14642 17442
rect 14642 17390 14644 17442
rect 14588 17388 14644 17390
rect 14364 16940 14420 16996
rect 14140 16604 14196 16660
rect 13916 16492 13972 16548
rect 13692 16210 13748 16212
rect 13692 16158 13694 16210
rect 13694 16158 13746 16210
rect 13746 16158 13748 16210
rect 13692 16156 13748 16158
rect 13916 15538 13972 15540
rect 13916 15486 13918 15538
rect 13918 15486 13970 15538
rect 13970 15486 13972 15538
rect 13916 15484 13972 15486
rect 13468 15314 13524 15316
rect 13468 15262 13470 15314
rect 13470 15262 13522 15314
rect 13522 15262 13524 15314
rect 13468 15260 13524 15262
rect 14700 16882 14756 16884
rect 14700 16830 14702 16882
rect 14702 16830 14754 16882
rect 14754 16830 14756 16882
rect 14700 16828 14756 16830
rect 14588 16268 14644 16324
rect 14476 15314 14532 15316
rect 14476 15262 14478 15314
rect 14478 15262 14530 15314
rect 14530 15262 14532 15314
rect 14476 15260 14532 15262
rect 14364 15148 14420 15204
rect 14028 14924 14084 14980
rect 14252 14700 14308 14756
rect 12236 14140 12292 14196
rect 12796 13858 12852 13860
rect 12796 13806 12798 13858
rect 12798 13806 12850 13858
rect 12850 13806 12852 13858
rect 12796 13804 12852 13806
rect 13244 13858 13300 13860
rect 13244 13806 13246 13858
rect 13246 13806 13298 13858
rect 13298 13806 13300 13858
rect 13244 13804 13300 13806
rect 14028 14530 14084 14532
rect 14028 14478 14030 14530
rect 14030 14478 14082 14530
rect 14082 14478 14084 14530
rect 14028 14476 14084 14478
rect 14700 15986 14756 15988
rect 14700 15934 14702 15986
rect 14702 15934 14754 15986
rect 14754 15934 14756 15986
rect 14700 15932 14756 15934
rect 15372 22204 15428 22260
rect 15932 29484 15988 29540
rect 16044 29148 16100 29204
rect 16604 29148 16660 29204
rect 16604 28924 16660 28980
rect 16492 28476 16548 28532
rect 16268 28252 16324 28308
rect 16044 27858 16100 27860
rect 16044 27806 16046 27858
rect 16046 27806 16098 27858
rect 16098 27806 16100 27858
rect 16044 27804 16100 27806
rect 16268 27746 16324 27748
rect 16268 27694 16270 27746
rect 16270 27694 16322 27746
rect 16322 27694 16324 27746
rect 16268 27692 16324 27694
rect 15932 26908 15988 26964
rect 16044 27244 16100 27300
rect 15932 25506 15988 25508
rect 15932 25454 15934 25506
rect 15934 25454 15986 25506
rect 15986 25454 15988 25506
rect 15932 25452 15988 25454
rect 16604 27804 16660 27860
rect 16492 26850 16548 26852
rect 16492 26798 16494 26850
rect 16494 26798 16546 26850
rect 16546 26798 16548 26850
rect 16492 26796 16548 26798
rect 16492 26348 16548 26404
rect 15820 24332 15876 24388
rect 15708 22540 15764 22596
rect 15820 22428 15876 22484
rect 16156 23884 16212 23940
rect 16268 24892 16324 24948
rect 16044 22428 16100 22484
rect 15708 20300 15764 20356
rect 15932 21308 15988 21364
rect 15708 19740 15764 19796
rect 15596 19628 15652 19684
rect 15148 18508 15204 18564
rect 15036 18284 15092 18340
rect 15260 18284 15316 18340
rect 15372 19068 15428 19124
rect 15148 17554 15204 17556
rect 15148 17502 15150 17554
rect 15150 17502 15202 17554
rect 15202 17502 15204 17554
rect 15148 17500 15204 17502
rect 15036 17388 15092 17444
rect 15148 16716 15204 16772
rect 16156 22370 16212 22372
rect 16156 22318 16158 22370
rect 16158 22318 16210 22370
rect 16210 22318 16212 22370
rect 16156 22316 16212 22318
rect 16380 23772 16436 23828
rect 16492 22428 16548 22484
rect 16268 21756 16324 21812
rect 16156 20802 16212 20804
rect 16156 20750 16158 20802
rect 16158 20750 16210 20802
rect 16210 20750 16212 20802
rect 16156 20748 16212 20750
rect 16380 21308 16436 21364
rect 16380 20300 16436 20356
rect 15932 19068 15988 19124
rect 15820 18338 15876 18340
rect 15820 18286 15822 18338
rect 15822 18286 15874 18338
rect 15874 18286 15876 18338
rect 15820 18284 15876 18286
rect 16044 18226 16100 18228
rect 16044 18174 16046 18226
rect 16046 18174 16098 18226
rect 16098 18174 16100 18226
rect 16044 18172 16100 18174
rect 15708 17836 15764 17892
rect 15372 17388 15428 17444
rect 15708 17164 15764 17220
rect 15596 17106 15652 17108
rect 15596 17054 15598 17106
rect 15598 17054 15650 17106
rect 15650 17054 15652 17106
rect 15596 17052 15652 17054
rect 15596 16604 15652 16660
rect 15372 16156 15428 16212
rect 14924 16098 14980 16100
rect 14924 16046 14926 16098
rect 14926 16046 14978 16098
rect 14978 16046 14980 16098
rect 14924 16044 14980 16046
rect 15148 15484 15204 15540
rect 14812 15426 14868 15428
rect 14812 15374 14814 15426
rect 14814 15374 14866 15426
rect 14866 15374 14868 15426
rect 14812 15372 14868 15374
rect 16380 18844 16436 18900
rect 16716 27020 16772 27076
rect 16716 22764 16772 22820
rect 17500 31500 17556 31556
rect 17052 30940 17108 30996
rect 18060 33404 18116 33460
rect 19404 33628 19460 33684
rect 19180 33234 19236 33236
rect 19180 33182 19182 33234
rect 19182 33182 19234 33234
rect 19234 33182 19236 33234
rect 19180 33180 19236 33182
rect 18396 33068 18452 33124
rect 18284 32844 18340 32900
rect 18844 32620 18900 32676
rect 21308 33964 21364 34020
rect 19964 33516 20020 33572
rect 20972 33516 21028 33572
rect 18956 32450 19012 32452
rect 18956 32398 18958 32450
rect 18958 32398 19010 32450
rect 19010 32398 19012 32450
rect 18956 32396 19012 32398
rect 19516 32396 19572 32452
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19628 32508 19684 32564
rect 19404 32284 19460 32340
rect 18284 31948 18340 32004
rect 17948 31554 18004 31556
rect 17948 31502 17950 31554
rect 17950 31502 18002 31554
rect 18002 31502 18004 31554
rect 17948 31500 18004 31502
rect 17612 30940 17668 30996
rect 17836 29820 17892 29876
rect 17388 29036 17444 29092
rect 17836 29372 17892 29428
rect 17836 28812 17892 28868
rect 17500 28642 17556 28644
rect 17500 28590 17502 28642
rect 17502 28590 17554 28642
rect 17554 28590 17556 28642
rect 17500 28588 17556 28590
rect 17164 28530 17220 28532
rect 17164 28478 17166 28530
rect 17166 28478 17218 28530
rect 17218 28478 17220 28530
rect 17164 28476 17220 28478
rect 17164 27244 17220 27300
rect 18060 29148 18116 29204
rect 17612 26684 17668 26740
rect 17276 26572 17332 26628
rect 17388 26514 17444 26516
rect 17388 26462 17390 26514
rect 17390 26462 17442 26514
rect 17442 26462 17444 26514
rect 17388 26460 17444 26462
rect 17948 26178 18004 26180
rect 17948 26126 17950 26178
rect 17950 26126 18002 26178
rect 18002 26126 18004 26178
rect 17948 26124 18004 26126
rect 17612 26012 17668 26068
rect 17052 25452 17108 25508
rect 16828 22316 16884 22372
rect 16828 22092 16884 22148
rect 16940 23436 16996 23492
rect 16940 21980 16996 22036
rect 17388 25730 17444 25732
rect 17388 25678 17390 25730
rect 17390 25678 17442 25730
rect 17442 25678 17444 25730
rect 17388 25676 17444 25678
rect 17276 25004 17332 25060
rect 17500 25116 17556 25172
rect 17164 23436 17220 23492
rect 18060 25900 18116 25956
rect 17836 25340 17892 25396
rect 17724 24780 17780 24836
rect 18060 24780 18116 24836
rect 17500 24556 17556 24612
rect 17388 23548 17444 23604
rect 17500 23996 17556 24052
rect 17052 22540 17108 22596
rect 16828 21308 16884 21364
rect 16604 20524 16660 20580
rect 16828 20300 16884 20356
rect 16940 20524 16996 20580
rect 16828 20018 16884 20020
rect 16828 19966 16830 20018
rect 16830 19966 16882 20018
rect 16882 19966 16884 20018
rect 16828 19964 16884 19966
rect 16716 19292 16772 19348
rect 16156 17666 16212 17668
rect 16156 17614 16158 17666
rect 16158 17614 16210 17666
rect 16210 17614 16212 17666
rect 16156 17612 16212 17614
rect 15820 17052 15876 17108
rect 15820 16156 15876 16212
rect 16044 17500 16100 17556
rect 16156 16604 16212 16660
rect 16716 18060 16772 18116
rect 16492 17836 16548 17892
rect 16716 17778 16772 17780
rect 16716 17726 16718 17778
rect 16718 17726 16770 17778
rect 16770 17726 16772 17778
rect 16716 17724 16772 17726
rect 16604 17666 16660 17668
rect 16604 17614 16606 17666
rect 16606 17614 16658 17666
rect 16658 17614 16660 17666
rect 16604 17612 16660 17614
rect 16380 17500 16436 17556
rect 16716 17554 16772 17556
rect 16716 17502 16718 17554
rect 16718 17502 16770 17554
rect 16770 17502 16772 17554
rect 16716 17500 16772 17502
rect 16380 16994 16436 16996
rect 16380 16942 16382 16994
rect 16382 16942 16434 16994
rect 16434 16942 16436 16994
rect 16380 16940 16436 16942
rect 17164 22370 17220 22372
rect 17164 22318 17166 22370
rect 17166 22318 17218 22370
rect 17218 22318 17220 22370
rect 17164 22316 17220 22318
rect 17500 22540 17556 22596
rect 18060 23436 18116 23492
rect 17836 22876 17892 22932
rect 17948 22988 18004 23044
rect 17500 22370 17556 22372
rect 17500 22318 17502 22370
rect 17502 22318 17554 22370
rect 17554 22318 17556 22370
rect 17500 22316 17556 22318
rect 17724 22258 17780 22260
rect 17724 22206 17726 22258
rect 17726 22206 17778 22258
rect 17778 22206 17780 22258
rect 17724 22204 17780 22206
rect 17612 21868 17668 21924
rect 17052 19964 17108 20020
rect 17388 21586 17444 21588
rect 17388 21534 17390 21586
rect 17390 21534 17442 21586
rect 17442 21534 17444 21586
rect 17388 21532 17444 21534
rect 17836 21532 17892 21588
rect 17388 21308 17444 21364
rect 18620 30994 18676 30996
rect 18620 30942 18622 30994
rect 18622 30942 18674 30994
rect 18674 30942 18676 30994
rect 18620 30940 18676 30942
rect 18396 30882 18452 30884
rect 18396 30830 18398 30882
rect 18398 30830 18450 30882
rect 18450 30830 18452 30882
rect 18396 30828 18452 30830
rect 18396 30604 18452 30660
rect 18844 29986 18900 29988
rect 18844 29934 18846 29986
rect 18846 29934 18898 29986
rect 18898 29934 18900 29986
rect 18844 29932 18900 29934
rect 18508 29708 18564 29764
rect 18620 29650 18676 29652
rect 18620 29598 18622 29650
rect 18622 29598 18674 29650
rect 18674 29598 18676 29650
rect 18620 29596 18676 29598
rect 18284 29372 18340 29428
rect 18396 28812 18452 28868
rect 19852 32732 19908 32788
rect 19740 31948 19796 32004
rect 20524 32450 20580 32452
rect 20524 32398 20526 32450
rect 20526 32398 20578 32450
rect 20578 32398 20580 32450
rect 20524 32396 20580 32398
rect 20300 32338 20356 32340
rect 20300 32286 20302 32338
rect 20302 32286 20354 32338
rect 20354 32286 20356 32338
rect 20300 32284 20356 32286
rect 20076 31836 20132 31892
rect 21196 32562 21252 32564
rect 21196 32510 21198 32562
rect 21198 32510 21250 32562
rect 21250 32510 21252 32562
rect 21196 32508 21252 32510
rect 20636 31612 20692 31668
rect 20748 32284 20804 32340
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20524 30716 20580 30772
rect 19852 30044 19908 30100
rect 19404 29820 19460 29876
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20636 29596 20692 29652
rect 18956 29148 19012 29204
rect 18732 28812 18788 28868
rect 18508 28476 18564 28532
rect 18284 28140 18340 28196
rect 18844 28700 18900 28756
rect 19068 28476 19124 28532
rect 18844 27692 18900 27748
rect 19068 27858 19124 27860
rect 19068 27806 19070 27858
rect 19070 27806 19122 27858
rect 19122 27806 19124 27858
rect 19068 27804 19124 27806
rect 18396 27356 18452 27412
rect 18508 27244 18564 27300
rect 18284 26236 18340 26292
rect 18396 27132 18452 27188
rect 19404 29426 19460 29428
rect 19404 29374 19406 29426
rect 19406 29374 19458 29426
rect 19458 29374 19460 29426
rect 19404 29372 19460 29374
rect 19292 28812 19348 28868
rect 20300 28588 20356 28644
rect 20188 28530 20244 28532
rect 20188 28478 20190 28530
rect 20190 28478 20242 28530
rect 20242 28478 20244 28530
rect 20188 28476 20244 28478
rect 19292 28364 19348 28420
rect 19852 28418 19908 28420
rect 19852 28366 19854 28418
rect 19854 28366 19906 28418
rect 19906 28366 19908 28418
rect 19852 28364 19908 28366
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20188 28028 20244 28084
rect 19852 27916 19908 27972
rect 19740 27356 19796 27412
rect 20300 27746 20356 27748
rect 20300 27694 20302 27746
rect 20302 27694 20354 27746
rect 20354 27694 20356 27746
rect 20300 27692 20356 27694
rect 20300 27186 20356 27188
rect 20300 27134 20302 27186
rect 20302 27134 20354 27186
rect 20354 27134 20356 27186
rect 20300 27132 20356 27134
rect 18284 25900 18340 25956
rect 18284 25004 18340 25060
rect 18284 24722 18340 24724
rect 18284 24670 18286 24722
rect 18286 24670 18338 24722
rect 18338 24670 18340 24722
rect 18284 24668 18340 24670
rect 19292 26402 19348 26404
rect 19292 26350 19294 26402
rect 19294 26350 19346 26402
rect 19346 26350 19348 26402
rect 19292 26348 19348 26350
rect 18508 25452 18564 25508
rect 18620 26124 18676 26180
rect 18732 26012 18788 26068
rect 18508 25004 18564 25060
rect 18508 24668 18564 24724
rect 18396 24556 18452 24612
rect 18620 24444 18676 24500
rect 19516 26124 19572 26180
rect 19404 26012 19460 26068
rect 19516 25564 19572 25620
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19852 26460 19908 26516
rect 19740 25394 19796 25396
rect 19740 25342 19742 25394
rect 19742 25342 19794 25394
rect 19794 25342 19796 25394
rect 19740 25340 19796 25342
rect 20412 26796 20468 26852
rect 19964 25564 20020 25620
rect 19964 25394 20020 25396
rect 19964 25342 19966 25394
rect 19966 25342 20018 25394
rect 20018 25342 20020 25394
rect 19964 25340 20020 25342
rect 20412 25900 20468 25956
rect 21308 31890 21364 31892
rect 21308 31838 21310 31890
rect 21310 31838 21362 31890
rect 21362 31838 21364 31890
rect 21308 31836 21364 31838
rect 21532 31778 21588 31780
rect 21532 31726 21534 31778
rect 21534 31726 21586 31778
rect 21586 31726 21588 31778
rect 21532 31724 21588 31726
rect 20972 31218 21028 31220
rect 20972 31166 20974 31218
rect 20974 31166 21026 31218
rect 21026 31166 21028 31218
rect 20972 31164 21028 31166
rect 21308 31106 21364 31108
rect 21308 31054 21310 31106
rect 21310 31054 21362 31106
rect 21362 31054 21364 31106
rect 21308 31052 21364 31054
rect 21084 30828 21140 30884
rect 20972 29372 21028 29428
rect 21532 30380 21588 30436
rect 22540 31890 22596 31892
rect 22540 31838 22542 31890
rect 22542 31838 22594 31890
rect 22594 31838 22596 31890
rect 22540 31836 22596 31838
rect 22764 31836 22820 31892
rect 22316 31612 22372 31668
rect 21980 31500 22036 31556
rect 22652 31554 22708 31556
rect 22652 31502 22654 31554
rect 22654 31502 22706 31554
rect 22706 31502 22708 31554
rect 22652 31500 22708 31502
rect 22204 31164 22260 31220
rect 22428 31052 22484 31108
rect 21980 30716 22036 30772
rect 22428 30268 22484 30324
rect 21868 29708 21924 29764
rect 21420 29538 21476 29540
rect 21420 29486 21422 29538
rect 21422 29486 21474 29538
rect 21474 29486 21476 29538
rect 21420 29484 21476 29486
rect 22652 31164 22708 31220
rect 22876 31164 22932 31220
rect 23100 31612 23156 31668
rect 23100 31052 23156 31108
rect 22988 30604 23044 30660
rect 22988 30098 23044 30100
rect 22988 30046 22990 30098
rect 22990 30046 23042 30098
rect 23042 30046 23044 30098
rect 22988 30044 23044 30046
rect 21868 29260 21924 29316
rect 21756 28754 21812 28756
rect 21756 28702 21758 28754
rect 21758 28702 21810 28754
rect 21810 28702 21812 28754
rect 21756 28700 21812 28702
rect 20748 27916 20804 27972
rect 21420 27356 21476 27412
rect 22428 28642 22484 28644
rect 22428 28590 22430 28642
rect 22430 28590 22482 28642
rect 22482 28590 22484 28642
rect 22428 28588 22484 28590
rect 22540 27468 22596 27524
rect 21980 27244 22036 27300
rect 22316 27298 22372 27300
rect 22316 27246 22318 27298
rect 22318 27246 22370 27298
rect 22370 27246 22372 27298
rect 22316 27244 22372 27246
rect 20636 27132 20692 27188
rect 21644 26850 21700 26852
rect 21644 26798 21646 26850
rect 21646 26798 21698 26850
rect 21698 26798 21700 26850
rect 21644 26796 21700 26798
rect 21532 26460 21588 26516
rect 22316 26962 22372 26964
rect 22316 26910 22318 26962
rect 22318 26910 22370 26962
rect 22370 26910 22372 26962
rect 22316 26908 22372 26910
rect 21980 26796 22036 26852
rect 21084 26290 21140 26292
rect 21084 26238 21086 26290
rect 21086 26238 21138 26290
rect 21138 26238 21140 26290
rect 21084 26236 21140 26238
rect 21308 25900 21364 25956
rect 20524 25506 20580 25508
rect 20524 25454 20526 25506
rect 20526 25454 20578 25506
rect 20578 25454 20580 25506
rect 20524 25452 20580 25454
rect 21644 25900 21700 25956
rect 20636 25564 20692 25620
rect 19180 25116 19236 25172
rect 19404 25228 19460 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19180 24834 19236 24836
rect 19180 24782 19182 24834
rect 19182 24782 19234 24834
rect 19234 24782 19236 24834
rect 19180 24780 19236 24782
rect 20412 25340 20468 25396
rect 19404 24444 19460 24500
rect 18508 23548 18564 23604
rect 18396 23212 18452 23268
rect 17948 21308 18004 21364
rect 18172 22428 18228 22484
rect 18284 22876 18340 22932
rect 17836 20412 17892 20468
rect 17724 20018 17780 20020
rect 17724 19966 17726 20018
rect 17726 19966 17778 20018
rect 17778 19966 17780 20018
rect 17724 19964 17780 19966
rect 18172 19852 18228 19908
rect 17276 18284 17332 18340
rect 17724 18508 17780 18564
rect 17500 17612 17556 17668
rect 17612 17106 17668 17108
rect 17612 17054 17614 17106
rect 17614 17054 17666 17106
rect 17666 17054 17668 17106
rect 17612 17052 17668 17054
rect 17948 18450 18004 18452
rect 17948 18398 17950 18450
rect 17950 18398 18002 18450
rect 18002 18398 18004 18450
rect 17948 18396 18004 18398
rect 18732 23660 18788 23716
rect 18956 23548 19012 23604
rect 19180 23548 19236 23604
rect 19964 24556 20020 24612
rect 20412 24444 20468 24500
rect 20300 23938 20356 23940
rect 20300 23886 20302 23938
rect 20302 23886 20354 23938
rect 20354 23886 20356 23938
rect 20300 23884 20356 23886
rect 20972 25452 21028 25508
rect 20748 25282 20804 25284
rect 20748 25230 20750 25282
rect 20750 25230 20802 25282
rect 20802 25230 20804 25282
rect 20748 25228 20804 25230
rect 19628 23772 19684 23828
rect 20412 23714 20468 23716
rect 20412 23662 20414 23714
rect 20414 23662 20466 23714
rect 20466 23662 20468 23714
rect 20412 23660 20468 23662
rect 19068 23324 19124 23380
rect 18732 22988 18788 23044
rect 18956 22876 19012 22932
rect 18732 22540 18788 22596
rect 18508 22482 18564 22484
rect 18508 22430 18510 22482
rect 18510 22430 18562 22482
rect 18562 22430 18564 22482
rect 18508 22428 18564 22430
rect 18508 22092 18564 22148
rect 19516 23212 19572 23268
rect 19404 22988 19460 23044
rect 19292 22092 19348 22148
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18844 21756 18900 21812
rect 18956 21644 19012 21700
rect 19404 21586 19460 21588
rect 19404 21534 19406 21586
rect 19406 21534 19458 21586
rect 19458 21534 19460 21586
rect 19404 21532 19460 21534
rect 18508 19292 18564 19348
rect 18284 19068 18340 19124
rect 18396 19180 18452 19236
rect 18284 18674 18340 18676
rect 18284 18622 18286 18674
rect 18286 18622 18338 18674
rect 18338 18622 18340 18674
rect 18284 18620 18340 18622
rect 18172 18562 18228 18564
rect 18172 18510 18174 18562
rect 18174 18510 18226 18562
rect 18226 18510 18228 18562
rect 18172 18508 18228 18510
rect 18508 18508 18564 18564
rect 18396 18284 18452 18340
rect 18396 17948 18452 18004
rect 18060 17442 18116 17444
rect 18060 17390 18062 17442
rect 18062 17390 18114 17442
rect 18114 17390 18116 17442
rect 18060 17388 18116 17390
rect 17948 17276 18004 17332
rect 16604 16882 16660 16884
rect 16604 16830 16606 16882
rect 16606 16830 16658 16882
rect 16658 16830 16660 16882
rect 16604 16828 16660 16830
rect 17836 16882 17892 16884
rect 17836 16830 17838 16882
rect 17838 16830 17890 16882
rect 17890 16830 17892 16882
rect 17836 16828 17892 16830
rect 18060 17052 18116 17108
rect 16380 16716 16436 16772
rect 17612 16268 17668 16324
rect 16380 16098 16436 16100
rect 16380 16046 16382 16098
rect 16382 16046 16434 16098
rect 16434 16046 16436 16098
rect 16380 16044 16436 16046
rect 15932 15932 15988 15988
rect 16156 15986 16212 15988
rect 16156 15934 16158 15986
rect 16158 15934 16210 15986
rect 16210 15934 16212 15986
rect 16156 15932 16212 15934
rect 15820 15820 15876 15876
rect 16044 15874 16100 15876
rect 16044 15822 16046 15874
rect 16046 15822 16098 15874
rect 16098 15822 16100 15874
rect 16044 15820 16100 15822
rect 17500 16098 17556 16100
rect 17500 16046 17502 16098
rect 17502 16046 17554 16098
rect 17554 16046 17556 16098
rect 17500 16044 17556 16046
rect 17052 15708 17108 15764
rect 16380 15596 16436 15652
rect 15372 14700 15428 14756
rect 15372 14530 15428 14532
rect 15372 14478 15374 14530
rect 15374 14478 15426 14530
rect 15426 14478 15428 14530
rect 15372 14476 15428 14478
rect 16380 15372 16436 15428
rect 16156 15314 16212 15316
rect 16156 15262 16158 15314
rect 16158 15262 16210 15314
rect 16210 15262 16212 15314
rect 16156 15260 16212 15262
rect 16268 14700 16324 14756
rect 16156 14642 16212 14644
rect 16156 14590 16158 14642
rect 16158 14590 16210 14642
rect 16210 14590 16212 14642
rect 16156 14588 16212 14590
rect 17164 15820 17220 15876
rect 18172 16828 18228 16884
rect 17276 15484 17332 15540
rect 16268 13970 16324 13972
rect 16268 13918 16270 13970
rect 16270 13918 16322 13970
rect 16322 13918 16324 13970
rect 16268 13916 16324 13918
rect 18620 17836 18676 17892
rect 18508 17500 18564 17556
rect 18508 15932 18564 15988
rect 19292 20802 19348 20804
rect 19292 20750 19294 20802
rect 19294 20750 19346 20802
rect 19346 20750 19348 20802
rect 19292 20748 19348 20750
rect 19404 20412 19460 20468
rect 19404 19964 19460 20020
rect 18844 19292 18900 19348
rect 19180 19122 19236 19124
rect 19180 19070 19182 19122
rect 19182 19070 19234 19122
rect 19234 19070 19236 19122
rect 19180 19068 19236 19070
rect 18844 18396 18900 18452
rect 18844 18172 18900 18228
rect 19180 18450 19236 18452
rect 19180 18398 19182 18450
rect 19182 18398 19234 18450
rect 19234 18398 19236 18450
rect 19180 18396 19236 18398
rect 19180 18060 19236 18116
rect 18956 17948 19012 18004
rect 18844 17666 18900 17668
rect 18844 17614 18846 17666
rect 18846 17614 18898 17666
rect 18898 17614 18900 17666
rect 18844 17612 18900 17614
rect 18956 17442 19012 17444
rect 18956 17390 18958 17442
rect 18958 17390 19010 17442
rect 19010 17390 19012 17442
rect 18956 17388 19012 17390
rect 18844 17276 18900 17332
rect 21308 25228 21364 25284
rect 21420 25340 21476 25396
rect 21196 23772 21252 23828
rect 21868 23996 21924 24052
rect 21420 23714 21476 23716
rect 21420 23662 21422 23714
rect 21422 23662 21474 23714
rect 21474 23662 21476 23714
rect 21420 23660 21476 23662
rect 20860 23100 20916 23156
rect 20076 22540 20132 22596
rect 19628 22428 19684 22484
rect 19852 22092 19908 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20636 22482 20692 22484
rect 20636 22430 20638 22482
rect 20638 22430 20690 22482
rect 20690 22430 20692 22482
rect 20636 22428 20692 22430
rect 20412 21084 20468 21140
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20748 21980 20804 22036
rect 20860 21868 20916 21924
rect 20860 21644 20916 21700
rect 20748 20972 20804 21028
rect 20524 20860 20580 20916
rect 20188 19906 20244 19908
rect 20188 19854 20190 19906
rect 20190 19854 20242 19906
rect 20242 19854 20244 19906
rect 20188 19852 20244 19854
rect 19964 19516 20020 19572
rect 21084 21980 21140 22036
rect 21308 21644 21364 21700
rect 21420 21756 21476 21812
rect 21308 21196 21364 21252
rect 21084 21084 21140 21140
rect 21420 20860 21476 20916
rect 19628 18956 19684 19012
rect 20300 19010 20356 19012
rect 20300 18958 20302 19010
rect 20302 18958 20354 19010
rect 20354 18958 20356 19010
rect 20300 18956 20356 18958
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20188 18844 20244 18900
rect 19964 18620 20020 18676
rect 19404 18172 19460 18228
rect 19628 17948 19684 18004
rect 18844 16156 18900 16212
rect 18620 15314 18676 15316
rect 18620 15262 18622 15314
rect 18622 15262 18674 15314
rect 18674 15262 18676 15314
rect 18620 15260 18676 15262
rect 19180 17052 19236 17108
rect 19068 16268 19124 16324
rect 20076 17948 20132 18004
rect 20076 17554 20132 17556
rect 20076 17502 20078 17554
rect 20078 17502 20130 17554
rect 20130 17502 20132 17554
rect 20076 17500 20132 17502
rect 19740 17388 19796 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 17106 19684 17108
rect 19628 17054 19630 17106
rect 19630 17054 19682 17106
rect 19682 17054 19684 17106
rect 19628 17052 19684 17054
rect 20300 18172 20356 18228
rect 19852 16940 19908 16996
rect 19516 16770 19572 16772
rect 19516 16718 19518 16770
rect 19518 16718 19570 16770
rect 19570 16718 19572 16770
rect 19516 16716 19572 16718
rect 19740 16098 19796 16100
rect 19740 16046 19742 16098
rect 19742 16046 19794 16098
rect 19794 16046 19796 16098
rect 19740 16044 19796 16046
rect 19404 15932 19460 15988
rect 19516 15484 19572 15540
rect 19628 15820 19684 15876
rect 20188 16770 20244 16772
rect 20188 16718 20190 16770
rect 20190 16718 20242 16770
rect 20242 16718 20244 16770
rect 20188 16716 20244 16718
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19740 15148 19796 15204
rect 18508 14588 18564 14644
rect 16940 13916 16996 13972
rect 18060 13970 18116 13972
rect 18060 13918 18062 13970
rect 18062 13918 18114 13970
rect 18114 13918 18116 13970
rect 18060 13916 18116 13918
rect 20412 17612 20468 17668
rect 20636 18172 20692 18228
rect 21868 22652 21924 22708
rect 21756 21810 21812 21812
rect 21756 21758 21758 21810
rect 21758 21758 21810 21810
rect 21810 21758 21812 21810
rect 21756 21756 21812 21758
rect 21644 20860 21700 20916
rect 20860 20412 20916 20468
rect 21868 20636 21924 20692
rect 21532 20130 21588 20132
rect 21532 20078 21534 20130
rect 21534 20078 21586 20130
rect 21586 20078 21588 20130
rect 21532 20076 21588 20078
rect 21420 19964 21476 20020
rect 21084 19906 21140 19908
rect 21084 19854 21086 19906
rect 21086 19854 21138 19906
rect 21138 19854 21140 19906
rect 21084 19852 21140 19854
rect 20860 19628 20916 19684
rect 21420 19292 21476 19348
rect 21532 19122 21588 19124
rect 21532 19070 21534 19122
rect 21534 19070 21586 19122
rect 21586 19070 21588 19122
rect 21532 19068 21588 19070
rect 20860 18396 20916 18452
rect 20972 17612 21028 17668
rect 20748 17388 20804 17444
rect 22988 28924 23044 28980
rect 23436 31836 23492 31892
rect 23660 31554 23716 31556
rect 23660 31502 23662 31554
rect 23662 31502 23714 31554
rect 23714 31502 23716 31554
rect 23660 31500 23716 31502
rect 23436 31106 23492 31108
rect 23436 31054 23438 31106
rect 23438 31054 23490 31106
rect 23490 31054 23492 31106
rect 23436 31052 23492 31054
rect 23436 30604 23492 30660
rect 23324 30380 23380 30436
rect 23324 29986 23380 29988
rect 23324 29934 23326 29986
rect 23326 29934 23378 29986
rect 23378 29934 23380 29986
rect 23324 29932 23380 29934
rect 23324 27858 23380 27860
rect 23324 27806 23326 27858
rect 23326 27806 23378 27858
rect 23378 27806 23380 27858
rect 23324 27804 23380 27806
rect 22988 27580 23044 27636
rect 23100 27186 23156 27188
rect 23100 27134 23102 27186
rect 23102 27134 23154 27186
rect 23154 27134 23156 27186
rect 23100 27132 23156 27134
rect 22204 26572 22260 26628
rect 22428 26572 22484 26628
rect 22876 26514 22932 26516
rect 22876 26462 22878 26514
rect 22878 26462 22930 26514
rect 22930 26462 22932 26514
rect 22876 26460 22932 26462
rect 22092 25116 22148 25172
rect 22204 23212 22260 23268
rect 22428 23266 22484 23268
rect 22428 23214 22430 23266
rect 22430 23214 22482 23266
rect 22482 23214 22484 23266
rect 22428 23212 22484 23214
rect 22316 23154 22372 23156
rect 22316 23102 22318 23154
rect 22318 23102 22370 23154
rect 22370 23102 22372 23154
rect 22316 23100 22372 23102
rect 22092 20860 22148 20916
rect 22764 24946 22820 24948
rect 22764 24894 22766 24946
rect 22766 24894 22818 24946
rect 22818 24894 22820 24946
rect 22764 24892 22820 24894
rect 22652 24668 22708 24724
rect 23324 27020 23380 27076
rect 23324 26684 23380 26740
rect 23212 24668 23268 24724
rect 22988 23100 23044 23156
rect 23100 24108 23156 24164
rect 22652 21756 22708 21812
rect 22428 21308 22484 21364
rect 22204 20524 22260 20580
rect 22876 22428 22932 22484
rect 23100 21980 23156 22036
rect 22764 20860 22820 20916
rect 22876 20524 22932 20580
rect 22652 20412 22708 20468
rect 22092 19906 22148 19908
rect 22092 19854 22094 19906
rect 22094 19854 22146 19906
rect 22146 19854 22148 19906
rect 22092 19852 22148 19854
rect 21868 19292 21924 19348
rect 21980 18956 22036 19012
rect 21308 18284 21364 18340
rect 21420 18060 21476 18116
rect 21308 17836 21364 17892
rect 21308 17052 21364 17108
rect 20524 16380 20580 16436
rect 20300 15874 20356 15876
rect 20300 15822 20302 15874
rect 20302 15822 20354 15874
rect 20354 15822 20356 15874
rect 20300 15820 20356 15822
rect 20748 16098 20804 16100
rect 20748 16046 20750 16098
rect 20750 16046 20802 16098
rect 20802 16046 20804 16098
rect 20748 16044 20804 16046
rect 20524 15372 20580 15428
rect 21644 17948 21700 18004
rect 21980 17724 22036 17780
rect 21644 17164 21700 17220
rect 21532 16380 21588 16436
rect 22428 19628 22484 19684
rect 22428 19404 22484 19460
rect 22204 17836 22260 17892
rect 22092 17164 22148 17220
rect 22652 18284 22708 18340
rect 22876 18396 22932 18452
rect 22540 17836 22596 17892
rect 22764 17666 22820 17668
rect 22764 17614 22766 17666
rect 22766 17614 22818 17666
rect 22818 17614 22820 17666
rect 22764 17612 22820 17614
rect 23324 24610 23380 24612
rect 23324 24558 23326 24610
rect 23326 24558 23378 24610
rect 23378 24558 23380 24610
rect 23324 24556 23380 24558
rect 23660 29426 23716 29428
rect 23660 29374 23662 29426
rect 23662 29374 23714 29426
rect 23714 29374 23716 29426
rect 23660 29372 23716 29374
rect 23660 28924 23716 28980
rect 23996 31388 24052 31444
rect 23996 31164 24052 31220
rect 23884 30940 23940 30996
rect 24220 31388 24276 31444
rect 24892 31554 24948 31556
rect 24892 31502 24894 31554
rect 24894 31502 24946 31554
rect 24946 31502 24948 31554
rect 24892 31500 24948 31502
rect 24444 31164 24500 31220
rect 25452 31218 25508 31220
rect 25452 31166 25454 31218
rect 25454 31166 25506 31218
rect 25506 31166 25508 31218
rect 25452 31164 25508 31166
rect 25228 31106 25284 31108
rect 25228 31054 25230 31106
rect 25230 31054 25282 31106
rect 25282 31054 25284 31106
rect 25228 31052 25284 31054
rect 23996 29260 24052 29316
rect 25340 30380 25396 30436
rect 24332 28812 24388 28868
rect 25340 29708 25396 29764
rect 24668 29372 24724 29428
rect 24556 28700 24612 28756
rect 23884 28642 23940 28644
rect 23884 28590 23886 28642
rect 23886 28590 23938 28642
rect 23938 28590 23940 28642
rect 23884 28588 23940 28590
rect 24108 28642 24164 28644
rect 24108 28590 24110 28642
rect 24110 28590 24162 28642
rect 24162 28590 24164 28642
rect 24108 28588 24164 28590
rect 24780 28588 24836 28644
rect 25452 28700 25508 28756
rect 23884 28364 23940 28420
rect 23548 27692 23604 27748
rect 23548 27244 23604 27300
rect 23660 27356 23716 27412
rect 23660 27020 23716 27076
rect 23660 26684 23716 26740
rect 23772 27132 23828 27188
rect 24108 27916 24164 27972
rect 23996 27356 24052 27412
rect 24108 27244 24164 27300
rect 23884 26908 23940 26964
rect 24108 26852 24164 26908
rect 23772 25788 23828 25844
rect 23548 25676 23604 25732
rect 23772 24892 23828 24948
rect 23548 23436 23604 23492
rect 23996 24834 24052 24836
rect 23996 24782 23998 24834
rect 23998 24782 24050 24834
rect 24050 24782 24052 24834
rect 23996 24780 24052 24782
rect 23884 23772 23940 23828
rect 23436 23212 23492 23268
rect 23548 22370 23604 22372
rect 23548 22318 23550 22370
rect 23550 22318 23602 22370
rect 23602 22318 23604 22370
rect 23548 22316 23604 22318
rect 23996 23100 24052 23156
rect 23884 22428 23940 22484
rect 24108 22764 24164 22820
rect 24332 27916 24388 27972
rect 25116 27916 25172 27972
rect 25228 27858 25284 27860
rect 25228 27806 25230 27858
rect 25230 27806 25282 27858
rect 25282 27806 25284 27858
rect 25228 27804 25284 27806
rect 25340 27468 25396 27524
rect 24780 27132 24836 27188
rect 24332 24556 24388 24612
rect 25228 26124 25284 26180
rect 24892 25506 24948 25508
rect 24892 25454 24894 25506
rect 24894 25454 24946 25506
rect 24946 25454 24948 25506
rect 24892 25452 24948 25454
rect 24668 25228 24724 25284
rect 25116 25228 25172 25284
rect 24780 24498 24836 24500
rect 24780 24446 24782 24498
rect 24782 24446 24834 24498
rect 24834 24446 24836 24498
rect 24780 24444 24836 24446
rect 24556 23826 24612 23828
rect 24556 23774 24558 23826
rect 24558 23774 24610 23826
rect 24610 23774 24612 23826
rect 24556 23772 24612 23774
rect 24332 23436 24388 23492
rect 24332 23266 24388 23268
rect 24332 23214 24334 23266
rect 24334 23214 24386 23266
rect 24386 23214 24388 23266
rect 24332 23212 24388 23214
rect 24108 22316 24164 22372
rect 24332 22204 24388 22260
rect 23660 22092 23716 22148
rect 23548 21644 23604 21700
rect 23324 20578 23380 20580
rect 23324 20526 23326 20578
rect 23326 20526 23378 20578
rect 23378 20526 23380 20578
rect 23324 20524 23380 20526
rect 23212 19346 23268 19348
rect 23212 19294 23214 19346
rect 23214 19294 23266 19346
rect 23266 19294 23268 19346
rect 23212 19292 23268 19294
rect 23100 18226 23156 18228
rect 23100 18174 23102 18226
rect 23102 18174 23154 18226
rect 23154 18174 23156 18226
rect 23100 18172 23156 18174
rect 22092 16940 22148 16996
rect 21980 16828 22036 16884
rect 22092 16492 22148 16548
rect 21644 15820 21700 15876
rect 21868 16098 21924 16100
rect 21868 16046 21870 16098
rect 21870 16046 21922 16098
rect 21922 16046 21924 16098
rect 21868 16044 21924 16046
rect 22540 16098 22596 16100
rect 22540 16046 22542 16098
rect 22542 16046 22594 16098
rect 22594 16046 22596 16098
rect 22540 16044 22596 16046
rect 22428 15874 22484 15876
rect 22428 15822 22430 15874
rect 22430 15822 22482 15874
rect 22482 15822 22484 15874
rect 22428 15820 22484 15822
rect 22092 15538 22148 15540
rect 22092 15486 22094 15538
rect 22094 15486 22146 15538
rect 22146 15486 22148 15538
rect 22092 15484 22148 15486
rect 20076 14476 20132 14532
rect 22316 15260 22372 15316
rect 19852 14252 19908 14308
rect 21980 14812 22036 14868
rect 20860 14252 20916 14308
rect 22204 14588 22260 14644
rect 21980 14418 22036 14420
rect 21980 14366 21982 14418
rect 21982 14366 22034 14418
rect 22034 14366 22036 14418
rect 21980 14364 22036 14366
rect 21868 14252 21924 14308
rect 19628 14140 19684 14196
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18956 13970 19012 13972
rect 18956 13918 18958 13970
rect 18958 13918 19010 13970
rect 19010 13918 19012 13970
rect 18956 13916 19012 13918
rect 13692 13858 13748 13860
rect 13692 13806 13694 13858
rect 13694 13806 13746 13858
rect 13746 13806 13748 13858
rect 13692 13804 13748 13806
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 8876 11452 8932 11508
rect 22540 14642 22596 14644
rect 22540 14590 22542 14642
rect 22542 14590 22594 14642
rect 22594 14590 22596 14642
rect 22540 14588 22596 14590
rect 22876 17052 22932 17108
rect 22988 17500 23044 17556
rect 22764 15372 22820 15428
rect 22652 14364 22708 14420
rect 23100 16098 23156 16100
rect 23100 16046 23102 16098
rect 23102 16046 23154 16098
rect 23154 16046 23156 16098
rect 23100 16044 23156 16046
rect 23100 15820 23156 15876
rect 23212 15426 23268 15428
rect 23212 15374 23214 15426
rect 23214 15374 23266 15426
rect 23266 15374 23268 15426
rect 23212 15372 23268 15374
rect 24220 21698 24276 21700
rect 24220 21646 24222 21698
rect 24222 21646 24274 21698
rect 24274 21646 24276 21698
rect 24220 21644 24276 21646
rect 23996 21586 24052 21588
rect 23996 21534 23998 21586
rect 23998 21534 24050 21586
rect 24050 21534 24052 21586
rect 23996 21532 24052 21534
rect 24556 21980 24612 22036
rect 23548 18620 23604 18676
rect 23660 19292 23716 19348
rect 25228 24892 25284 24948
rect 25228 24722 25284 24724
rect 25228 24670 25230 24722
rect 25230 24670 25282 24722
rect 25282 24670 25284 24722
rect 25228 24668 25284 24670
rect 26908 32620 26964 32676
rect 26124 28812 26180 28868
rect 25564 27804 25620 27860
rect 25788 25394 25844 25396
rect 25788 25342 25790 25394
rect 25790 25342 25842 25394
rect 25842 25342 25844 25394
rect 25788 25340 25844 25342
rect 26236 28252 26292 28308
rect 26124 27858 26180 27860
rect 26124 27806 26126 27858
rect 26126 27806 26178 27858
rect 26178 27806 26180 27858
rect 26124 27804 26180 27806
rect 26012 27468 26068 27524
rect 26348 27468 26404 27524
rect 26236 27074 26292 27076
rect 26236 27022 26238 27074
rect 26238 27022 26290 27074
rect 26290 27022 26292 27074
rect 26236 27020 26292 27022
rect 28140 28252 28196 28308
rect 27356 27804 27412 27860
rect 26684 26514 26740 26516
rect 26684 26462 26686 26514
rect 26686 26462 26738 26514
rect 26738 26462 26740 26514
rect 26684 26460 26740 26462
rect 26796 26402 26852 26404
rect 26796 26350 26798 26402
rect 26798 26350 26850 26402
rect 26850 26350 26852 26402
rect 26796 26348 26852 26350
rect 26236 26290 26292 26292
rect 26236 26238 26238 26290
rect 26238 26238 26290 26290
rect 26290 26238 26292 26290
rect 26236 26236 26292 26238
rect 27580 26460 27636 26516
rect 28364 27020 28420 27076
rect 27468 26236 27524 26292
rect 26908 24220 26964 24276
rect 25116 22988 25172 23044
rect 25004 21980 25060 22036
rect 23884 20130 23940 20132
rect 23884 20078 23886 20130
rect 23886 20078 23938 20130
rect 23938 20078 23940 20130
rect 23884 20076 23940 20078
rect 24444 20188 24500 20244
rect 24108 19458 24164 19460
rect 24108 19406 24110 19458
rect 24110 19406 24162 19458
rect 24162 19406 24164 19458
rect 24108 19404 24164 19406
rect 23996 19122 24052 19124
rect 23996 19070 23998 19122
rect 23998 19070 24050 19122
rect 24050 19070 24052 19122
rect 23996 19068 24052 19070
rect 23884 18396 23940 18452
rect 23772 15820 23828 15876
rect 23324 15260 23380 15316
rect 24108 18172 24164 18228
rect 24108 17612 24164 17668
rect 25004 19964 25060 20020
rect 27356 25282 27412 25284
rect 27356 25230 27358 25282
rect 27358 25230 27410 25282
rect 27410 25230 27412 25282
rect 27356 25228 27412 25230
rect 27244 24780 27300 24836
rect 27244 24444 27300 24500
rect 27020 23212 27076 23268
rect 24668 19234 24724 19236
rect 24668 19182 24670 19234
rect 24670 19182 24722 19234
rect 24722 19182 24724 19234
rect 24668 19180 24724 19182
rect 25340 22764 25396 22820
rect 25452 22146 25508 22148
rect 25452 22094 25454 22146
rect 25454 22094 25506 22146
rect 25506 22094 25508 22146
rect 25452 22092 25508 22094
rect 25564 21980 25620 22036
rect 28140 24050 28196 24052
rect 28140 23998 28142 24050
rect 28142 23998 28194 24050
rect 28194 23998 28196 24050
rect 28140 23996 28196 23998
rect 27804 23154 27860 23156
rect 27804 23102 27806 23154
rect 27806 23102 27858 23154
rect 27858 23102 27860 23154
rect 27804 23100 27860 23102
rect 26012 22764 26068 22820
rect 26124 22876 26180 22932
rect 25788 21532 25844 21588
rect 25676 20748 25732 20804
rect 26236 21586 26292 21588
rect 26236 21534 26238 21586
rect 26238 21534 26290 21586
rect 26290 21534 26292 21586
rect 26236 21532 26292 21534
rect 25788 20412 25844 20468
rect 26460 22876 26516 22932
rect 26572 22764 26628 22820
rect 28140 23212 28196 23268
rect 28140 22876 28196 22932
rect 27692 21980 27748 22036
rect 26796 21756 26852 21812
rect 27356 21532 27412 21588
rect 26796 20802 26852 20804
rect 26796 20750 26798 20802
rect 26798 20750 26850 20802
rect 26850 20750 26852 20802
rect 26796 20748 26852 20750
rect 28476 26402 28532 26404
rect 28476 26350 28478 26402
rect 28478 26350 28530 26402
rect 28530 26350 28532 26402
rect 28476 26348 28532 26350
rect 28700 23324 28756 23380
rect 28364 22988 28420 23044
rect 28476 22428 28532 22484
rect 30380 29820 30436 29876
rect 30268 25452 30324 25508
rect 28924 22930 28980 22932
rect 28924 22878 28926 22930
rect 28926 22878 28978 22930
rect 28978 22878 28980 22930
rect 28924 22876 28980 22878
rect 28700 20860 28756 20916
rect 26236 19852 26292 19908
rect 27692 20018 27748 20020
rect 27692 19966 27694 20018
rect 27694 19966 27746 20018
rect 27746 19966 27748 20018
rect 27692 19964 27748 19966
rect 29484 19906 29540 19908
rect 29484 19854 29486 19906
rect 29486 19854 29538 19906
rect 29538 19854 29540 19906
rect 29484 19852 29540 19854
rect 26684 19740 26740 19796
rect 24556 18508 24612 18564
rect 24444 17836 24500 17892
rect 25004 18396 25060 18452
rect 25676 17666 25732 17668
rect 25676 17614 25678 17666
rect 25678 17614 25730 17666
rect 25730 17614 25732 17666
rect 25676 17612 25732 17614
rect 24780 16770 24836 16772
rect 24780 16718 24782 16770
rect 24782 16718 24834 16770
rect 24834 16718 24836 16770
rect 24780 16716 24836 16718
rect 32844 26348 32900 26404
rect 34412 37100 34468 37156
rect 35980 37154 36036 37156
rect 35980 37102 35982 37154
rect 35982 37102 36034 37154
rect 36034 37102 36036 37154
rect 35980 37100 36036 37102
rect 36428 37100 36484 37156
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34412 23996 34468 24052
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 30380 20076 30436 20132
rect 37660 19852 37716 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 30268 16716 30324 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 23884 15036 23940 15092
rect 26012 15372 26068 15428
rect 24668 15036 24724 15092
rect 23100 14812 23156 14868
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 22876 11564 22932 11620
rect 22316 11340 22372 11396
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 6300 9212 6356 9268
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4844 7644 4900 7700
rect 4060 7420 4116 7476
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 3724 6300 3780 6356
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 2492 6076 2548 6132
rect 1708 5740 1764 5796
rect 1708 5180 1764 5236
rect 1260 4732 1316 4788
rect 2492 5794 2548 5796
rect 2492 5742 2494 5794
rect 2494 5742 2546 5794
rect 2546 5742 2548 5794
rect 2492 5740 2548 5742
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 1708 4844 1764 4900
rect 2492 4844 2548 4900
rect 1708 4284 1764 4340
rect 2044 4732 2100 4788
rect 1708 3442 1764 3444
rect 1708 3390 1710 3442
rect 1710 3390 1762 3442
rect 1762 3390 1764 3442
rect 1708 3388 1764 3390
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 2492 3442 2548 3444
rect 2492 3390 2494 3442
rect 2494 3390 2546 3442
rect 2546 3390 2548 3442
rect 2492 3388 2548 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
<< metal3 >>
rect 0 38388 800 38416
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 0 38332 3388 38388
rect 0 38304 800 38332
rect 3332 38164 3388 38332
rect 15922 38220 15932 38276
rect 15988 38220 17164 38276
rect 17220 38220 17230 38276
rect 22642 38220 22652 38276
rect 22708 38220 25564 38276
rect 25620 38220 25630 38276
rect 32722 38220 32732 38276
rect 32788 38220 33852 38276
rect 33908 38220 33918 38276
rect 36082 38220 36092 38276
rect 36148 38220 37324 38276
rect 37380 38220 37390 38276
rect 3332 38108 4284 38164
rect 4340 38108 7756 38164
rect 7812 38108 7822 38164
rect 10994 38108 11004 38164
rect 11060 38108 13132 38164
rect 13188 38108 13692 38164
rect 13748 38108 13758 38164
rect 5954 37996 5964 38052
rect 6020 37996 7308 38052
rect 7364 37996 7374 38052
rect 12562 37996 12572 38052
rect 12628 37996 14252 38052
rect 14308 37996 15036 38052
rect 15092 37996 15102 38052
rect 19506 37996 19516 38052
rect 19572 37996 19964 38052
rect 20020 37996 28700 38052
rect 28756 37996 28766 38052
rect 2370 37884 2380 37940
rect 2436 37884 8204 37940
rect 8260 37884 8270 37940
rect 9538 37884 9548 37940
rect 9604 37884 13468 37940
rect 13524 37884 13534 37940
rect 21298 37884 21308 37940
rect 21364 37884 21756 37940
rect 21812 37884 21822 37940
rect 2258 37772 2268 37828
rect 2324 37772 3948 37828
rect 4004 37772 4014 37828
rect 20962 37772 20972 37828
rect 21028 37772 21644 37828
rect 21700 37772 21710 37828
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 6402 37548 6412 37604
rect 6468 37548 9548 37604
rect 9604 37548 9614 37604
rect 0 37492 800 37520
rect 0 37436 2380 37492
rect 2436 37436 2446 37492
rect 6514 37436 6524 37492
rect 6580 37436 8652 37492
rect 8708 37436 13468 37492
rect 13524 37436 14700 37492
rect 14756 37436 14766 37492
rect 26002 37436 26012 37492
rect 26068 37436 27244 37492
rect 27300 37436 27310 37492
rect 0 37408 800 37436
rect 2706 37324 2716 37380
rect 2772 37324 3388 37380
rect 3444 37324 6748 37380
rect 6804 37324 6814 37380
rect 3154 37212 3164 37268
rect 3220 37212 5236 37268
rect 5394 37212 5404 37268
rect 5460 37212 5852 37268
rect 5908 37212 10220 37268
rect 10276 37212 10286 37268
rect 5180 37156 5236 37212
rect 2706 37100 2716 37156
rect 2772 37100 3388 37156
rect 5180 37100 6300 37156
rect 6356 37100 6366 37156
rect 6850 37100 6860 37156
rect 6916 37100 9996 37156
rect 10052 37100 10062 37156
rect 34402 37100 34412 37156
rect 34468 37100 35980 37156
rect 36036 37100 36428 37156
rect 36484 37100 36494 37156
rect 3332 37044 3388 37100
rect 3332 36988 6524 37044
rect 6580 36988 6590 37044
rect 7746 36988 7756 37044
rect 7812 36988 11004 37044
rect 11060 36988 11070 37044
rect 13346 36988 13356 37044
rect 13412 36988 14308 37044
rect 14252 36932 14308 36988
rect 2034 36876 2044 36932
rect 2100 36876 2940 36932
rect 2996 36876 3836 36932
rect 3892 36876 3902 36932
rect 14242 36876 14252 36932
rect 14308 36876 14318 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 12338 36764 12348 36820
rect 12404 36764 15148 36820
rect 15204 36764 15214 36820
rect 3490 36652 3500 36708
rect 3556 36652 4844 36708
rect 4900 36652 11900 36708
rect 11956 36652 11966 36708
rect 14130 36652 14140 36708
rect 14196 36652 15260 36708
rect 15316 36652 15326 36708
rect 0 36596 800 36624
rect 0 36540 1764 36596
rect 4050 36540 4060 36596
rect 4116 36540 5964 36596
rect 6020 36540 6030 36596
rect 6402 36540 6412 36596
rect 6468 36540 7308 36596
rect 7364 36540 12796 36596
rect 12852 36540 15428 36596
rect 0 36512 800 36540
rect 1708 36372 1764 36540
rect 2594 36428 2604 36484
rect 2660 36428 4284 36484
rect 4340 36428 4350 36484
rect 5282 36428 5292 36484
rect 5348 36428 5740 36484
rect 5796 36428 6972 36484
rect 7028 36428 7038 36484
rect 8194 36428 8204 36484
rect 8260 36428 12012 36484
rect 12068 36428 12078 36484
rect 12898 36428 12908 36484
rect 12964 36428 13692 36484
rect 13748 36428 14028 36484
rect 14084 36428 14094 36484
rect 14690 36428 14700 36484
rect 14756 36428 15148 36484
rect 15204 36428 15214 36484
rect 15372 36372 15428 36540
rect 1708 36316 4956 36372
rect 5012 36316 5022 36372
rect 5740 36316 8148 36372
rect 13794 36316 13804 36372
rect 13860 36316 14588 36372
rect 14644 36316 14654 36372
rect 15250 36316 15260 36372
rect 15316 36316 15428 36372
rect 5740 36148 5796 36316
rect 8092 36260 8148 36316
rect 6402 36204 6412 36260
rect 6468 36204 6478 36260
rect 8082 36204 8092 36260
rect 8148 36204 8158 36260
rect 924 36092 2156 36148
rect 2212 36092 5796 36148
rect 0 35700 800 35728
rect 924 35700 980 36092
rect 6412 36036 6468 36204
rect 14242 36092 14252 36148
rect 14308 36092 15596 36148
rect 15652 36092 16044 36148
rect 16100 36092 16110 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 1138 35980 1148 36036
rect 1204 35980 6468 36036
rect 15138 35980 15148 36036
rect 15204 35980 19628 36036
rect 19684 35980 19694 36036
rect 1586 35868 1596 35924
rect 1652 35868 6860 35924
rect 6916 35868 6926 35924
rect 1810 35756 1820 35812
rect 1876 35756 3388 35812
rect 4386 35756 4396 35812
rect 4452 35756 4956 35812
rect 5012 35756 5022 35812
rect 7298 35756 7308 35812
rect 7364 35756 7374 35812
rect 0 35644 980 35700
rect 3332 35700 3388 35756
rect 7308 35700 7364 35756
rect 3332 35644 3948 35700
rect 4004 35644 7364 35700
rect 10994 35644 11004 35700
rect 11060 35644 11788 35700
rect 11844 35644 12572 35700
rect 12628 35644 12638 35700
rect 0 35616 800 35644
rect 1932 35532 2604 35588
rect 2660 35532 3612 35588
rect 3668 35532 3678 35588
rect 6066 35532 6076 35588
rect 6132 35532 17388 35588
rect 17444 35532 17454 35588
rect 0 34804 800 34832
rect 1932 34804 1988 35532
rect 5058 35420 5068 35476
rect 5124 35420 6412 35476
rect 6468 35420 8204 35476
rect 8260 35420 12236 35476
rect 12292 35420 12302 35476
rect 7634 35308 7644 35364
rect 7700 35308 8652 35364
rect 8708 35308 8718 35364
rect 16482 35308 16492 35364
rect 16548 35308 17836 35364
rect 17892 35308 17902 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 8642 34972 8652 35028
rect 8708 34972 10780 35028
rect 10836 34972 14252 35028
rect 14308 34972 14318 35028
rect 2370 34860 2380 34916
rect 2436 34860 2446 34916
rect 8754 34860 8764 34916
rect 8820 34860 16380 34916
rect 16436 34860 16446 34916
rect 0 34748 1988 34804
rect 2380 34804 2436 34860
rect 2380 34748 2828 34804
rect 2884 34748 2894 34804
rect 3332 34748 4844 34804
rect 4900 34748 6524 34804
rect 6580 34748 6590 34804
rect 11778 34748 11788 34804
rect 11844 34748 12908 34804
rect 12964 34748 12974 34804
rect 0 34720 800 34748
rect 3332 34692 3388 34748
rect 2594 34636 2604 34692
rect 2660 34636 3388 34692
rect 3826 34636 3836 34692
rect 3892 34636 4732 34692
rect 4788 34636 4798 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 1922 34412 1932 34468
rect 1988 34412 2268 34468
rect 2324 34412 2334 34468
rect 2930 34412 2940 34468
rect 2996 34412 6188 34468
rect 6244 34412 8204 34468
rect 8260 34412 8270 34468
rect 7858 34300 7868 34356
rect 7924 34300 15148 34356
rect 2258 34188 2268 34244
rect 2324 34188 3388 34244
rect 3444 34188 3454 34244
rect 15092 34132 15148 34300
rect 2034 34076 2044 34132
rect 2100 34076 3052 34132
rect 3108 34076 3118 34132
rect 6290 34076 6300 34132
rect 6356 34076 6366 34132
rect 8418 34076 8428 34132
rect 8484 34076 9772 34132
rect 9828 34076 9838 34132
rect 13906 34076 13916 34132
rect 13972 34076 14700 34132
rect 14756 34076 14766 34132
rect 15092 34076 16044 34132
rect 16100 34076 16492 34132
rect 16548 34076 16558 34132
rect 2818 33964 2828 34020
rect 2884 33964 3164 34020
rect 3220 33964 5628 34020
rect 5684 33964 5694 34020
rect 0 33908 800 33936
rect 6300 33908 6356 34076
rect 12450 33964 12460 34020
rect 12516 33964 13580 34020
rect 13636 33964 13646 34020
rect 15698 33964 15708 34020
rect 15764 33964 19628 34020
rect 19684 33964 21308 34020
rect 21364 33964 21374 34020
rect 0 33852 1596 33908
rect 1652 33852 1662 33908
rect 4274 33852 4284 33908
rect 4340 33852 7868 33908
rect 7924 33852 7934 33908
rect 14130 33852 14140 33908
rect 14196 33852 15148 33908
rect 15204 33852 15214 33908
rect 0 33824 800 33852
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 11442 33628 11452 33684
rect 11508 33628 19404 33684
rect 19460 33628 19470 33684
rect 5842 33516 5852 33572
rect 5908 33516 6748 33572
rect 6804 33516 6814 33572
rect 14018 33516 14028 33572
rect 14084 33516 14252 33572
rect 14308 33516 16268 33572
rect 16324 33516 16334 33572
rect 19954 33516 19964 33572
rect 20020 33516 20972 33572
rect 21028 33516 21038 33572
rect 3490 33404 3500 33460
rect 3556 33404 7084 33460
rect 7140 33404 7150 33460
rect 15586 33404 15596 33460
rect 15652 33404 17052 33460
rect 17108 33404 18060 33460
rect 18116 33404 18126 33460
rect 1820 33292 2156 33348
rect 2212 33292 2222 33348
rect 4946 33292 4956 33348
rect 5012 33292 5628 33348
rect 5684 33292 5694 33348
rect 10098 33292 10108 33348
rect 10164 33292 11788 33348
rect 11844 33292 11854 33348
rect 0 33012 800 33040
rect 1820 33012 1876 33292
rect 2482 33180 2492 33236
rect 2548 33180 6300 33236
rect 6356 33180 6366 33236
rect 9538 33180 9548 33236
rect 9604 33180 10332 33236
rect 10388 33180 10398 33236
rect 11218 33180 11228 33236
rect 11284 33180 11452 33236
rect 11508 33180 11518 33236
rect 15250 33180 15260 33236
rect 15316 33180 19180 33236
rect 19236 33180 19246 33236
rect 2258 33068 2268 33124
rect 2324 33068 2828 33124
rect 2884 33068 2894 33124
rect 5170 33068 5180 33124
rect 5236 33068 10780 33124
rect 10836 33068 13580 33124
rect 13636 33068 13646 33124
rect 15026 33068 15036 33124
rect 15092 33068 15484 33124
rect 15540 33068 15550 33124
rect 15708 33012 15764 33180
rect 16370 33068 16380 33124
rect 16436 33068 17500 33124
rect 17556 33068 18396 33124
rect 18452 33068 18462 33124
rect 0 32956 1876 33012
rect 4274 32956 4284 33012
rect 4340 32956 6860 33012
rect 6916 32956 6926 33012
rect 7746 32956 7756 33012
rect 7812 32956 15764 33012
rect 0 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 12450 32844 12460 32900
rect 12516 32844 17276 32900
rect 17332 32844 18284 32900
rect 18340 32844 18350 32900
rect 3612 32732 4396 32788
rect 4452 32732 4462 32788
rect 13682 32732 13692 32788
rect 13748 32732 15372 32788
rect 15428 32732 15438 32788
rect 16818 32732 16828 32788
rect 16884 32732 19852 32788
rect 19908 32732 19918 32788
rect 3612 32676 3668 32732
rect 2482 32620 2492 32676
rect 2548 32620 3612 32676
rect 3668 32620 3678 32676
rect 11452 32620 16492 32676
rect 16548 32620 17388 32676
rect 17444 32620 17454 32676
rect 18834 32620 18844 32676
rect 18900 32620 26908 32676
rect 26964 32620 26974 32676
rect 11452 32340 11508 32620
rect 14130 32508 14140 32564
rect 14196 32508 15036 32564
rect 15092 32508 15102 32564
rect 19618 32508 19628 32564
rect 19684 32508 21196 32564
rect 21252 32508 21262 32564
rect 14578 32396 14588 32452
rect 14644 32396 15484 32452
rect 15540 32396 15550 32452
rect 18610 32396 18620 32452
rect 18676 32396 18956 32452
rect 19012 32396 19516 32452
rect 19572 32396 20524 32452
rect 20580 32396 20590 32452
rect 8306 32284 8316 32340
rect 8372 32284 10108 32340
rect 10164 32284 11452 32340
rect 11508 32284 11518 32340
rect 16230 32284 16268 32340
rect 16324 32284 16334 32340
rect 19394 32284 19404 32340
rect 19460 32284 20300 32340
rect 20356 32284 20748 32340
rect 20804 32284 20814 32340
rect 6402 32172 6412 32228
rect 6468 32172 9996 32228
rect 10052 32172 10062 32228
rect 11004 32172 16044 32228
rect 16100 32172 16110 32228
rect 0 32116 800 32144
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 0 32060 3948 32116
rect 4004 32060 4014 32116
rect 4956 32060 5292 32116
rect 5348 32060 5358 32116
rect 0 32032 800 32060
rect 4956 32004 5012 32060
rect 11004 32004 11060 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 2258 31948 2268 32004
rect 2324 31948 3276 32004
rect 3332 31948 3342 32004
rect 3714 31948 3724 32004
rect 3780 31948 4732 32004
rect 4788 31948 5012 32004
rect 5170 31948 5180 32004
rect 5236 31948 11004 32004
rect 11060 31948 11070 32004
rect 15586 31948 15596 32004
rect 15652 31948 16268 32004
rect 16324 31948 18284 32004
rect 18340 31948 19740 32004
rect 19796 31948 19806 32004
rect 3490 31836 3500 31892
rect 3556 31836 6524 31892
rect 6580 31836 7868 31892
rect 7924 31836 7934 31892
rect 11106 31836 11116 31892
rect 11172 31836 12348 31892
rect 12404 31836 12796 31892
rect 12852 31836 13244 31892
rect 13300 31836 13310 31892
rect 16034 31836 16044 31892
rect 16100 31836 16940 31892
rect 16996 31836 17006 31892
rect 20066 31836 20076 31892
rect 20132 31836 21308 31892
rect 21364 31836 21374 31892
rect 21970 31836 21980 31892
rect 22036 31836 22540 31892
rect 22596 31836 22606 31892
rect 22754 31836 22764 31892
rect 22820 31836 23436 31892
rect 23492 31836 23502 31892
rect 3378 31724 3388 31780
rect 3444 31724 4844 31780
rect 4900 31724 6636 31780
rect 6692 31724 8876 31780
rect 8932 31724 8942 31780
rect 13010 31724 13020 31780
rect 13076 31724 21532 31780
rect 21588 31724 21598 31780
rect 3826 31612 3836 31668
rect 3892 31612 6188 31668
rect 6244 31612 6254 31668
rect 7074 31612 7084 31668
rect 7140 31612 9380 31668
rect 9538 31612 9548 31668
rect 9604 31612 11228 31668
rect 11284 31612 11294 31668
rect 11452 31612 15148 31668
rect 15204 31612 15372 31668
rect 15428 31612 15438 31668
rect 15586 31612 15596 31668
rect 15652 31612 16380 31668
rect 16436 31612 16446 31668
rect 20626 31612 20636 31668
rect 20692 31612 22316 31668
rect 22372 31612 23100 31668
rect 23156 31612 23166 31668
rect 9324 31556 9380 31612
rect 11452 31556 11508 31612
rect 23436 31556 23492 31836
rect 2594 31500 2604 31556
rect 2660 31500 5628 31556
rect 5684 31500 7868 31556
rect 7924 31500 8540 31556
rect 8596 31500 8606 31556
rect 9324 31500 11508 31556
rect 11666 31500 11676 31556
rect 11732 31500 12012 31556
rect 12068 31500 13356 31556
rect 13412 31500 13422 31556
rect 16034 31500 16044 31556
rect 16100 31500 17500 31556
rect 17556 31500 17948 31556
rect 18004 31500 18014 31556
rect 21970 31500 21980 31556
rect 22036 31500 22652 31556
rect 22708 31500 22718 31556
rect 23436 31500 23660 31556
rect 23716 31500 24892 31556
rect 24948 31500 24958 31556
rect 22652 31444 22708 31500
rect 5954 31388 5964 31444
rect 6020 31388 7420 31444
rect 7476 31388 8316 31444
rect 8372 31388 8382 31444
rect 9986 31388 9996 31444
rect 10052 31388 19684 31444
rect 22652 31388 23996 31444
rect 24052 31388 24220 31444
rect 24276 31388 24286 31444
rect 15026 31276 15036 31332
rect 15092 31276 15148 31332
rect 15204 31276 16604 31332
rect 16660 31276 16670 31332
rect 0 31220 800 31248
rect 19628 31220 19684 31388
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 0 31164 2492 31220
rect 2548 31164 2558 31220
rect 19628 31164 20972 31220
rect 21028 31164 22204 31220
rect 22260 31164 22652 31220
rect 22708 31164 22718 31220
rect 22866 31164 22876 31220
rect 22932 31164 23996 31220
rect 24052 31164 24444 31220
rect 24500 31164 25452 31220
rect 25508 31164 25518 31220
rect 0 31136 800 31164
rect 2034 31052 2044 31108
rect 2100 31052 3612 31108
rect 3668 31052 3678 31108
rect 11330 31052 11340 31108
rect 11396 31052 14140 31108
rect 14196 31052 15148 31108
rect 15204 31052 15214 31108
rect 21298 31052 21308 31108
rect 21364 31052 22428 31108
rect 22484 31052 23100 31108
rect 23156 31052 23166 31108
rect 23426 31052 23436 31108
rect 23492 31052 25228 31108
rect 25284 31052 25294 31108
rect 23100 30996 23156 31052
rect 1698 30940 1708 30996
rect 1764 30940 1932 30996
rect 1988 30940 1998 30996
rect 6850 30940 6860 30996
rect 6916 30940 10220 30996
rect 10276 30940 11452 30996
rect 11508 30940 11518 30996
rect 12338 30940 12348 30996
rect 12404 30940 13692 30996
rect 13748 30940 13758 30996
rect 14700 30940 17052 30996
rect 17108 30940 17118 30996
rect 17602 30940 17612 30996
rect 17668 30940 18620 30996
rect 18676 30940 18686 30996
rect 23100 30940 23884 30996
rect 23940 30940 23950 30996
rect 14700 30884 14756 30940
rect 4722 30828 4732 30884
rect 4788 30828 6524 30884
rect 6580 30828 7532 30884
rect 7588 30828 7598 30884
rect 9874 30828 9884 30884
rect 9940 30828 12516 30884
rect 12898 30828 12908 30884
rect 12964 30828 14700 30884
rect 14756 30828 14766 30884
rect 16706 30828 16716 30884
rect 16772 30828 18396 30884
rect 18452 30828 21084 30884
rect 21140 30828 21150 30884
rect 12460 30772 12516 30828
rect 10210 30716 10220 30772
rect 10276 30716 11116 30772
rect 11172 30716 11182 30772
rect 12460 30716 20524 30772
rect 20580 30716 21980 30772
rect 22036 30716 22046 30772
rect 16370 30604 16380 30660
rect 16436 30604 18396 30660
rect 18452 30604 18462 30660
rect 22978 30604 22988 30660
rect 23044 30604 23436 30660
rect 23492 30604 23502 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 10322 30492 10332 30548
rect 10388 30492 15148 30548
rect 15204 30492 15214 30548
rect 2034 30380 2044 30436
rect 2100 30380 3948 30436
rect 4004 30380 4014 30436
rect 4274 30380 4284 30436
rect 4340 30380 6972 30436
rect 7028 30380 8988 30436
rect 9044 30380 9054 30436
rect 10546 30380 10556 30436
rect 10612 30380 11340 30436
rect 11396 30380 11406 30436
rect 14242 30380 14252 30436
rect 14308 30380 16380 30436
rect 16436 30380 16446 30436
rect 21522 30380 21532 30436
rect 21588 30380 23324 30436
rect 23380 30380 25340 30436
rect 25396 30380 25406 30436
rect 0 30324 800 30352
rect 0 30268 1932 30324
rect 1988 30268 1998 30324
rect 3042 30268 3052 30324
rect 3108 30268 3118 30324
rect 4498 30268 4508 30324
rect 4564 30268 6076 30324
rect 6132 30268 6412 30324
rect 6468 30268 6478 30324
rect 7298 30268 7308 30324
rect 7364 30268 8204 30324
rect 8260 30268 8270 30324
rect 8418 30268 8428 30324
rect 8484 30268 9996 30324
rect 10052 30268 11004 30324
rect 11060 30268 11070 30324
rect 14354 30268 14364 30324
rect 14420 30268 16492 30324
rect 16548 30268 16558 30324
rect 22418 30268 22428 30324
rect 22484 30268 23044 30324
rect 0 30240 800 30268
rect 2818 29932 2828 29988
rect 2884 29932 2894 29988
rect 2828 29876 2884 29932
rect 3052 29876 3108 30268
rect 8204 30212 8260 30268
rect 5170 30156 5180 30212
rect 5236 30156 6636 30212
rect 6692 30156 7868 30212
rect 7924 30156 7934 30212
rect 8204 30156 8652 30212
rect 8708 30156 8718 30212
rect 9090 30156 9100 30212
rect 9156 30156 10444 30212
rect 10500 30156 10510 30212
rect 12422 30156 12460 30212
rect 12516 30156 12526 30212
rect 15362 30156 15372 30212
rect 15428 30156 15932 30212
rect 15988 30156 15998 30212
rect 22988 30100 23044 30268
rect 9426 30044 9436 30100
rect 9492 30044 9884 30100
rect 9940 30044 9950 30100
rect 11890 30044 11900 30100
rect 11956 30044 14700 30100
rect 14756 30044 14766 30100
rect 17164 30044 19852 30100
rect 19908 30044 19918 30100
rect 22978 30044 22988 30100
rect 23044 30044 23054 30100
rect 17164 29988 17220 30044
rect 3602 29932 3612 29988
rect 3668 29932 4844 29988
rect 4900 29932 4910 29988
rect 9314 29932 9324 29988
rect 9380 29932 9548 29988
rect 9604 29932 9614 29988
rect 12226 29932 12236 29988
rect 12292 29932 17220 29988
rect 18834 29932 18844 29988
rect 18900 29932 22316 29988
rect 22372 29932 22382 29988
rect 23314 29932 23324 29988
rect 23380 29932 26908 29988
rect 26852 29876 26908 29932
rect 1698 29820 1708 29876
rect 1764 29820 1774 29876
rect 2594 29820 2604 29876
rect 2660 29820 2884 29876
rect 3042 29820 3052 29876
rect 3108 29820 3118 29876
rect 12534 29820 12572 29876
rect 12628 29820 12638 29876
rect 16034 29820 16044 29876
rect 16100 29820 16492 29876
rect 16548 29820 16558 29876
rect 17826 29820 17836 29876
rect 17892 29820 18004 29876
rect 18946 29820 18956 29876
rect 19012 29820 19404 29876
rect 19460 29820 19470 29876
rect 26852 29820 30380 29876
rect 30436 29820 30446 29876
rect 1708 29652 1764 29820
rect 17948 29764 18004 29820
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 7858 29708 7868 29764
rect 7924 29708 12124 29764
rect 12180 29708 12190 29764
rect 13234 29708 13244 29764
rect 13300 29708 13580 29764
rect 13636 29708 14588 29764
rect 14644 29708 14654 29764
rect 17948 29708 18508 29764
rect 18564 29708 18900 29764
rect 21858 29708 21868 29764
rect 21924 29708 25340 29764
rect 25396 29708 25406 29764
rect 18844 29652 18900 29708
rect 1148 29596 1764 29652
rect 3826 29596 3836 29652
rect 3892 29596 6188 29652
rect 6244 29596 6972 29652
rect 7028 29596 7038 29652
rect 8754 29596 8764 29652
rect 8820 29596 18620 29652
rect 18676 29596 18686 29652
rect 18844 29596 20636 29652
rect 20692 29596 20702 29652
rect 0 29428 800 29456
rect 1148 29428 1204 29596
rect 1362 29484 1372 29540
rect 1428 29484 2044 29540
rect 2100 29484 2110 29540
rect 3332 29484 4956 29540
rect 5012 29484 5022 29540
rect 5170 29484 5180 29540
rect 5236 29484 9772 29540
rect 9828 29484 9838 29540
rect 12786 29484 12796 29540
rect 12852 29484 13692 29540
rect 13748 29484 13758 29540
rect 13906 29484 13916 29540
rect 13972 29484 14924 29540
rect 14980 29484 14990 29540
rect 15922 29484 15932 29540
rect 15988 29484 21028 29540
rect 21382 29484 21420 29540
rect 21476 29484 21486 29540
rect 3332 29428 3388 29484
rect 13692 29428 13748 29484
rect 20972 29428 21028 29484
rect 0 29372 1204 29428
rect 2370 29372 2380 29428
rect 2436 29372 3388 29428
rect 3602 29372 3612 29428
rect 3668 29372 3948 29428
rect 4004 29372 4396 29428
rect 4452 29372 4462 29428
rect 7634 29372 7644 29428
rect 7700 29372 8652 29428
rect 8708 29372 9548 29428
rect 9604 29372 9614 29428
rect 9986 29372 9996 29428
rect 10052 29372 10444 29428
rect 10500 29372 10510 29428
rect 11890 29372 11900 29428
rect 11956 29372 13636 29428
rect 13692 29372 14028 29428
rect 14084 29372 14094 29428
rect 15138 29372 15148 29428
rect 15204 29372 17836 29428
rect 17892 29372 17902 29428
rect 18274 29372 18284 29428
rect 18340 29372 19404 29428
rect 19460 29372 19470 29428
rect 20962 29372 20972 29428
rect 21028 29372 21038 29428
rect 23650 29372 23660 29428
rect 23716 29372 24668 29428
rect 24724 29372 24734 29428
rect 0 29344 800 29372
rect 13580 29316 13636 29372
rect 3490 29260 3500 29316
rect 3556 29260 4172 29316
rect 4228 29260 4238 29316
rect 7746 29260 7756 29316
rect 7812 29260 7822 29316
rect 8306 29260 8316 29316
rect 8372 29260 8876 29316
rect 8932 29260 8942 29316
rect 11218 29260 11228 29316
rect 11284 29260 12012 29316
rect 12068 29260 12078 29316
rect 13206 29260 13244 29316
rect 13300 29260 13310 29316
rect 13570 29260 13580 29316
rect 13636 29260 14588 29316
rect 14644 29260 14654 29316
rect 15092 29260 21868 29316
rect 21924 29260 23996 29316
rect 24052 29260 24062 29316
rect 3490 29036 3500 29092
rect 3556 29036 4284 29092
rect 4340 29036 4350 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 7756 28980 7812 29260
rect 8876 29204 8932 29260
rect 15092 29204 15148 29260
rect 8876 29148 11340 29204
rect 11396 29148 11406 29204
rect 11666 29148 11676 29204
rect 11732 29148 15148 29204
rect 15250 29148 15260 29204
rect 15316 29148 15708 29204
rect 15764 29148 16044 29204
rect 16100 29148 16110 29204
rect 16594 29148 16604 29204
rect 16660 29148 18060 29204
rect 18116 29148 18126 29204
rect 18946 29148 18956 29204
rect 19012 29148 21644 29204
rect 21700 29148 21710 29204
rect 10322 29036 10332 29092
rect 10388 29036 12460 29092
rect 12516 29036 12526 29092
rect 13122 29036 13132 29092
rect 13188 29036 13468 29092
rect 13524 29036 13534 29092
rect 14354 29036 14364 29092
rect 14420 29036 14700 29092
rect 14756 29036 17388 29092
rect 17444 29036 17454 29092
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 7756 28924 16604 28980
rect 16660 28924 16670 28980
rect 17612 28924 22988 28980
rect 23044 28924 23660 28980
rect 23716 28924 23726 28980
rect 17612 28868 17668 28924
rect 8306 28812 8316 28868
rect 8372 28812 12180 28868
rect 13794 28812 13804 28868
rect 13860 28812 17668 28868
rect 17826 28812 17836 28868
rect 17892 28812 18396 28868
rect 18452 28812 18462 28868
rect 18722 28812 18732 28868
rect 18788 28812 19292 28868
rect 19348 28812 19358 28868
rect 24322 28812 24332 28868
rect 24388 28812 26124 28868
rect 26180 28812 26190 28868
rect 5058 28700 5068 28756
rect 5124 28700 6748 28756
rect 6804 28700 7756 28756
rect 7812 28700 8092 28756
rect 8148 28700 10668 28756
rect 10724 28700 10734 28756
rect 10994 28700 11004 28756
rect 11060 28700 11900 28756
rect 11956 28700 11966 28756
rect 12124 28644 12180 28812
rect 12450 28700 12460 28756
rect 12516 28700 15372 28756
rect 15428 28700 15438 28756
rect 18834 28700 18844 28756
rect 18900 28700 21756 28756
rect 21812 28700 21822 28756
rect 24546 28700 24556 28756
rect 24612 28700 25452 28756
rect 25508 28700 25518 28756
rect 3826 28588 3836 28644
rect 3892 28588 4284 28644
rect 4340 28588 5628 28644
rect 5684 28588 5694 28644
rect 9762 28588 9772 28644
rect 9828 28588 11452 28644
rect 11508 28588 11518 28644
rect 12124 28588 13356 28644
rect 13412 28588 13422 28644
rect 17490 28588 17500 28644
rect 17556 28588 20300 28644
rect 20356 28588 20366 28644
rect 22418 28588 22428 28644
rect 22484 28588 23884 28644
rect 23940 28588 23950 28644
rect 24098 28588 24108 28644
rect 24164 28588 24780 28644
rect 24836 28588 24846 28644
rect 0 28532 800 28560
rect 19068 28532 19124 28588
rect 0 28476 1820 28532
rect 1876 28476 2828 28532
rect 2884 28476 2894 28532
rect 5730 28476 5740 28532
rect 5796 28476 6412 28532
rect 6468 28476 6478 28532
rect 7970 28476 7980 28532
rect 8036 28476 11564 28532
rect 11620 28476 11630 28532
rect 14018 28476 14028 28532
rect 14084 28476 15708 28532
rect 15764 28476 15774 28532
rect 16482 28476 16492 28532
rect 16548 28476 17164 28532
rect 17220 28476 17230 28532
rect 18498 28476 18508 28532
rect 18564 28476 18574 28532
rect 19058 28476 19068 28532
rect 19124 28476 19134 28532
rect 19404 28476 20188 28532
rect 20244 28476 20254 28532
rect 0 28448 800 28476
rect 18508 28420 18564 28476
rect 19404 28420 19460 28476
rect 8418 28364 8428 28420
rect 8484 28364 9660 28420
rect 9716 28364 12236 28420
rect 12292 28364 12302 28420
rect 12562 28364 12572 28420
rect 12628 28364 13356 28420
rect 13412 28364 13422 28420
rect 14214 28364 14252 28420
rect 14308 28364 14318 28420
rect 18508 28364 19292 28420
rect 19348 28364 19460 28420
rect 19842 28364 19852 28420
rect 19908 28364 23884 28420
rect 23940 28364 23950 28420
rect 10322 28252 10332 28308
rect 10388 28252 11228 28308
rect 11284 28252 15484 28308
rect 15540 28252 16268 28308
rect 16324 28252 16334 28308
rect 26226 28252 26236 28308
rect 26292 28252 28140 28308
rect 28196 28252 28206 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 13570 28140 13580 28196
rect 13636 28140 14140 28196
rect 14196 28140 18284 28196
rect 18340 28140 18350 28196
rect 8866 28028 8876 28084
rect 8932 28028 12460 28084
rect 12516 28028 20188 28084
rect 20244 28028 20254 28084
rect 1932 27916 2604 27972
rect 2660 27916 3276 27972
rect 3332 27916 3342 27972
rect 4834 27916 4844 27972
rect 4900 27916 6524 27972
rect 6580 27916 6590 27972
rect 13682 27916 13692 27972
rect 13748 27916 14980 27972
rect 19842 27916 19852 27972
rect 19908 27916 20748 27972
rect 20804 27916 20814 27972
rect 22306 27916 22316 27972
rect 22372 27916 24108 27972
rect 24164 27916 24332 27972
rect 24388 27916 24398 27972
rect 25106 27916 25116 27972
rect 25172 27916 25620 27972
rect 0 27636 800 27664
rect 1932 27636 1988 27916
rect 14924 27860 14980 27916
rect 25564 27860 25620 27916
rect 14924 27804 15148 27860
rect 15204 27804 15708 27860
rect 15764 27804 15774 27860
rect 16034 27804 16044 27860
rect 16100 27804 16604 27860
rect 16660 27804 16670 27860
rect 19030 27804 19068 27860
rect 19124 27804 19134 27860
rect 23314 27804 23324 27860
rect 23380 27804 25228 27860
rect 25284 27804 25294 27860
rect 25554 27804 25564 27860
rect 25620 27804 26124 27860
rect 26180 27804 27356 27860
rect 27412 27804 27422 27860
rect 7186 27692 7196 27748
rect 7252 27692 12908 27748
rect 12964 27692 14028 27748
rect 14084 27692 14094 27748
rect 14354 27692 14364 27748
rect 14420 27692 14924 27748
rect 14980 27692 14990 27748
rect 16258 27692 16268 27748
rect 16324 27692 18844 27748
rect 18900 27692 18910 27748
rect 20290 27692 20300 27748
rect 20356 27692 21308 27748
rect 21364 27692 21374 27748
rect 23492 27636 23548 27748
rect 23604 27692 23614 27748
rect 0 27580 1988 27636
rect 15474 27580 15484 27636
rect 15540 27580 22204 27636
rect 22260 27580 22988 27636
rect 23044 27580 23548 27636
rect 0 27552 800 27580
rect 8092 27468 22540 27524
rect 22596 27468 22606 27524
rect 25330 27468 25340 27524
rect 25396 27468 26012 27524
rect 26068 27468 26348 27524
rect 26404 27468 26414 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 8092 27188 8148 27468
rect 13570 27356 13580 27412
rect 13636 27356 18396 27412
rect 18452 27356 18462 27412
rect 19730 27356 19740 27412
rect 19796 27356 21420 27412
rect 21476 27356 21486 27412
rect 10658 27244 10668 27300
rect 10724 27244 11340 27300
rect 11396 27244 15484 27300
rect 15540 27244 15550 27300
rect 15698 27244 15708 27300
rect 15764 27244 16044 27300
rect 16100 27244 16110 27300
rect 17154 27244 17164 27300
rect 17220 27244 18508 27300
rect 18564 27244 18574 27300
rect 21970 27244 21980 27300
rect 22036 27244 22316 27300
rect 22372 27244 22382 27300
rect 22540 27188 22596 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 23650 27356 23660 27412
rect 23716 27356 23996 27412
rect 24052 27356 24062 27412
rect 23538 27244 23548 27300
rect 23604 27244 24108 27300
rect 24164 27244 24174 27300
rect 4946 27132 4956 27188
rect 5012 27132 8092 27188
rect 8148 27132 8158 27188
rect 14018 27132 14028 27188
rect 14084 27132 14812 27188
rect 14868 27132 14878 27188
rect 15026 27132 15036 27188
rect 15092 27132 18396 27188
rect 18452 27132 18462 27188
rect 20290 27132 20300 27188
rect 20356 27132 20636 27188
rect 20692 27132 20702 27188
rect 22540 27132 23100 27188
rect 23156 27132 23772 27188
rect 23828 27132 24780 27188
rect 24836 27132 24846 27188
rect 3154 27020 3164 27076
rect 3220 27020 3836 27076
rect 3892 27020 3902 27076
rect 5058 27020 5068 27076
rect 5124 27020 5740 27076
rect 5796 27020 5806 27076
rect 10658 27020 10668 27076
rect 10724 27020 11228 27076
rect 11284 27020 11294 27076
rect 12786 27020 12796 27076
rect 12852 27020 15148 27076
rect 15204 27020 15214 27076
rect 16706 27020 16716 27076
rect 16772 27020 23324 27076
rect 23380 27020 23390 27076
rect 23650 27020 23660 27076
rect 23716 27020 26236 27076
rect 26292 27020 28364 27076
rect 28420 27020 28430 27076
rect 11778 26908 11788 26964
rect 11844 26908 12852 26964
rect 14476 26908 15932 26964
rect 15988 26908 15998 26964
rect 22278 26908 22316 26964
rect 22372 26908 22382 26964
rect 23874 26908 23884 26964
rect 23940 26908 24164 26964
rect 12786 26852 12796 26908
rect 12852 26852 12862 26908
rect 14476 26852 14532 26908
rect 24098 26852 24108 26908
rect 24164 26852 24174 26908
rect 1698 26796 1708 26852
rect 1764 26796 1774 26852
rect 14466 26796 14476 26852
rect 14532 26796 14542 26852
rect 15138 26796 15148 26852
rect 15204 26796 15540 26852
rect 16482 26796 16492 26852
rect 16548 26796 20244 26852
rect 20402 26796 20412 26852
rect 20468 26796 21644 26852
rect 21700 26796 21710 26852
rect 21942 26796 21980 26852
rect 22036 26796 22046 26852
rect 0 26740 800 26768
rect 1708 26740 1764 26796
rect 15484 26740 15540 26796
rect 20188 26740 20244 26796
rect 0 26684 1764 26740
rect 8978 26684 8988 26740
rect 9044 26684 9436 26740
rect 9492 26684 9502 26740
rect 15474 26684 15484 26740
rect 15540 26684 15550 26740
rect 16930 26684 16940 26740
rect 16996 26684 17612 26740
rect 17668 26684 17678 26740
rect 20188 26684 23324 26740
rect 23380 26684 23660 26740
rect 23716 26684 23726 26740
rect 0 26656 800 26684
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 6626 26572 6636 26628
rect 6692 26572 7308 26628
rect 7364 26572 7374 26628
rect 8418 26572 8428 26628
rect 8484 26572 10780 26628
rect 10836 26572 13020 26628
rect 13076 26572 17276 26628
rect 17332 26572 17342 26628
rect 22166 26572 22204 26628
rect 22260 26572 22270 26628
rect 22418 26572 22428 26628
rect 22484 26572 23548 26628
rect 2258 26460 2268 26516
rect 2324 26460 2604 26516
rect 2660 26460 3276 26516
rect 3332 26460 3342 26516
rect 9286 26460 9324 26516
rect 9380 26460 9390 26516
rect 12114 26460 12124 26516
rect 12180 26460 13580 26516
rect 13636 26460 13646 26516
rect 14242 26460 14252 26516
rect 14308 26460 17388 26516
rect 17444 26460 17454 26516
rect 19618 26460 19628 26516
rect 19684 26460 19852 26516
rect 19908 26460 19918 26516
rect 21522 26460 21532 26516
rect 21588 26460 22876 26516
rect 22932 26460 22942 26516
rect 23492 26404 23548 26572
rect 26674 26460 26684 26516
rect 26740 26460 27580 26516
rect 27636 26460 27646 26516
rect 7186 26348 7196 26404
rect 7252 26348 7262 26404
rect 9986 26348 9996 26404
rect 10052 26348 13244 26404
rect 13300 26348 13310 26404
rect 13458 26348 13468 26404
rect 13524 26348 15372 26404
rect 15428 26348 16492 26404
rect 16548 26348 16558 26404
rect 19254 26348 19292 26404
rect 19348 26348 19358 26404
rect 23492 26348 26796 26404
rect 26852 26348 26862 26404
rect 28466 26348 28476 26404
rect 28532 26348 32844 26404
rect 32900 26348 32910 26404
rect 7196 26292 7252 26348
rect 2594 26236 2604 26292
rect 2660 26236 7252 26292
rect 11554 26236 11564 26292
rect 11620 26236 13132 26292
rect 13188 26236 15596 26292
rect 15652 26236 15662 26292
rect 18274 26236 18284 26292
rect 18340 26236 18732 26292
rect 18788 26236 18798 26292
rect 18946 26236 18956 26292
rect 19012 26236 19516 26292
rect 19572 26236 19582 26292
rect 21074 26236 21084 26292
rect 21140 26236 26236 26292
rect 26292 26236 27468 26292
rect 27524 26236 27534 26292
rect 3378 26124 3388 26180
rect 3444 26124 4060 26180
rect 4116 26124 5964 26180
rect 6020 26124 6030 26180
rect 8082 26124 8092 26180
rect 8148 26124 9548 26180
rect 9604 26124 9614 26180
rect 10994 26124 11004 26180
rect 11060 26124 13580 26180
rect 13636 26124 13646 26180
rect 17938 26124 17948 26180
rect 18004 26124 18620 26180
rect 18676 26124 18686 26180
rect 19506 26124 19516 26180
rect 19572 26124 25228 26180
rect 25284 26124 25294 26180
rect 10770 26012 10780 26068
rect 10836 26012 14476 26068
rect 14532 26012 15148 26068
rect 17602 26012 17612 26068
rect 17668 26012 18732 26068
rect 18788 26012 18798 26068
rect 19394 26012 19404 26068
rect 19460 26012 19628 26068
rect 19684 26012 19694 26068
rect 15092 25956 15148 26012
rect 15092 25900 18060 25956
rect 18116 25900 18126 25956
rect 18274 25900 18284 25956
rect 18340 25900 20412 25956
rect 20468 25900 20478 25956
rect 21270 25900 21308 25956
rect 21364 25900 21374 25956
rect 21606 25900 21644 25956
rect 21700 25900 21710 25956
rect 0 25844 800 25872
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 0 25788 2380 25844
rect 2436 25788 2446 25844
rect 12908 25788 23772 25844
rect 23828 25788 23838 25844
rect 0 25760 800 25788
rect 10966 25676 11004 25732
rect 11060 25676 11070 25732
rect 12908 25620 12964 25788
rect 13570 25676 13580 25732
rect 13636 25676 15988 25732
rect 17378 25676 17388 25732
rect 17444 25676 23548 25732
rect 23604 25676 23614 25732
rect 2146 25564 2156 25620
rect 2212 25564 4508 25620
rect 4564 25564 4574 25620
rect 5058 25564 5068 25620
rect 5124 25564 5852 25620
rect 5908 25564 5918 25620
rect 12898 25564 12908 25620
rect 12964 25564 12974 25620
rect 15932 25508 15988 25676
rect 18834 25564 18844 25620
rect 18900 25564 19516 25620
rect 19572 25564 19582 25620
rect 19954 25564 19964 25620
rect 20020 25564 20636 25620
rect 20692 25564 20702 25620
rect 4610 25452 4620 25508
rect 4676 25452 6188 25508
rect 6244 25452 6254 25508
rect 7298 25452 7308 25508
rect 7364 25452 11788 25508
rect 11844 25452 11854 25508
rect 14018 25452 14028 25508
rect 14084 25452 14812 25508
rect 14868 25452 14878 25508
rect 15922 25452 15932 25508
rect 15988 25452 15998 25508
rect 17042 25452 17052 25508
rect 17108 25452 18508 25508
rect 18564 25452 19796 25508
rect 20514 25452 20524 25508
rect 20580 25452 20972 25508
rect 21028 25452 21038 25508
rect 24882 25452 24892 25508
rect 24948 25452 30268 25508
rect 30324 25452 30334 25508
rect 19740 25396 19796 25452
rect 4498 25340 4508 25396
rect 4564 25340 5516 25396
rect 5572 25340 5582 25396
rect 6514 25340 6524 25396
rect 6580 25340 17836 25396
rect 17892 25340 19180 25396
rect 19236 25340 19246 25396
rect 19730 25340 19740 25396
rect 19796 25340 19806 25396
rect 19954 25340 19964 25396
rect 20020 25340 20188 25396
rect 20244 25340 20412 25396
rect 20468 25340 20478 25396
rect 21410 25340 21420 25396
rect 21476 25340 25788 25396
rect 25844 25340 25854 25396
rect 2034 25228 2044 25284
rect 2100 25228 3220 25284
rect 3378 25228 3388 25284
rect 3444 25228 5292 25284
rect 5348 25228 5358 25284
rect 6626 25228 6636 25284
rect 6692 25228 7420 25284
rect 7476 25228 7756 25284
rect 7812 25228 7822 25284
rect 9090 25228 9100 25284
rect 9156 25228 9996 25284
rect 10052 25228 10062 25284
rect 13458 25228 13468 25284
rect 13524 25228 15372 25284
rect 15428 25228 15438 25284
rect 16940 25228 19404 25284
rect 19460 25228 19470 25284
rect 19628 25228 20244 25284
rect 20738 25228 20748 25284
rect 20804 25228 21308 25284
rect 21364 25228 21374 25284
rect 24658 25228 24668 25284
rect 24724 25228 25116 25284
rect 25172 25228 27356 25284
rect 27412 25228 27422 25284
rect 3164 25060 3220 25228
rect 16940 25172 16996 25228
rect 12898 25116 12908 25172
rect 12964 25116 13356 25172
rect 13412 25116 13422 25172
rect 16930 25116 16940 25172
rect 16996 25116 17006 25172
rect 17490 25116 17500 25172
rect 17556 25116 19180 25172
rect 19236 25116 19246 25172
rect 19628 25060 19684 25228
rect 20188 25172 20244 25228
rect 20188 25116 22092 25172
rect 22148 25116 22158 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 3154 25004 3164 25060
rect 3220 25004 3230 25060
rect 8642 25004 8652 25060
rect 8708 25004 9884 25060
rect 9940 25004 9950 25060
rect 11676 25004 17276 25060
rect 17332 25004 18284 25060
rect 18340 25004 18350 25060
rect 18498 25004 18508 25060
rect 18564 25004 19684 25060
rect 0 24948 800 24976
rect 11676 24948 11732 25004
rect 0 24892 1820 24948
rect 1876 24892 1886 24948
rect 4022 24892 4060 24948
rect 4116 24892 4126 24948
rect 4946 24892 4956 24948
rect 5012 24892 5628 24948
rect 5684 24892 5694 24948
rect 8866 24892 8876 24948
rect 8932 24892 11676 24948
rect 11732 24892 11742 24948
rect 14578 24892 14588 24948
rect 14644 24892 15372 24948
rect 15428 24892 15438 24948
rect 16230 24892 16268 24948
rect 16324 24892 16334 24948
rect 17724 24892 22764 24948
rect 22820 24892 23772 24948
rect 23828 24892 25228 24948
rect 25284 24892 25294 24948
rect 0 24864 800 24892
rect 17724 24836 17780 24892
rect 5058 24780 5068 24836
rect 5124 24780 6076 24836
rect 6132 24780 6412 24836
rect 6468 24780 6478 24836
rect 17686 24780 17724 24836
rect 17780 24780 17790 24836
rect 18050 24780 18060 24836
rect 18116 24780 18956 24836
rect 19012 24780 19022 24836
rect 19170 24780 19180 24836
rect 19236 24780 19274 24836
rect 23986 24780 23996 24836
rect 24052 24780 27244 24836
rect 27300 24780 27310 24836
rect 4162 24668 4172 24724
rect 4228 24668 5852 24724
rect 5908 24668 7532 24724
rect 7588 24668 7598 24724
rect 8306 24668 8316 24724
rect 8372 24668 10668 24724
rect 10724 24668 10734 24724
rect 13234 24668 13244 24724
rect 13300 24668 14252 24724
rect 14308 24668 18284 24724
rect 18340 24668 18508 24724
rect 18564 24668 18574 24724
rect 22642 24668 22652 24724
rect 22708 24668 23212 24724
rect 23268 24668 25228 24724
rect 25284 24668 25294 24724
rect 7410 24556 7420 24612
rect 7476 24556 8764 24612
rect 8820 24556 8830 24612
rect 14018 24556 14028 24612
rect 14084 24556 15148 24612
rect 17490 24556 17500 24612
rect 17556 24556 18396 24612
rect 18452 24556 18462 24612
rect 18722 24556 18732 24612
rect 18788 24556 19180 24612
rect 19236 24556 19964 24612
rect 20020 24556 20030 24612
rect 23314 24556 23324 24612
rect 23380 24556 24332 24612
rect 24388 24556 24398 24612
rect 3602 24444 3612 24500
rect 3668 24444 4060 24500
rect 4116 24444 4126 24500
rect 4610 24444 4620 24500
rect 4676 24444 4844 24500
rect 4900 24444 4910 24500
rect 7634 24444 7644 24500
rect 7700 24444 12684 24500
rect 12740 24444 12750 24500
rect 8082 24332 8092 24388
rect 8148 24332 10220 24388
rect 10276 24332 12348 24388
rect 12404 24332 12414 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 15092 24276 15148 24556
rect 18498 24444 18508 24500
rect 18564 24444 18620 24500
rect 18676 24444 19404 24500
rect 19460 24444 20412 24500
rect 20468 24444 20478 24500
rect 24770 24444 24780 24500
rect 24836 24444 27244 24500
rect 27300 24444 27310 24500
rect 15810 24332 15820 24388
rect 15876 24332 20188 24388
rect 20244 24332 20254 24388
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 9202 24220 9212 24276
rect 9268 24220 9996 24276
rect 10052 24220 10062 24276
rect 15092 24220 26908 24276
rect 26964 24220 26974 24276
rect 3490 24108 3500 24164
rect 3556 24108 3948 24164
rect 4004 24108 4014 24164
rect 10770 24108 10780 24164
rect 10836 24108 23100 24164
rect 23156 24108 23166 24164
rect 0 24052 800 24080
rect 0 23996 1708 24052
rect 1764 23996 2940 24052
rect 2996 23996 3006 24052
rect 7858 23996 7868 24052
rect 7924 23996 14924 24052
rect 14980 23996 14990 24052
rect 17490 23996 17500 24052
rect 17556 23996 21868 24052
rect 21924 23996 21934 24052
rect 28130 23996 28140 24052
rect 28196 23996 34412 24052
rect 34468 23996 34478 24052
rect 0 23968 800 23996
rect 3938 23884 3948 23940
rect 4004 23884 8428 23940
rect 8484 23884 8494 23940
rect 11190 23884 11228 23940
rect 11284 23884 11294 23940
rect 12674 23884 12684 23940
rect 12740 23884 14140 23940
rect 14196 23884 14206 23940
rect 14690 23884 14700 23940
rect 14756 23884 15148 23940
rect 16146 23884 16156 23940
rect 16212 23884 20300 23940
rect 20356 23884 21308 23940
rect 21364 23884 21374 23940
rect 15092 23828 15148 23884
rect 4162 23772 4172 23828
rect 4228 23772 4620 23828
rect 4676 23772 5628 23828
rect 5684 23772 5694 23828
rect 6636 23772 13468 23828
rect 13524 23772 13534 23828
rect 15092 23772 16380 23828
rect 16436 23772 16446 23828
rect 17612 23772 19628 23828
rect 19684 23772 21196 23828
rect 21252 23772 21262 23828
rect 23874 23772 23884 23828
rect 23940 23772 24556 23828
rect 24612 23772 24622 23828
rect 6636 23716 6692 23772
rect 17612 23716 17668 23772
rect 4050 23660 4060 23716
rect 4116 23660 4732 23716
rect 4788 23660 4798 23716
rect 6626 23660 6636 23716
rect 6692 23660 6702 23716
rect 6962 23660 6972 23716
rect 7028 23660 17668 23716
rect 18722 23660 18732 23716
rect 18788 23660 20412 23716
rect 20468 23660 20478 23716
rect 21382 23660 21420 23716
rect 21476 23660 21486 23716
rect 4806 23548 4844 23604
rect 4900 23548 4910 23604
rect 10210 23548 10220 23604
rect 10276 23548 13244 23604
rect 13300 23548 13310 23604
rect 14130 23548 14140 23604
rect 14196 23548 17388 23604
rect 17444 23548 17454 23604
rect 18470 23548 18508 23604
rect 18564 23548 18574 23604
rect 18834 23548 18844 23604
rect 18900 23548 18956 23604
rect 19012 23548 19022 23604
rect 19170 23548 19180 23604
rect 19236 23548 19274 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 5954 23436 5964 23492
rect 6020 23436 9884 23492
rect 9940 23436 10444 23492
rect 10500 23436 10510 23492
rect 10994 23436 11004 23492
rect 11060 23436 11452 23492
rect 11508 23436 11518 23492
rect 16902 23436 16940 23492
rect 16996 23436 17006 23492
rect 17154 23436 17164 23492
rect 17220 23436 17500 23492
rect 17556 23436 17566 23492
rect 18050 23436 18060 23492
rect 18116 23436 19684 23492
rect 23538 23436 23548 23492
rect 23604 23436 24332 23492
rect 24388 23436 24398 23492
rect 19628 23380 19684 23436
rect 2706 23324 2716 23380
rect 2772 23324 3612 23380
rect 3668 23324 3678 23380
rect 6850 23324 6860 23380
rect 6916 23324 8204 23380
rect 8260 23324 8270 23380
rect 9426 23324 9436 23380
rect 9492 23324 9502 23380
rect 10770 23324 10780 23380
rect 10836 23324 11116 23380
rect 11172 23324 11182 23380
rect 16594 23324 16604 23380
rect 16660 23324 19068 23380
rect 19124 23324 19134 23380
rect 19618 23324 19628 23380
rect 19684 23324 19694 23380
rect 22204 23324 28700 23380
rect 28756 23324 28766 23380
rect 9436 23268 9492 23324
rect 22204 23268 22260 23324
rect 6402 23212 6412 23268
rect 6468 23212 9492 23268
rect 10182 23212 10220 23268
rect 10276 23212 10286 23268
rect 11116 23212 18396 23268
rect 18452 23212 19516 23268
rect 19572 23212 19582 23268
rect 22194 23212 22204 23268
rect 22260 23212 22270 23268
rect 22418 23212 22428 23268
rect 22484 23212 23436 23268
rect 23492 23212 23502 23268
rect 24322 23212 24332 23268
rect 24388 23212 27020 23268
rect 27076 23212 28140 23268
rect 28196 23212 28206 23268
rect 0 23156 800 23184
rect 0 23100 1932 23156
rect 1988 23100 1998 23156
rect 4946 23100 4956 23156
rect 5012 23100 7756 23156
rect 7812 23100 7822 23156
rect 9090 23100 9100 23156
rect 9156 23100 9660 23156
rect 9716 23100 9726 23156
rect 0 23072 800 23100
rect 11116 23044 11172 23212
rect 11330 23100 11340 23156
rect 11396 23100 14476 23156
rect 14532 23100 14542 23156
rect 14914 23100 14924 23156
rect 14980 23100 20860 23156
rect 20916 23100 20926 23156
rect 22306 23100 22316 23156
rect 22372 23100 22988 23156
rect 23044 23100 23054 23156
rect 23986 23100 23996 23156
rect 24052 23100 27804 23156
rect 27860 23100 27870 23156
rect 7410 22988 7420 23044
rect 7476 22988 8876 23044
rect 8932 22988 8942 23044
rect 11106 22988 11116 23044
rect 11172 22988 11182 23044
rect 12348 22988 17948 23044
rect 18004 22988 18014 23044
rect 18722 22988 18732 23044
rect 18788 22988 19404 23044
rect 19460 22988 19470 23044
rect 25106 22988 25116 23044
rect 25172 22988 28364 23044
rect 28420 22988 28430 23044
rect 8082 22876 8092 22932
rect 8148 22876 9772 22932
rect 9828 22876 11228 22932
rect 11284 22876 12124 22932
rect 12180 22876 12190 22932
rect 12348 22820 12404 22988
rect 13234 22876 13244 22932
rect 13300 22876 17164 22932
rect 17220 22876 17230 22932
rect 17826 22876 17836 22932
rect 17892 22876 18284 22932
rect 18340 22876 18350 22932
rect 18946 22876 18956 22932
rect 19012 22876 26124 22932
rect 26180 22876 26460 22932
rect 26516 22876 26526 22932
rect 28130 22876 28140 22932
rect 28196 22876 28924 22932
rect 28980 22876 28990 22932
rect 5058 22764 5068 22820
rect 5124 22764 6076 22820
rect 6132 22764 8540 22820
rect 8596 22764 8606 22820
rect 8866 22764 8876 22820
rect 8932 22764 12404 22820
rect 12562 22764 12572 22820
rect 12628 22764 12908 22820
rect 12964 22764 12974 22820
rect 16706 22764 16716 22820
rect 16772 22764 23548 22820
rect 24098 22764 24108 22820
rect 24164 22764 25340 22820
rect 25396 22764 25406 22820
rect 26002 22764 26012 22820
rect 26068 22764 26572 22820
rect 26628 22764 26638 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 7522 22652 7532 22708
rect 7588 22652 21868 22708
rect 21924 22652 21934 22708
rect 3378 22540 3388 22596
rect 3444 22540 3482 22596
rect 15670 22540 15708 22596
rect 15764 22540 15774 22596
rect 17042 22540 17052 22596
rect 17108 22540 17500 22596
rect 17556 22540 17566 22596
rect 18722 22540 18732 22596
rect 18788 22540 20076 22596
rect 20132 22540 20142 22596
rect 23492 22484 23548 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 4162 22428 4172 22484
rect 4228 22428 6972 22484
rect 7028 22428 7038 22484
rect 10994 22428 11004 22484
rect 11060 22428 13580 22484
rect 13636 22428 13646 22484
rect 13794 22428 13804 22484
rect 13860 22428 14364 22484
rect 14420 22428 14430 22484
rect 15810 22428 15820 22484
rect 15876 22428 16044 22484
rect 16100 22428 16492 22484
rect 16548 22428 16558 22484
rect 18162 22428 18172 22484
rect 18228 22428 18508 22484
rect 18564 22428 18574 22484
rect 19590 22428 19628 22484
rect 19684 22428 19694 22484
rect 20626 22428 20636 22484
rect 20692 22428 22876 22484
rect 22932 22428 22942 22484
rect 23492 22428 23884 22484
rect 23940 22428 24220 22484
rect 24276 22428 28476 22484
rect 28532 22428 28542 22484
rect 1810 22316 1820 22372
rect 1876 22316 1886 22372
rect 2370 22316 2380 22372
rect 2436 22316 2940 22372
rect 2996 22316 4284 22372
rect 4340 22316 4350 22372
rect 5730 22316 5740 22372
rect 5796 22316 6412 22372
rect 6468 22316 6478 22372
rect 8978 22316 8988 22372
rect 9044 22316 16156 22372
rect 16212 22316 16222 22372
rect 16818 22316 16828 22372
rect 16884 22316 17164 22372
rect 17220 22316 17230 22372
rect 17490 22316 17500 22372
rect 17556 22316 23548 22372
rect 23604 22316 23614 22372
rect 24070 22316 24108 22372
rect 24164 22316 24174 22372
rect 0 22260 800 22288
rect 1820 22260 1876 22316
rect 23548 22260 23604 22316
rect 0 22204 1876 22260
rect 3686 22204 3724 22260
rect 3780 22204 3790 22260
rect 12450 22204 12460 22260
rect 12516 22204 15372 22260
rect 15428 22204 17724 22260
rect 17780 22204 17790 22260
rect 23548 22204 24332 22260
rect 24388 22204 24398 22260
rect 0 22176 800 22204
rect 2034 22092 2044 22148
rect 2100 22092 4172 22148
rect 4228 22092 4238 22148
rect 4834 22092 4844 22148
rect 4900 22092 5740 22148
rect 5796 22092 5806 22148
rect 10098 22092 10108 22148
rect 10164 22092 11004 22148
rect 11060 22092 11564 22148
rect 11620 22092 14812 22148
rect 14868 22092 14878 22148
rect 16818 22092 16828 22148
rect 16884 22092 18508 22148
rect 18564 22092 19292 22148
rect 19348 22092 19358 22148
rect 19842 22092 19852 22148
rect 19908 22092 20188 22148
rect 20244 22092 20254 22148
rect 23650 22092 23660 22148
rect 23716 22092 25452 22148
rect 25508 22092 25518 22148
rect 3938 21980 3948 22036
rect 4004 21980 5516 22036
rect 5572 21980 5582 22036
rect 10630 21980 10668 22036
rect 10724 21980 10734 22036
rect 16930 21980 16940 22036
rect 16996 21980 19348 22036
rect 20738 21980 20748 22036
rect 20804 21980 21084 22036
rect 21140 21980 21150 22036
rect 23090 21980 23100 22036
rect 23156 21980 24556 22036
rect 24612 21980 25004 22036
rect 25060 21980 25564 22036
rect 25620 21980 27692 22036
rect 27748 21980 27758 22036
rect 2370 21868 2380 21924
rect 2436 21868 7308 21924
rect 7364 21868 7374 21924
rect 12898 21868 12908 21924
rect 12964 21868 13244 21924
rect 13300 21868 13310 21924
rect 13906 21868 13916 21924
rect 13972 21868 17612 21924
rect 17668 21868 17678 21924
rect 3826 21756 3836 21812
rect 3892 21756 4060 21812
rect 4116 21756 4126 21812
rect 4722 21756 4732 21812
rect 4788 21756 6188 21812
rect 6244 21756 6254 21812
rect 8278 21756 8316 21812
rect 8372 21756 8382 21812
rect 11666 21756 11676 21812
rect 11732 21756 12460 21812
rect 12516 21756 12526 21812
rect 16258 21756 16268 21812
rect 16324 21756 18844 21812
rect 18900 21756 18910 21812
rect 19292 21700 19348 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 20822 21868 20860 21924
rect 20916 21868 20926 21924
rect 19506 21756 19516 21812
rect 19572 21756 21420 21812
rect 21476 21756 21486 21812
rect 21718 21756 21756 21812
rect 21812 21756 21822 21812
rect 22642 21756 22652 21812
rect 22708 21756 26796 21812
rect 26852 21756 26862 21812
rect 2034 21644 2044 21700
rect 2100 21644 4844 21700
rect 4900 21644 5852 21700
rect 5908 21644 5918 21700
rect 12114 21644 12124 21700
rect 12180 21644 13580 21700
rect 13636 21644 13646 21700
rect 14018 21644 14028 21700
rect 14084 21644 15708 21700
rect 15764 21644 15774 21700
rect 18946 21644 18956 21700
rect 19012 21644 20860 21700
rect 20916 21644 20926 21700
rect 21298 21644 21308 21700
rect 21364 21644 23548 21700
rect 23604 21644 23614 21700
rect 24182 21644 24220 21700
rect 24276 21644 24286 21700
rect 13580 21588 13636 21644
rect 2818 21532 2828 21588
rect 2884 21532 3164 21588
rect 3220 21532 3230 21588
rect 3378 21532 3388 21588
rect 3444 21532 4284 21588
rect 4340 21532 4350 21588
rect 7186 21532 7196 21588
rect 7252 21532 8652 21588
rect 8708 21532 9660 21588
rect 9716 21532 9726 21588
rect 10546 21532 10556 21588
rect 10612 21532 12572 21588
rect 12628 21532 13524 21588
rect 13580 21532 14140 21588
rect 14196 21532 17388 21588
rect 17444 21532 17454 21588
rect 17826 21532 17836 21588
rect 17892 21532 19404 21588
rect 19460 21532 19470 21588
rect 23986 21532 23996 21588
rect 24052 21532 24062 21588
rect 25778 21532 25788 21588
rect 25844 21532 26236 21588
rect 26292 21532 27356 21588
rect 27412 21532 27422 21588
rect 13468 21476 13524 21532
rect 23996 21476 24052 21532
rect 2258 21420 2268 21476
rect 2324 21420 2716 21476
rect 2772 21420 2782 21476
rect 6626 21420 6636 21476
rect 6692 21420 12124 21476
rect 12180 21420 12190 21476
rect 13468 21420 14532 21476
rect 0 21364 800 21392
rect 0 21308 1596 21364
rect 1652 21308 1662 21364
rect 11218 21308 11228 21364
rect 11284 21308 11564 21364
rect 11620 21308 13804 21364
rect 13860 21308 13870 21364
rect 0 21280 800 21308
rect 12786 21196 12796 21252
rect 12852 21196 14028 21252
rect 14084 21196 14094 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 5142 21084 5180 21140
rect 5236 21084 5246 21140
rect 7298 21084 7308 21140
rect 7364 21084 13860 21140
rect 3826 20972 3836 21028
rect 3892 20972 6412 21028
rect 6468 20972 6478 21028
rect 11190 20972 11228 21028
rect 11284 20972 11294 21028
rect 13570 20972 13580 21028
rect 13636 20972 13646 21028
rect 2370 20860 2380 20916
rect 2436 20860 2940 20916
rect 2996 20860 3006 20916
rect 3266 20860 3276 20916
rect 3332 20860 7756 20916
rect 7812 20860 7822 20916
rect 13580 20804 13636 20972
rect 13804 20916 13860 21084
rect 14476 21028 14532 21420
rect 15932 21420 24052 21476
rect 15932 21364 15988 21420
rect 15922 21308 15932 21364
rect 15988 21308 15998 21364
rect 16370 21308 16380 21364
rect 16436 21308 16828 21364
rect 16884 21308 17388 21364
rect 17444 21308 17454 21364
rect 17938 21308 17948 21364
rect 18004 21308 22428 21364
rect 22484 21308 22494 21364
rect 16380 21140 16436 21308
rect 21270 21196 21308 21252
rect 21364 21196 21374 21252
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 14690 21084 14700 21140
rect 14756 21084 16436 21140
rect 20402 21084 20412 21140
rect 20468 21084 21084 21140
rect 21140 21084 21150 21140
rect 14476 20972 20580 21028
rect 20738 20972 20748 21028
rect 20804 20972 21700 21028
rect 20524 20916 20580 20972
rect 21644 20916 21700 20972
rect 13804 20860 14364 20916
rect 14420 20860 14700 20916
rect 14756 20860 14766 20916
rect 20514 20860 20524 20916
rect 20580 20860 21420 20916
rect 21476 20860 21486 20916
rect 21634 20860 21644 20916
rect 21700 20860 21710 20916
rect 22082 20860 22092 20916
rect 22148 20860 22764 20916
rect 22820 20860 28700 20916
rect 28756 20860 28766 20916
rect 1250 20748 1260 20804
rect 1316 20748 2436 20804
rect 3042 20748 3052 20804
rect 3108 20748 8204 20804
rect 8260 20748 8270 20804
rect 13580 20748 15148 20804
rect 15204 20748 15214 20804
rect 15698 20748 15708 20804
rect 15764 20748 16156 20804
rect 16212 20748 16222 20804
rect 17154 20748 17164 20804
rect 17220 20748 19292 20804
rect 19348 20748 19358 20804
rect 25666 20748 25676 20804
rect 25732 20748 26796 20804
rect 26852 20748 26862 20804
rect 2380 20692 2436 20748
rect 1698 20636 1708 20692
rect 1764 20636 1774 20692
rect 2380 20636 5180 20692
rect 5236 20636 5852 20692
rect 5908 20636 5918 20692
rect 13458 20636 13468 20692
rect 13524 20636 21868 20692
rect 21924 20636 21934 20692
rect 1708 20580 1764 20636
rect 1708 20524 3164 20580
rect 3220 20524 3230 20580
rect 3378 20524 3388 20580
rect 3444 20524 3724 20580
rect 3780 20524 3790 20580
rect 9762 20524 9772 20580
rect 9828 20524 10444 20580
rect 10500 20524 10510 20580
rect 10770 20524 10780 20580
rect 10836 20524 15148 20580
rect 16566 20524 16604 20580
rect 16660 20524 16670 20580
rect 16930 20524 16940 20580
rect 16996 20524 22204 20580
rect 22260 20524 22270 20580
rect 22866 20524 22876 20580
rect 22932 20524 23324 20580
rect 23380 20524 23390 20580
rect 0 20468 800 20496
rect 15092 20468 15148 20524
rect 0 20412 1708 20468
rect 1764 20412 1774 20468
rect 10210 20412 10220 20468
rect 10276 20412 13860 20468
rect 15092 20412 17836 20468
rect 17892 20412 17902 20468
rect 19394 20412 19404 20468
rect 19460 20412 19628 20468
rect 19684 20412 19694 20468
rect 20822 20412 20860 20468
rect 20916 20412 20926 20468
rect 22642 20412 22652 20468
rect 22708 20412 25788 20468
rect 25844 20412 25854 20468
rect 0 20384 800 20412
rect 13804 20356 13860 20412
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 10434 20300 10444 20356
rect 10500 20300 10668 20356
rect 10724 20300 10734 20356
rect 13794 20300 13804 20356
rect 13860 20300 15036 20356
rect 15092 20300 15102 20356
rect 15670 20300 15708 20356
rect 15764 20300 15774 20356
rect 16370 20300 16380 20356
rect 16436 20300 16828 20356
rect 16884 20300 16894 20356
rect 6178 20188 6188 20244
rect 6244 20188 7644 20244
rect 7700 20188 7710 20244
rect 9762 20188 9772 20244
rect 9828 20188 24444 20244
rect 24500 20188 24510 20244
rect 2818 20076 2828 20132
rect 2884 20076 5404 20132
rect 5460 20076 5470 20132
rect 9874 20076 9884 20132
rect 9940 20076 10780 20132
rect 10836 20076 10846 20132
rect 12450 20076 12460 20132
rect 12516 20076 21532 20132
rect 21588 20076 21598 20132
rect 23874 20076 23884 20132
rect 23940 20076 30380 20132
rect 30436 20076 30446 20132
rect 2370 19964 2380 20020
rect 2436 19964 3612 20020
rect 3668 19964 3678 20020
rect 4834 19964 4844 20020
rect 4900 19964 4956 20020
rect 5012 19964 5022 20020
rect 5618 19964 5628 20020
rect 5684 19964 15148 20020
rect 15204 19964 15214 20020
rect 16706 19964 16716 20020
rect 16772 19964 16828 20020
rect 16884 19964 17052 20020
rect 17108 19964 17118 20020
rect 17714 19964 17724 20020
rect 17780 19964 17790 20020
rect 19394 19964 19404 20020
rect 19460 19964 21420 20020
rect 21476 19964 21486 20020
rect 24994 19964 25004 20020
rect 25060 19964 27692 20020
rect 27748 19964 27758 20020
rect 17724 19908 17780 19964
rect 3042 19852 3052 19908
rect 3108 19852 4396 19908
rect 4452 19852 4462 19908
rect 6402 19852 6412 19908
rect 6468 19852 6478 19908
rect 8838 19852 8876 19908
rect 8932 19852 8942 19908
rect 9090 19852 9100 19908
rect 9156 19852 17780 19908
rect 18162 19852 18172 19908
rect 18228 19852 20188 19908
rect 20244 19852 20254 19908
rect 21046 19852 21084 19908
rect 21140 19852 21150 19908
rect 22082 19852 22092 19908
rect 22148 19852 26236 19908
rect 26292 19852 26302 19908
rect 29474 19852 29484 19908
rect 29540 19852 37660 19908
rect 37716 19852 37726 19908
rect 6412 19796 6468 19852
rect 1698 19740 1708 19796
rect 1764 19740 6468 19796
rect 15698 19740 15708 19796
rect 15764 19740 26684 19796
rect 26740 19740 26750 19796
rect 15586 19628 15596 19684
rect 15652 19628 17724 19684
rect 17780 19628 17790 19684
rect 20850 19628 20860 19684
rect 20916 19628 22428 19684
rect 22484 19628 22494 19684
rect 0 19572 800 19600
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 0 19516 2380 19572
rect 2436 19516 2446 19572
rect 14018 19516 14028 19572
rect 14084 19516 19964 19572
rect 20020 19516 20030 19572
rect 0 19488 800 19516
rect 11330 19404 11340 19460
rect 11396 19404 12348 19460
rect 12404 19404 12414 19460
rect 21644 19404 22428 19460
rect 22484 19404 22494 19460
rect 24070 19404 24108 19460
rect 24164 19404 24174 19460
rect 21644 19348 21700 19404
rect 6962 19292 6972 19348
rect 7028 19292 16716 19348
rect 16772 19292 16782 19348
rect 18060 19292 18508 19348
rect 18564 19292 18574 19348
rect 18834 19292 18844 19348
rect 18900 19292 21420 19348
rect 21476 19292 21700 19348
rect 21858 19292 21868 19348
rect 21924 19292 23212 19348
rect 23268 19292 23660 19348
rect 23716 19292 23726 19348
rect 18060 19236 18116 19292
rect 2706 19180 2716 19236
rect 2772 19180 5292 19236
rect 5348 19180 5358 19236
rect 9538 19180 9548 19236
rect 9604 19180 12908 19236
rect 12964 19180 12974 19236
rect 13654 19180 13692 19236
rect 13748 19180 13758 19236
rect 13990 19180 14028 19236
rect 14084 19180 14094 19236
rect 14802 19180 14812 19236
rect 14868 19180 18116 19236
rect 18386 19180 18396 19236
rect 18452 19180 24668 19236
rect 24724 19180 24734 19236
rect 1698 19068 1708 19124
rect 1764 19068 5740 19124
rect 5796 19068 5806 19124
rect 10770 19068 10780 19124
rect 10836 19068 11228 19124
rect 11284 19068 12796 19124
rect 12852 19068 12862 19124
rect 15362 19068 15372 19124
rect 15428 19068 15932 19124
rect 15988 19068 15998 19124
rect 18274 19068 18284 19124
rect 18340 19068 19180 19124
rect 19236 19068 19246 19124
rect 20524 19068 21532 19124
rect 21588 19068 21598 19124
rect 23986 19068 23996 19124
rect 24052 19068 24062 19124
rect 3826 18956 3836 19012
rect 3892 18956 4844 19012
rect 4900 18956 4910 19012
rect 9314 18956 9324 19012
rect 9380 18956 10332 19012
rect 10388 18956 10398 19012
rect 10994 18956 11004 19012
rect 11060 18956 11900 19012
rect 11956 18956 19628 19012
rect 19684 18956 20300 19012
rect 20356 18956 20366 19012
rect 10332 18900 10388 18956
rect 20524 18900 20580 19068
rect 23996 19012 24052 19068
rect 21970 18956 21980 19012
rect 22036 18956 24052 19012
rect 2706 18844 2716 18900
rect 2772 18844 2782 18900
rect 10332 18844 10780 18900
rect 10836 18844 10846 18900
rect 12348 18844 16380 18900
rect 16436 18844 16446 18900
rect 20178 18844 20188 18900
rect 20244 18844 20580 18900
rect 2716 18788 2772 18844
rect 12348 18788 12404 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 2258 18732 2268 18788
rect 2324 18732 2772 18788
rect 8754 18732 8764 18788
rect 8820 18732 12348 18788
rect 12404 18732 12414 18788
rect 0 18676 800 18704
rect 0 18620 1708 18676
rect 1764 18620 1774 18676
rect 2370 18620 2380 18676
rect 2436 18620 3052 18676
rect 3108 18620 3118 18676
rect 4162 18620 4172 18676
rect 4228 18620 8876 18676
rect 8932 18620 8942 18676
rect 9538 18620 9548 18676
rect 9604 18620 10556 18676
rect 10612 18620 10622 18676
rect 15260 18620 18284 18676
rect 18340 18620 18350 18676
rect 19058 18620 19068 18676
rect 19124 18620 19964 18676
rect 20020 18620 20030 18676
rect 0 18592 800 18620
rect 15260 18564 15316 18620
rect 2930 18508 2940 18564
rect 2996 18508 3948 18564
rect 4004 18508 4508 18564
rect 4564 18508 4574 18564
rect 5058 18508 5068 18564
rect 5124 18508 5180 18564
rect 5236 18508 5852 18564
rect 5908 18508 5918 18564
rect 15138 18508 15148 18564
rect 15204 18508 15316 18564
rect 17714 18508 17724 18564
rect 17780 18508 18172 18564
rect 18228 18508 18238 18564
rect 18498 18508 18508 18564
rect 18564 18508 21812 18564
rect 21756 18452 21812 18508
rect 8978 18396 8988 18452
rect 9044 18396 9548 18452
rect 9604 18396 9614 18452
rect 9762 18396 9772 18452
rect 9828 18396 10108 18452
rect 10164 18396 10174 18452
rect 14018 18396 14028 18452
rect 14084 18396 14588 18452
rect 14644 18396 14654 18452
rect 17938 18396 17948 18452
rect 18004 18396 18844 18452
rect 18900 18396 18910 18452
rect 19170 18396 19180 18452
rect 19236 18396 20860 18452
rect 20916 18396 20926 18452
rect 21756 18396 22876 18452
rect 22932 18396 22942 18452
rect 23492 18340 23548 18676
rect 23604 18620 23614 18676
rect 23996 18564 24052 18956
rect 23996 18508 24556 18564
rect 24612 18508 24622 18564
rect 23874 18396 23884 18452
rect 23940 18396 25004 18452
rect 25060 18396 25070 18452
rect 15026 18284 15036 18340
rect 15092 18284 15260 18340
rect 15316 18284 15326 18340
rect 15810 18284 15820 18340
rect 15876 18284 17276 18340
rect 17332 18284 17342 18340
rect 18386 18284 18396 18340
rect 18452 18284 21308 18340
rect 21364 18284 22652 18340
rect 22708 18284 22718 18340
rect 22876 18284 23548 18340
rect 7522 18172 7532 18228
rect 7588 18172 16044 18228
rect 16100 18172 16110 18228
rect 18834 18172 18844 18228
rect 18900 18172 19404 18228
rect 19460 18172 19470 18228
rect 20290 18172 20300 18228
rect 20356 18172 20636 18228
rect 20692 18172 20702 18228
rect 22876 18116 22932 18284
rect 23090 18172 23100 18228
rect 23156 18172 24108 18228
rect 24164 18172 24174 18228
rect 16706 18060 16716 18116
rect 16772 18060 19180 18116
rect 19236 18060 19246 18116
rect 21410 18060 21420 18116
rect 21476 18060 22932 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 2342 17948 2380 18004
rect 2436 17948 2446 18004
rect 11330 17948 11340 18004
rect 11396 17948 18396 18004
rect 18452 17948 18462 18004
rect 18946 17948 18956 18004
rect 19012 17948 19628 18004
rect 19684 17948 19694 18004
rect 20066 17948 20076 18004
rect 20132 17948 20188 18004
rect 20244 17948 20254 18004
rect 20636 17948 21644 18004
rect 21700 17948 21710 18004
rect 20636 17892 20692 17948
rect 5282 17836 5292 17892
rect 5348 17836 12012 17892
rect 12068 17836 12078 17892
rect 15698 17836 15708 17892
rect 15764 17836 16492 17892
rect 16548 17836 16558 17892
rect 18582 17836 18620 17892
rect 18676 17836 20692 17892
rect 21270 17836 21308 17892
rect 21364 17836 21374 17892
rect 22194 17836 22204 17892
rect 22260 17836 22540 17892
rect 22596 17836 24444 17892
rect 24500 17836 24510 17892
rect 0 17780 800 17808
rect 0 17724 1708 17780
rect 1764 17724 4620 17780
rect 4676 17724 4686 17780
rect 8082 17724 8092 17780
rect 8148 17724 13580 17780
rect 13636 17724 13646 17780
rect 14130 17724 14140 17780
rect 14196 17724 16156 17780
rect 16212 17724 16436 17780
rect 16706 17724 16716 17780
rect 16772 17724 21980 17780
rect 22036 17724 22046 17780
rect 0 17696 800 17724
rect 16380 17668 16436 17724
rect 1922 17612 1932 17668
rect 1988 17612 3276 17668
rect 3332 17612 3342 17668
rect 3826 17612 3836 17668
rect 3892 17612 8764 17668
rect 8820 17612 8830 17668
rect 11218 17612 11228 17668
rect 11284 17612 12012 17668
rect 12068 17612 12078 17668
rect 13010 17612 13020 17668
rect 13076 17612 13468 17668
rect 13524 17612 16156 17668
rect 16212 17612 16222 17668
rect 16380 17612 16604 17668
rect 16660 17612 17500 17668
rect 17556 17612 17566 17668
rect 18834 17612 18844 17668
rect 18900 17612 20412 17668
rect 20468 17612 20478 17668
rect 20962 17612 20972 17668
rect 21028 17612 22764 17668
rect 22820 17612 22830 17668
rect 24098 17612 24108 17668
rect 24164 17612 25676 17668
rect 25732 17612 25742 17668
rect 15138 17500 15148 17556
rect 15204 17500 15242 17556
rect 16034 17500 16044 17556
rect 16100 17500 16380 17556
rect 16436 17500 16446 17556
rect 16678 17500 16716 17556
rect 16772 17500 16782 17556
rect 18498 17500 18508 17556
rect 18564 17500 20076 17556
rect 20132 17500 22988 17556
rect 23044 17500 23054 17556
rect 10994 17388 11004 17444
rect 11060 17388 14140 17444
rect 14196 17388 14206 17444
rect 14578 17388 14588 17444
rect 14644 17388 15036 17444
rect 15092 17388 15372 17444
rect 15428 17388 18060 17444
rect 18116 17388 18956 17444
rect 19012 17388 19022 17444
rect 19730 17388 19740 17444
rect 19796 17388 20748 17444
rect 20804 17388 20814 17444
rect 1932 17276 5404 17332
rect 5460 17276 5470 17332
rect 8306 17276 8316 17332
rect 8372 17276 13356 17332
rect 13412 17276 13422 17332
rect 16594 17276 16604 17332
rect 16660 17276 17948 17332
rect 18004 17276 18844 17332
rect 18900 17276 18910 17332
rect 1932 17220 1988 17276
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 1922 17164 1932 17220
rect 1988 17164 1998 17220
rect 15670 17164 15708 17220
rect 15764 17164 15774 17220
rect 21634 17164 21644 17220
rect 21700 17164 22092 17220
rect 22148 17164 22158 17220
rect 3798 17052 3836 17108
rect 3892 17052 3902 17108
rect 4050 17052 4060 17108
rect 4116 17052 4284 17108
rect 4340 17052 4732 17108
rect 4788 17052 4798 17108
rect 7186 17052 7196 17108
rect 7252 17052 8652 17108
rect 8708 17052 8718 17108
rect 8978 17052 8988 17108
rect 9044 17052 9660 17108
rect 9716 17052 10668 17108
rect 10724 17052 11564 17108
rect 11620 17052 11630 17108
rect 13458 17052 13468 17108
rect 13524 17052 13692 17108
rect 13748 17052 13758 17108
rect 14018 17052 14028 17108
rect 14084 17052 15596 17108
rect 15652 17052 15662 17108
rect 15810 17052 15820 17108
rect 15876 17052 17612 17108
rect 17668 17052 18060 17108
rect 18116 17052 18126 17108
rect 18834 17052 18844 17108
rect 18900 17052 19180 17108
rect 19236 17052 19246 17108
rect 19618 17052 19628 17108
rect 19684 17052 21308 17108
rect 21364 17052 21374 17108
rect 21634 17052 21644 17108
rect 21700 17052 22876 17108
rect 22932 17052 22942 17108
rect 3938 16940 3948 16996
rect 4004 16940 7868 16996
rect 7924 16940 7934 16996
rect 10098 16940 10108 16996
rect 10164 16940 11228 16996
rect 11284 16940 11452 16996
rect 11508 16940 11518 16996
rect 12562 16940 12572 16996
rect 12628 16940 14364 16996
rect 14420 16940 16380 16996
rect 16436 16940 16446 16996
rect 19842 16940 19852 16996
rect 19908 16940 20188 16996
rect 20244 16940 22092 16996
rect 22148 16940 22158 16996
rect 0 16884 800 16912
rect 11452 16884 11508 16940
rect 0 16828 1708 16884
rect 1764 16828 1774 16884
rect 3826 16828 3836 16884
rect 3892 16828 6860 16884
rect 6916 16828 6926 16884
rect 7746 16828 7756 16884
rect 7812 16828 8988 16884
rect 9044 16828 10444 16884
rect 10500 16828 10510 16884
rect 10668 16828 10780 16884
rect 10836 16828 10846 16884
rect 11452 16828 12460 16884
rect 12516 16828 12526 16884
rect 14690 16828 14700 16884
rect 14756 16828 16604 16884
rect 16660 16828 16670 16884
rect 16828 16828 17836 16884
rect 17892 16828 17902 16884
rect 18162 16828 18172 16884
rect 18228 16828 21980 16884
rect 22036 16828 22046 16884
rect 0 16800 800 16828
rect 10668 16772 10724 16828
rect 16828 16772 16884 16828
rect 2258 16716 2268 16772
rect 2324 16716 2492 16772
rect 2548 16716 3164 16772
rect 3220 16716 3230 16772
rect 3602 16716 3612 16772
rect 3668 16716 4508 16772
rect 4564 16716 4574 16772
rect 4834 16716 4844 16772
rect 4900 16716 7420 16772
rect 7476 16716 7486 16772
rect 9958 16716 9996 16772
rect 10052 16716 10062 16772
rect 10658 16716 10668 16772
rect 10724 16716 10734 16772
rect 15026 16716 15036 16772
rect 15092 16716 15148 16772
rect 15204 16716 15214 16772
rect 16370 16716 16380 16772
rect 16436 16716 16884 16772
rect 19506 16716 19516 16772
rect 19572 16716 20188 16772
rect 20244 16716 20254 16772
rect 24770 16716 24780 16772
rect 24836 16716 30268 16772
rect 30324 16716 30334 16772
rect 13570 16604 13580 16660
rect 13636 16604 14140 16660
rect 14196 16604 14206 16660
rect 15586 16604 15596 16660
rect 15652 16604 16156 16660
rect 16212 16604 16222 16660
rect 13906 16492 13916 16548
rect 13972 16492 22092 16548
rect 22148 16492 22158 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 7858 16380 7868 16436
rect 7924 16380 9436 16436
rect 9492 16380 20524 16436
rect 20580 16380 21532 16436
rect 21588 16380 21598 16436
rect 3266 16268 3276 16324
rect 3332 16268 5068 16324
rect 5124 16268 5628 16324
rect 5684 16268 5694 16324
rect 12226 16268 12236 16324
rect 12292 16268 13244 16324
rect 13300 16268 13310 16324
rect 14578 16268 14588 16324
rect 14644 16268 17612 16324
rect 17668 16268 19068 16324
rect 19124 16268 19134 16324
rect 3714 16156 3724 16212
rect 3780 16156 4844 16212
rect 4900 16156 4910 16212
rect 11666 16156 11676 16212
rect 11732 16156 13692 16212
rect 13748 16156 13758 16212
rect 15362 16156 15372 16212
rect 15428 16156 15820 16212
rect 15876 16156 15886 16212
rect 18806 16156 18844 16212
rect 18900 16156 18910 16212
rect 1362 16044 1372 16100
rect 1428 16044 3612 16100
rect 3668 16044 3678 16100
rect 5170 16044 5180 16100
rect 5236 16044 5852 16100
rect 5908 16044 5918 16100
rect 10434 16044 10444 16100
rect 10500 16044 10780 16100
rect 10836 16044 10846 16100
rect 11778 16044 11788 16100
rect 11844 16044 12460 16100
rect 12516 16044 12526 16100
rect 13234 16044 13244 16100
rect 13300 16044 14924 16100
rect 14980 16044 16380 16100
rect 16436 16044 16446 16100
rect 17462 16044 17500 16100
rect 17556 16044 17566 16100
rect 19730 16044 19740 16100
rect 19796 16044 20748 16100
rect 20804 16044 21868 16100
rect 21924 16044 21934 16100
rect 22530 16044 22540 16100
rect 22596 16044 23100 16100
rect 23156 16044 23166 16100
rect 0 15988 800 16016
rect 0 15932 1484 15988
rect 1540 15932 1550 15988
rect 3154 15932 3164 15988
rect 3220 15932 4620 15988
rect 4676 15932 4686 15988
rect 8194 15932 8204 15988
rect 8260 15932 9212 15988
rect 9268 15932 9278 15988
rect 10210 15932 10220 15988
rect 10276 15932 12236 15988
rect 12292 15932 12302 15988
rect 14690 15932 14700 15988
rect 14756 15932 15932 15988
rect 15988 15932 15998 15988
rect 16146 15932 16156 15988
rect 16212 15932 16250 15988
rect 18498 15932 18508 15988
rect 18564 15932 19404 15988
rect 19460 15932 19470 15988
rect 0 15904 800 15932
rect 6066 15820 6076 15876
rect 6132 15820 8540 15876
rect 8596 15820 8606 15876
rect 10770 15820 10780 15876
rect 10836 15820 11900 15876
rect 11956 15820 11966 15876
rect 12562 15820 12572 15876
rect 12628 15820 15820 15876
rect 15876 15820 15886 15876
rect 16034 15820 16044 15876
rect 16100 15820 17164 15876
rect 17220 15820 17230 15876
rect 19618 15820 19628 15876
rect 19684 15820 20300 15876
rect 20356 15820 20366 15876
rect 21606 15820 21644 15876
rect 21700 15820 21710 15876
rect 22418 15820 22428 15876
rect 22484 15820 23100 15876
rect 23156 15820 23772 15876
rect 23828 15820 23838 15876
rect 1698 15708 1708 15764
rect 1764 15708 2492 15764
rect 2548 15708 2558 15764
rect 3602 15708 3612 15764
rect 3668 15708 4172 15764
rect 4228 15708 4238 15764
rect 7970 15708 7980 15764
rect 8036 15708 8652 15764
rect 8708 15708 10556 15764
rect 10612 15708 17052 15764
rect 17108 15708 17118 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 4022 15596 4060 15652
rect 4116 15596 4126 15652
rect 14018 15596 14028 15652
rect 14084 15596 16380 15652
rect 16436 15596 16446 15652
rect 10882 15484 10892 15540
rect 10948 15484 11676 15540
rect 11732 15484 11742 15540
rect 13010 15484 13020 15540
rect 13076 15484 13916 15540
rect 13972 15484 13982 15540
rect 10994 15372 11004 15428
rect 11060 15372 11228 15428
rect 11284 15372 12908 15428
rect 12964 15372 14812 15428
rect 14868 15372 14878 15428
rect 15092 15316 15148 15540
rect 15204 15484 17276 15540
rect 17332 15484 19516 15540
rect 19572 15484 22092 15540
rect 22148 15484 22158 15540
rect 16370 15372 16380 15428
rect 16436 15372 20524 15428
rect 20580 15372 20590 15428
rect 22754 15372 22764 15428
rect 22820 15372 23212 15428
rect 23268 15372 26012 15428
rect 26068 15372 26078 15428
rect 2370 15260 2380 15316
rect 2436 15260 2446 15316
rect 4610 15260 4620 15316
rect 4676 15260 7196 15316
rect 7252 15260 7262 15316
rect 12562 15260 12572 15316
rect 12628 15260 13468 15316
rect 13524 15260 13534 15316
rect 14466 15260 14476 15316
rect 14532 15260 15148 15316
rect 16146 15260 16156 15316
rect 16212 15260 18620 15316
rect 18676 15260 18686 15316
rect 22306 15260 22316 15316
rect 22372 15260 23324 15316
rect 23380 15260 23390 15316
rect 0 15092 800 15120
rect 2380 15092 2436 15260
rect 3276 15148 4956 15204
rect 5012 15148 5022 15204
rect 11666 15148 11676 15204
rect 11732 15148 14364 15204
rect 14420 15148 19740 15204
rect 19796 15148 19806 15204
rect 0 15036 2996 15092
rect 0 15008 800 15036
rect 2940 14980 2996 15036
rect 2930 14924 2940 14980
rect 2996 14924 3006 14980
rect 3276 14868 3332 15148
rect 12786 15036 12796 15092
rect 12852 15036 23884 15092
rect 23940 15036 23950 15092
rect 24658 15036 24668 15092
rect 24724 15036 24734 15092
rect 24668 14980 24724 15036
rect 14018 14924 14028 14980
rect 14084 14924 24724 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 3042 14812 3052 14868
rect 3108 14812 3332 14868
rect 21970 14812 21980 14868
rect 22036 14812 23100 14868
rect 23156 14812 23166 14868
rect 3826 14700 3836 14756
rect 3892 14700 5292 14756
rect 5348 14700 5358 14756
rect 14242 14700 14252 14756
rect 14308 14700 15372 14756
rect 15428 14700 16268 14756
rect 16324 14700 22036 14756
rect 2818 14588 2828 14644
rect 2884 14588 15148 14644
rect 15204 14588 15214 14644
rect 16146 14588 16156 14644
rect 16212 14588 18508 14644
rect 18564 14588 18574 14644
rect 14018 14476 14028 14532
rect 14084 14476 15372 14532
rect 15428 14476 15438 14532
rect 15596 14476 20076 14532
rect 20132 14476 20142 14532
rect 15596 14420 15652 14476
rect 21980 14420 22036 14700
rect 22194 14588 22204 14644
rect 22260 14588 22540 14644
rect 22596 14588 22606 14644
rect 1474 14364 1484 14420
rect 1540 14364 2492 14420
rect 2548 14364 2558 14420
rect 9986 14364 9996 14420
rect 10052 14364 15652 14420
rect 15708 14364 21588 14420
rect 21970 14364 21980 14420
rect 22036 14364 22652 14420
rect 22708 14364 22718 14420
rect 15708 14308 15764 14364
rect 21532 14308 21588 14364
rect 9874 14252 9884 14308
rect 9940 14252 15764 14308
rect 19842 14252 19852 14308
rect 19908 14252 20860 14308
rect 20916 14252 20926 14308
rect 21532 14252 21868 14308
rect 21924 14252 21934 14308
rect 0 14196 800 14224
rect 0 14140 1708 14196
rect 1764 14140 3388 14196
rect 3444 14140 3454 14196
rect 12226 14140 12236 14196
rect 12292 14140 19628 14196
rect 19684 14140 19694 14196
rect 0 14112 800 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 2034 13916 2044 13972
rect 2100 13916 3836 13972
rect 3892 13916 3902 13972
rect 10322 13916 10332 13972
rect 10388 13916 16268 13972
rect 16324 13916 16940 13972
rect 16996 13916 17006 13972
rect 18050 13916 18060 13972
rect 18116 13916 18956 13972
rect 19012 13916 19022 13972
rect 1138 13804 1148 13860
rect 1204 13804 12796 13860
rect 12852 13804 13244 13860
rect 13300 13804 13692 13860
rect 13748 13804 13758 13860
rect 3332 13692 6972 13748
rect 7028 13692 7038 13748
rect 1698 13580 1708 13636
rect 1764 13580 2940 13636
rect 2996 13580 3006 13636
rect 3332 13524 3388 13692
rect 2044 13468 3388 13524
rect 2044 13412 2100 13468
rect 2034 13356 2044 13412
rect 2100 13356 2110 13412
rect 0 13300 800 13328
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 0 13244 1708 13300
rect 1764 13244 1774 13300
rect 0 13216 800 13244
rect 3826 13132 3836 13188
rect 3892 13132 19292 13188
rect 19348 13132 19358 13188
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 0 12404 800 12432
rect 0 12348 1708 12404
rect 1764 12348 2492 12404
rect 2548 12348 2558 12404
rect 0 12320 800 12348
rect 1698 12012 1708 12068
rect 1764 12012 2492 12068
rect 2548 12012 2558 12068
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 8082 11564 8092 11620
rect 8148 11564 22876 11620
rect 22932 11564 22942 11620
rect 0 11508 800 11536
rect 0 11452 1708 11508
rect 1764 11452 1774 11508
rect 8866 11452 8876 11508
rect 8932 11452 21084 11508
rect 21140 11452 21150 11508
rect 0 11424 800 11452
rect 4050 11340 4060 11396
rect 4116 11340 22316 11396
rect 22372 11340 22382 11396
rect 1698 11116 1708 11172
rect 1764 11116 2492 11172
rect 2548 11116 2558 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 0 10612 800 10640
rect 0 10556 1708 10612
rect 1764 10556 1774 10612
rect 0 10528 800 10556
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 0 9716 800 9744
rect 0 9660 1932 9716
rect 1988 9660 2492 9716
rect 2548 9660 2558 9716
rect 0 9632 800 9660
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 2034 9212 2044 9268
rect 2100 9212 6300 9268
rect 6356 9212 6366 9268
rect 0 8820 800 8848
rect 0 8764 1708 8820
rect 1764 8764 2492 8820
rect 2548 8764 2558 8820
rect 0 8736 800 8764
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 2034 8092 2044 8148
rect 2100 8092 3724 8148
rect 3780 8092 3790 8148
rect 0 7924 800 7952
rect 0 7868 1708 7924
rect 1764 7868 2492 7924
rect 2548 7868 2558 7924
rect 0 7840 800 7868
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 2034 7644 2044 7700
rect 2100 7644 4844 7700
rect 4900 7644 4910 7700
rect 2034 7420 2044 7476
rect 2100 7420 4060 7476
rect 4116 7420 4126 7476
rect 0 7028 800 7056
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 0 6972 1708 7028
rect 1764 6972 2492 7028
rect 2548 6972 2558 7028
rect 0 6944 800 6972
rect 2146 6300 2156 6356
rect 2212 6300 3724 6356
rect 3780 6300 3790 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 0 6132 800 6160
rect 0 6076 1708 6132
rect 1764 6076 2492 6132
rect 2548 6076 2558 6132
rect 0 6048 800 6076
rect 1698 5740 1708 5796
rect 1764 5740 2492 5796
rect 2548 5740 2558 5796
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 0 5236 800 5264
rect 0 5180 1708 5236
rect 1764 5180 1774 5236
rect 0 5152 800 5180
rect 1698 4844 1708 4900
rect 1764 4844 2492 4900
rect 2548 4844 2558 4900
rect 1250 4732 1260 4788
rect 1316 4732 2044 4788
rect 2100 4732 2110 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 0 4340 800 4368
rect 0 4284 1708 4340
rect 1764 4284 1774 4340
rect 0 4256 800 4284
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 0 3444 800 3472
rect 0 3388 1708 3444
rect 1764 3388 2492 3444
rect 2548 3388 2558 3444
rect 0 3360 800 3388
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 21756 37884 21812 37940
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 15148 36428 15204 36484
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 15148 35980 15204 36036
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 19628 33964 19684 34020
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 14252 33516 14308 33572
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 18620 32396 18676 32452
rect 16268 32284 16324 32340
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 21980 31836 22036 31892
rect 15148 31276 15204 31332
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 12460 30156 12516 30212
rect 9324 29932 9380 29988
rect 22316 29932 22372 29988
rect 12572 29820 12628 29876
rect 18956 29820 19012 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 21420 29484 21476 29540
rect 13244 29260 13300 29316
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 21644 29148 21700 29204
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 8316 28812 8372 28868
rect 13804 28812 13860 28868
rect 13356 28588 13412 28644
rect 12572 28364 12628 28420
rect 14252 28364 14308 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 8876 28028 8932 28084
rect 12460 28028 12516 28084
rect 22316 27916 22372 27972
rect 15148 27804 15204 27860
rect 19068 27804 19124 27860
rect 21308 27692 21364 27748
rect 22204 27580 22260 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 22316 26908 22372 26964
rect 21980 26796 22036 26852
rect 16940 26684 16996 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 10780 26572 10836 26628
rect 22204 26572 22260 26628
rect 9324 26460 9380 26516
rect 19628 26460 19684 26516
rect 15372 26348 15428 26404
rect 19292 26348 19348 26404
rect 18732 26236 18788 26292
rect 18956 26236 19012 26292
rect 19516 26236 19572 26292
rect 19628 26012 19684 26068
rect 21308 25900 21364 25956
rect 21644 25900 21700 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 11004 25676 11060 25732
rect 18844 25564 18900 25620
rect 19180 25340 19236 25396
rect 20188 25340 20244 25396
rect 16940 25116 16996 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4060 24892 4116 24948
rect 16268 24892 16324 24948
rect 17724 24780 17780 24836
rect 18956 24780 19012 24836
rect 19180 24780 19236 24836
rect 13244 24668 13300 24724
rect 18732 24556 18788 24612
rect 19180 24556 19236 24612
rect 4844 24444 4900 24500
rect 10220 24332 10276 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 18508 24444 18564 24500
rect 20188 24332 20244 24388
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 11228 23884 11284 23940
rect 21308 23884 21364 23940
rect 4060 23660 4116 23716
rect 21420 23660 21476 23716
rect 4844 23548 4900 23604
rect 18508 23548 18564 23604
rect 18844 23548 18900 23604
rect 19180 23548 19236 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 11004 23436 11060 23492
rect 16940 23436 16996 23492
rect 17500 23436 17556 23492
rect 3612 23324 3668 23380
rect 16604 23324 16660 23380
rect 19628 23324 19684 23380
rect 10220 23212 10276 23268
rect 17164 22876 17220 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 3388 22540 3444 22596
rect 15708 22540 15764 22596
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19628 22428 19684 22484
rect 24220 22428 24276 22484
rect 24108 22316 24164 22372
rect 3724 22204 3780 22260
rect 20188 22092 20244 22148
rect 10668 21980 10724 22036
rect 2380 21868 2436 21924
rect 4060 21756 4116 21812
rect 8316 21756 8372 21812
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 20860 21868 20916 21924
rect 19516 21756 19572 21812
rect 21756 21756 21812 21812
rect 4844 21644 4900 21700
rect 15708 21644 15764 21700
rect 24220 21644 24276 21700
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 5180 21084 5236 21140
rect 11228 20972 11284 21028
rect 21308 21196 21364 21252
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 15708 20748 15764 20804
rect 17164 20748 17220 20804
rect 3388 20524 3444 20580
rect 16604 20524 16660 20580
rect 19628 20412 19684 20468
rect 20860 20412 20916 20468
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 10668 20300 10724 20356
rect 15036 20300 15092 20356
rect 15708 20300 15764 20356
rect 4844 19964 4900 20020
rect 16716 19964 16772 20020
rect 8876 19852 8932 19908
rect 21084 19852 21140 19908
rect 17724 19628 17780 19684
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 24108 19404 24164 19460
rect 13692 19180 13748 19236
rect 14028 19180 14084 19236
rect 20188 18844 20244 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 19068 18620 19124 18676
rect 5180 18508 5236 18564
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 2380 17948 2436 18004
rect 20188 17948 20244 18004
rect 18620 17836 18676 17892
rect 21308 17836 21364 17892
rect 16156 17724 16212 17780
rect 15148 17500 15204 17556
rect 16716 17500 16772 17556
rect 16604 17276 16660 17332
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 15708 17164 15764 17220
rect 3836 17052 3892 17108
rect 13692 17052 13748 17108
rect 18844 17052 18900 17108
rect 21644 17052 21700 17108
rect 20188 16940 20244 16996
rect 10780 16828 10836 16884
rect 3612 16716 3668 16772
rect 9996 16716 10052 16772
rect 15036 16716 15092 16772
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 18844 16156 18900 16212
rect 17500 16044 17556 16100
rect 16156 15932 16212 15988
rect 21644 15820 21700 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4060 15596 4116 15652
rect 14028 15596 14084 15652
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 15148 14588 15204 14644
rect 15372 14476 15428 14532
rect 9996 14364 10052 14420
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 3836 13132 3892 13188
rect 19292 13132 19348 13188
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 21084 11452 21140 11508
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 3724 8092 3780 8148
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 19808 37660 20128 38476
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 15148 36484 15204 36494
rect 15148 36036 15204 36428
rect 15148 35970 15204 35980
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 19628 34020 19684 34030
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 14252 33572 14308 33582
rect 12460 30212 12516 30222
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 9324 29988 9380 29998
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4060 24948 4116 24958
rect 4060 23716 4116 24892
rect 4060 23650 4116 23660
rect 4448 24332 4768 25844
rect 8316 28868 8372 28878
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 3612 23380 3668 23390
rect 3388 22596 3444 22606
rect 2380 21924 2436 21934
rect 2380 18004 2436 21868
rect 3388 20580 3444 22540
rect 3388 20514 3444 20524
rect 2380 17938 2436 17948
rect 3612 16772 3668 23324
rect 4448 22764 4768 24276
rect 4844 24500 4900 24510
rect 4844 23604 4900 24444
rect 4844 23538 4900 23548
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 3612 16706 3668 16716
rect 3724 22260 3780 22270
rect 3724 8148 3780 22204
rect 4060 21812 4116 21822
rect 3836 17108 3892 17118
rect 3836 13188 3892 17052
rect 4060 15652 4116 21756
rect 4060 15586 4116 15596
rect 4448 21196 4768 22708
rect 8316 21812 8372 28812
rect 8316 21746 8372 21756
rect 8876 28084 8932 28094
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4844 21700 4900 21710
rect 4844 20020 4900 21644
rect 4844 19954 4900 19964
rect 5180 21140 5236 21150
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 5180 18564 5236 21084
rect 8876 19908 8932 28028
rect 9324 26516 9380 29932
rect 12460 28084 12516 30156
rect 12572 29876 12628 29886
rect 12572 28420 12628 29820
rect 12572 28354 12628 28364
rect 13244 29316 13300 29326
rect 12460 28018 12516 28028
rect 9324 26450 9380 26460
rect 10780 26628 10836 26638
rect 10220 24388 10276 24398
rect 10220 23268 10276 24332
rect 10220 23202 10276 23212
rect 10668 22036 10724 22046
rect 10668 20356 10724 21980
rect 10668 20290 10724 20300
rect 8876 19842 8932 19852
rect 5180 18498 5236 18508
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 10780 16884 10836 26572
rect 11004 25732 11060 25742
rect 11004 23492 11060 25676
rect 13244 24724 13300 29260
rect 13804 28868 13860 28878
rect 13804 28738 13860 28812
rect 13356 28682 13860 28738
rect 13356 28644 13412 28682
rect 13356 28578 13412 28588
rect 14252 28420 14308 33516
rect 18620 32452 18676 32462
rect 16268 32340 16324 32350
rect 14252 28354 14308 28364
rect 15148 31332 15204 31342
rect 15148 27860 15204 31276
rect 15148 27794 15204 27804
rect 13244 24658 13300 24668
rect 15372 26404 15428 26414
rect 11004 23426 11060 23436
rect 11228 23940 11284 23950
rect 11228 21028 11284 23884
rect 11228 20962 11284 20972
rect 15036 20356 15092 20366
rect 13692 19236 13748 19246
rect 13692 17108 13748 19180
rect 13692 17042 13748 17052
rect 14028 19236 14084 19246
rect 10780 16818 10836 16828
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 3836 13122 3892 13132
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 9996 16772 10052 16782
rect 9996 14420 10052 16716
rect 14028 15652 14084 19180
rect 15036 16772 15092 20300
rect 15036 16706 15092 16716
rect 15148 17556 15204 17566
rect 14028 15586 14084 15596
rect 15148 14644 15204 17500
rect 15148 14578 15204 14588
rect 15372 14532 15428 26348
rect 16268 24948 16324 32284
rect 16268 24882 16324 24892
rect 16940 26740 16996 26750
rect 16940 25172 16996 26684
rect 16940 23492 16996 25116
rect 17724 24836 17780 24846
rect 16940 23426 16996 23436
rect 17500 23492 17556 23502
rect 16604 23380 16660 23390
rect 15708 22596 15764 22606
rect 15708 21700 15764 22540
rect 15708 20804 15764 21644
rect 15708 20738 15764 20748
rect 16604 20580 16660 23324
rect 17164 22932 17220 22942
rect 17164 20804 17220 22876
rect 17164 20738 17220 20748
rect 15708 20356 15764 20366
rect 15708 17220 15764 20300
rect 15708 17154 15764 17164
rect 16156 17780 16212 17790
rect 16156 15988 16212 17724
rect 16604 17332 16660 20524
rect 16716 20020 16772 20030
rect 16716 17556 16772 19964
rect 16716 17490 16772 17500
rect 16604 17266 16660 17276
rect 17500 16100 17556 23436
rect 17724 19684 17780 24780
rect 18508 24500 18564 24510
rect 18508 23604 18564 24444
rect 18508 23538 18564 23548
rect 17724 19618 17780 19628
rect 18620 17892 18676 32396
rect 18956 29876 19012 29886
rect 18732 26292 18788 26302
rect 18732 24612 18788 26236
rect 18956 26292 19012 29820
rect 18732 24546 18788 24556
rect 18844 25620 18900 25630
rect 18844 23604 18900 25564
rect 18956 24836 19012 26236
rect 18956 24770 19012 24780
rect 19068 27860 19124 27870
rect 18844 23538 18900 23548
rect 19068 18676 19124 27804
rect 19628 26516 19684 33964
rect 19628 26450 19684 26460
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 21756 37940 21812 37950
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 21420 29540 21476 29550
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19292 26404 19348 26414
rect 19180 25396 19236 25406
rect 19180 24836 19236 25340
rect 19180 24770 19236 24780
rect 19180 24612 19236 24622
rect 19180 23604 19236 24556
rect 19180 23538 19236 23548
rect 19068 18610 19124 18620
rect 18620 17826 18676 17836
rect 18844 17108 18900 17118
rect 18844 16212 18900 17052
rect 18844 16146 18900 16156
rect 17500 16034 17556 16044
rect 16156 15922 16212 15932
rect 15372 14466 15428 14476
rect 9996 14354 10052 14364
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 3724 8082 3780 8092
rect 4448 11788 4768 13300
rect 19292 13188 19348 26348
rect 19516 26292 19572 26302
rect 19516 21812 19572 26236
rect 19516 21746 19572 21756
rect 19628 26068 19684 26078
rect 19628 23380 19684 26012
rect 19628 22484 19684 23324
rect 19628 20468 19684 22428
rect 19628 20402 19684 20412
rect 19808 25116 20128 26628
rect 21308 27748 21364 27758
rect 21308 25956 21364 27692
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 20188 25396 20244 25406
rect 20188 24388 20244 25340
rect 20188 24322 20244 24332
rect 21308 23940 21364 25900
rect 21308 23874 21364 23884
rect 21420 23716 21476 29484
rect 21644 29204 21700 29214
rect 21644 25956 21700 29148
rect 21644 25890 21700 25900
rect 21420 23650 21476 23660
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19292 13122 19348 13132
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 20188 22148 20244 22158
rect 20188 18900 20244 22092
rect 20860 21924 20916 21934
rect 20860 20468 20916 21868
rect 21756 21812 21812 37884
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 21980 31892 22036 31902
rect 21980 26852 22036 31836
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 22316 29988 22372 29998
rect 22316 27972 22372 29932
rect 21980 26786 22036 26796
rect 22204 27636 22260 27646
rect 22204 26628 22260 27580
rect 22316 26964 22372 27916
rect 22316 26898 22372 26908
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 22204 26562 22260 26572
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 24220 22484 24276 22494
rect 21756 21746 21812 21756
rect 24108 22372 24164 22382
rect 20860 20402 20916 20412
rect 21308 21252 21364 21262
rect 20188 18834 20244 18844
rect 21084 19908 21140 19918
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 20188 18004 20244 18014
rect 20188 16996 20244 17948
rect 20188 16930 20244 16940
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 21084 11508 21140 19852
rect 21308 17892 21364 21196
rect 24108 19460 24164 22316
rect 24220 21700 24276 22428
rect 24220 21634 24276 21644
rect 24108 19394 24164 19404
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 21308 17826 21364 17836
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 21644 17108 21700 17118
rect 21644 15876 21700 17052
rect 21644 15810 21700 15820
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 21084 11442 21140 11452
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _386_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _387_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3696 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _388_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5712 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _389_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3136 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _390_
timestamp 1698431365
transform 1 0 2016 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _391_
timestamp 1698431365
transform 1 0 6384 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _392_
timestamp 1698431365
transform 1 0 7952 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _393_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _394_
timestamp 1698431365
transform 1 0 11536 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _395_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _396_
timestamp 1698431365
transform 1 0 1792 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _397_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3696 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _398_
timestamp 1698431365
transform -1 0 3360 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _399_
timestamp 1698431365
transform 1 0 2800 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _400_
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _401_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4032 0 -1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _402_
timestamp 1698431365
transform 1 0 16352 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _403_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19712 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _404_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22848 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _405_
timestamp 1698431365
transform 1 0 2016 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _406_
timestamp 1698431365
transform -1 0 3360 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _407_
timestamp 1698431365
transform -1 0 3136 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _408_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _409_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5264 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _410_
timestamp 1698431365
transform 1 0 16800 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _411_
timestamp 1698431365
transform -1 0 3808 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _412_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12432 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _413_
timestamp 1698431365
transform 1 0 2800 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  _414_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12768 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _415_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6720 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _416_
timestamp 1698431365
transform 1 0 2352 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _417_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4144 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _418_
timestamp 1698431365
transform 1 0 8960 0 1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _419_
timestamp 1698431365
transform 1 0 14672 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _420_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17920 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _421_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4592 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _422_
timestamp 1698431365
transform -1 0 5264 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _423_
timestamp 1698431365
transform 1 0 13776 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _424_
timestamp 1698431365
transform 1 0 4592 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _425_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4592 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _426_
timestamp 1698431365
transform 1 0 17024 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _427_
timestamp 1698431365
transform -1 0 21392 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _428_
timestamp 1698431365
transform 1 0 18704 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _429_
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _430_
timestamp 1698431365
transform 1 0 2016 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _431_
timestamp 1698431365
transform -1 0 4592 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _432_
timestamp 1698431365
transform 1 0 3808 0 -1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _433_
timestamp 1698431365
transform 1 0 13776 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _434_
timestamp 1698431365
transform 1 0 20272 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _435_
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _436_
timestamp 1698431365
transform 1 0 1904 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _437_
timestamp 1698431365
transform 1 0 7728 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _438_
timestamp 1698431365
transform 1 0 10976 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _439_
timestamp 1698431365
transform 1 0 18368 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _440_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _441_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _442_
timestamp 1698431365
transform -1 0 15344 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _443_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18928 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _444_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20720 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _445_
timestamp 1698431365
transform -1 0 4480 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _446_
timestamp 1698431365
transform -1 0 2800 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _447_
timestamp 1698431365
transform 1 0 2800 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _448_
timestamp 1698431365
transform -1 0 4480 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _449_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _450_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11088 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _451_
timestamp 1698431365
transform 1 0 13888 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _452_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6608 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _453_
timestamp 1698431365
transform 1 0 10304 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _454_
timestamp 1698431365
transform 1 0 14560 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _455_
timestamp 1698431365
transform -1 0 16464 0 -1 36064
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _456_
timestamp 1698431365
transform -1 0 14448 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _457_
timestamp 1698431365
transform 1 0 13440 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _458_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _459_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11424 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _460_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23072 0 -1 23520
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _461_
timestamp 1698431365
transform 1 0 7056 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _462_
timestamp 1698431365
transform 1 0 8288 0 1 36064
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _463_
timestamp 1698431365
transform 1 0 11872 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _464_
timestamp 1698431365
transform -1 0 12880 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _465_
timestamp 1698431365
transform 1 0 3360 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _466_
timestamp 1698431365
transform 1 0 4480 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _467_
timestamp 1698431365
transform 1 0 2688 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _468_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8400 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _469_
timestamp 1698431365
transform -1 0 17248 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _470_
timestamp 1698431365
transform -1 0 6944 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _471_
timestamp 1698431365
transform 1 0 11200 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _472_
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _473_
timestamp 1698431365
transform -1 0 15792 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _474_
timestamp 1698431365
transform -1 0 15120 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _475_
timestamp 1698431365
transform 1 0 13216 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _476_
timestamp 1698431365
transform 1 0 11536 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _477_
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _478_
timestamp 1698431365
transform 1 0 12320 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _479_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _480_
timestamp 1698431365
transform -1 0 9184 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _481_
timestamp 1698431365
transform -1 0 3136 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _482_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _483_
timestamp 1698431365
transform -1 0 6384 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _484_
timestamp 1698431365
transform -1 0 5264 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _485_
timestamp 1698431365
transform -1 0 6160 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _486_
timestamp 1698431365
transform 1 0 3024 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _487_
timestamp 1698431365
transform 1 0 9744 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _488_
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _489_
timestamp 1698431365
transform 1 0 8736 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _490_
timestamp 1698431365
transform 1 0 9296 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _491_
timestamp 1698431365
transform 1 0 9408 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _492_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8512 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _493_
timestamp 1698431365
transform 1 0 3696 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _494_
timestamp 1698431365
transform 1 0 1680 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _495_
timestamp 1698431365
transform -1 0 6832 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _496_
timestamp 1698431365
transform 1 0 3584 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _497_
timestamp 1698431365
transform -1 0 5264 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _498_
timestamp 1698431365
transform -1 0 6160 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _499_
timestamp 1698431365
transform 1 0 1904 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _500_
timestamp 1698431365
transform 1 0 2576 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _501_
timestamp 1698431365
transform -1 0 10528 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _502_
timestamp 1698431365
transform -1 0 8624 0 -1 32928
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _503_
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _504_
timestamp 1698431365
transform -1 0 19264 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _505_
timestamp 1698431365
transform 1 0 3136 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _506_
timestamp 1698431365
transform 1 0 3136 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _507_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3808 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _508_
timestamp 1698431365
transform -1 0 10528 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _509_
timestamp 1698431365
transform -1 0 6160 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _510_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5712 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _511_
timestamp 1698431365
transform -1 0 8400 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _512_
timestamp 1698431365
transform -1 0 16016 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _513_
timestamp 1698431365
transform 1 0 8400 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _514_
timestamp 1698431365
transform 1 0 10528 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _515_
timestamp 1698431365
transform 1 0 10304 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _516_
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _517_
timestamp 1698431365
transform -1 0 13776 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _518_
timestamp 1698431365
transform -1 0 18256 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _519_
timestamp 1698431365
transform 1 0 18032 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _520_
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _521_
timestamp 1698431365
transform 1 0 11200 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _522_
timestamp 1698431365
transform -1 0 11088 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _523_
timestamp 1698431365
transform 1 0 19936 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _524_
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _525_
timestamp 1698431365
transform 1 0 7840 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _526_
timestamp 1698431365
transform 1 0 16128 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _527_
timestamp 1698431365
transform 1 0 6944 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _528_
timestamp 1698431365
transform 1 0 8512 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _529_
timestamp 1698431365
transform -1 0 18816 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _530_
timestamp 1698431365
transform 1 0 14896 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _531_
timestamp 1698431365
transform -1 0 16240 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _532_
timestamp 1698431365
transform 1 0 15120 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _533_
timestamp 1698431365
transform -1 0 19600 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _534_
timestamp 1698431365
transform -1 0 7168 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _535_
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _536_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _537_
timestamp 1698431365
transform -1 0 20048 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _538_
timestamp 1698431365
transform 1 0 19936 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _539_
timestamp 1698431365
transform -1 0 7840 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _540_
timestamp 1698431365
transform 1 0 19040 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _541_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19600 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _542_
timestamp 1698431365
transform 1 0 16240 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _543_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10640 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _544_
timestamp 1698431365
transform 1 0 4368 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _545_
timestamp 1698431365
transform -1 0 8064 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _546_
timestamp 1698431365
transform -1 0 6944 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _547_
timestamp 1698431365
transform -1 0 7952 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _548_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11200 0 -1 31360
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _549_
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _550_
timestamp 1698431365
transform 1 0 25536 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _551_
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _552_
timestamp 1698431365
transform 1 0 12992 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _553_
timestamp 1698431365
transform 1 0 13888 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _554_
timestamp 1698431365
transform -1 0 14560 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _555_
timestamp 1698431365
transform 1 0 14560 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _556_
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _557_
timestamp 1698431365
transform 1 0 15232 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _558_
timestamp 1698431365
transform 1 0 16352 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _559_
timestamp 1698431365
transform 1 0 14896 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _560_
timestamp 1698431365
transform 1 0 11984 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _561_
timestamp 1698431365
transform -1 0 16912 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _562_
timestamp 1698431365
transform -1 0 18368 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _563_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17920 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _564_
timestamp 1698431365
transform 1 0 18256 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _565_
timestamp 1698431365
transform -1 0 20160 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _566_
timestamp 1698431365
transform 1 0 4256 0 -1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _567_
timestamp 1698431365
transform -1 0 18256 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _568_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _569_
timestamp 1698431365
transform -1 0 8736 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _570_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9296 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _571_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _572_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _573_
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _574_
timestamp 1698431365
transform -1 0 15456 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _575_
timestamp 1698431365
transform -1 0 14896 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _576_
timestamp 1698431365
transform 1 0 10080 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _577_
timestamp 1698431365
transform -1 0 11760 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _578_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17696 0 1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _579_
timestamp 1698431365
transform 1 0 13440 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _580_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13776 0 1 29792
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _581_
timestamp 1698431365
transform 1 0 24192 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _582_
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _583_
timestamp 1698431365
transform 1 0 9744 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _584_
timestamp 1698431365
transform 1 0 10416 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _585_
timestamp 1698431365
transform -1 0 12096 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _586_
timestamp 1698431365
transform 1 0 12096 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _587_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _588_
timestamp 1698431365
transform 1 0 23856 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _589_
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _590_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _591_
timestamp 1698431365
transform -1 0 16800 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _592_
timestamp 1698431365
transform 1 0 12096 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _593_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14672 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _594_
timestamp 1698431365
transform -1 0 24192 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _595_
timestamp 1698431365
transform -1 0 25872 0 1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _596_
timestamp 1698431365
transform 1 0 21504 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _597_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _598_
timestamp 1698431365
transform 1 0 13552 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _599_
timestamp 1698431365
transform -1 0 22288 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _600_
timestamp 1698431365
transform -1 0 23072 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _601_
timestamp 1698431365
transform 1 0 8176 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _602_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _603_
timestamp 1698431365
transform 1 0 22400 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _604_
timestamp 1698431365
transform 1 0 22400 0 1 17248
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _605_
timestamp 1698431365
transform 1 0 17024 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _606_
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _607_
timestamp 1698431365
transform 1 0 20048 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _608_
timestamp 1698431365
transform -1 0 16352 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _609_
timestamp 1698431365
transform 1 0 19824 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _610_
timestamp 1698431365
transform 1 0 18256 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _611_
timestamp 1698431365
transform -1 0 20160 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _612_
timestamp 1698431365
transform 1 0 19488 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _613_
timestamp 1698431365
transform 1 0 21280 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _614_
timestamp 1698431365
transform -1 0 24080 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _615_
timestamp 1698431365
transform 1 0 23072 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _616_
timestamp 1698431365
transform 1 0 11760 0 -1 26656
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _617_
timestamp 1698431365
transform -1 0 24304 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _618_
timestamp 1698431365
transform -1 0 23296 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _619_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _620_
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _621_
timestamp 1698431365
transform 1 0 8288 0 1 26656
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _622_
timestamp 1698431365
transform 1 0 14896 0 1 23520
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _623_
timestamp 1698431365
transform 1 0 3360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _624_
timestamp 1698431365
transform 1 0 4368 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _625_
timestamp 1698431365
transform 1 0 7280 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _626_
timestamp 1698431365
transform 1 0 16016 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _627_
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _628_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15008 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _629_
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _630_
timestamp 1698431365
transform 1 0 14560 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _631_
timestamp 1698431365
transform 1 0 16016 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _632_
timestamp 1698431365
transform -1 0 7056 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _633_
timestamp 1698431365
transform 1 0 17696 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _634_
timestamp 1698431365
transform 1 0 12880 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _635_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _636_
timestamp 1698431365
transform -1 0 5152 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _637_
timestamp 1698431365
transform -1 0 5264 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _638_
timestamp 1698431365
transform 1 0 2576 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _639_
timestamp 1698431365
transform 1 0 15456 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _640_
timestamp 1698431365
transform 1 0 14896 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _641_
timestamp 1698431365
transform 1 0 14784 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _642_
timestamp 1698431365
transform 1 0 15680 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _643_
timestamp 1698431365
transform -1 0 23072 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _644_
timestamp 1698431365
transform -1 0 21504 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _645_
timestamp 1698431365
transform 1 0 19600 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _646_
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _647_
timestamp 1698431365
transform 1 0 4592 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _648_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _649_
timestamp 1698431365
transform -1 0 16016 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _650_
timestamp 1698431365
transform 1 0 11760 0 -1 23520
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _651_
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _652_
timestamp 1698431365
transform 1 0 8624 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _653_
timestamp 1698431365
transform 1 0 15680 0 1 21952
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _654_
timestamp 1698431365
transform 1 0 23520 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _655_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _656_
timestamp 1698431365
transform -1 0 23632 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _657_
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _658_
timestamp 1698431365
transform 1 0 23184 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _659_
timestamp 1698431365
transform 1 0 21504 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _660_
timestamp 1698431365
transform 1 0 22736 0 1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _661_
timestamp 1698431365
transform 1 0 24528 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _662_
timestamp 1698431365
transform -1 0 20272 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _663_
timestamp 1698431365
transform 1 0 15680 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _664_
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _665_
timestamp 1698431365
transform 1 0 14896 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _666_
timestamp 1698431365
transform 1 0 11424 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _667_
timestamp 1698431365
transform 1 0 18256 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _668_
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _669_
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _670_
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _671_
timestamp 1698431365
transform -1 0 9184 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _672_
timestamp 1698431365
transform -1 0 17920 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _673_
timestamp 1698431365
transform 1 0 17360 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _674_
timestamp 1698431365
transform 1 0 15568 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _675_
timestamp 1698431365
transform 1 0 15680 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _676_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _677_
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _678_
timestamp 1698431365
transform 1 0 2576 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _679_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8064 0 1 21952
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _680_
timestamp 1698431365
transform -1 0 13888 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _681_
timestamp 1698431365
transform -1 0 12768 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _682_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _683_
timestamp 1698431365
transform -1 0 5264 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _684_
timestamp 1698431365
transform -1 0 10304 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _685_
timestamp 1698431365
transform 1 0 7728 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _686_
timestamp 1698431365
transform 1 0 8288 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _687_
timestamp 1698431365
transform 1 0 3584 0 -1 15680
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _688_
timestamp 1698431365
transform -1 0 9296 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _689_
timestamp 1698431365
transform -1 0 24528 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _690_
timestamp 1698431365
transform 1 0 23184 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _691_
timestamp 1698431365
transform 1 0 27104 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _692_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20048 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _693_
timestamp 1698431365
transform -1 0 28000 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _694_
timestamp 1698431365
transform 1 0 22288 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _695_
timestamp 1698431365
transform 1 0 19040 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _696_
timestamp 1698431365
transform 1 0 11088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _697_
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _698_
timestamp 1698431365
transform 1 0 20272 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _699_
timestamp 1698431365
transform 1 0 18816 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _700_
timestamp 1698431365
transform 1 0 20048 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _701_
timestamp 1698431365
transform 1 0 11312 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _702_
timestamp 1698431365
transform 1 0 3584 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _703_
timestamp 1698431365
transform 1 0 11312 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _704_
timestamp 1698431365
transform 1 0 2352 0 1 18816
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _705_
timestamp 1698431365
transform 1 0 21168 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _706_
timestamp 1698431365
transform -1 0 10864 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _707_
timestamp 1698431365
transform -1 0 4480 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _708_
timestamp 1698431365
transform 1 0 7728 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _709_
timestamp 1698431365
transform -1 0 22176 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _710_
timestamp 1698431365
transform 1 0 16016 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _711_
timestamp 1698431365
transform 1 0 21840 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _712_
timestamp 1698431365
transform 1 0 19152 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _713_
timestamp 1698431365
transform -1 0 20720 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _714_
timestamp 1698431365
transform 1 0 18480 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _715_
timestamp 1698431365
transform 1 0 17920 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _716_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23408 0 1 26656
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _717_
timestamp 1698431365
transform 1 0 25424 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _718_
timestamp 1698431365
transform -1 0 26880 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _719_
timestamp 1698431365
transform 1 0 25424 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _720_
timestamp 1698431365
transform 1 0 25760 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _721_
timestamp 1698431365
transform 1 0 28000 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _722_
timestamp 1698431365
transform 1 0 18928 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _723_
timestamp 1698431365
transform 1 0 25200 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _724_
timestamp 1698431365
transform -1 0 4368 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _725_
timestamp 1698431365
transform -1 0 4368 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _726_
timestamp 1698431365
transform 1 0 10528 0 -1 18816
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _727_
timestamp 1698431365
transform -1 0 10304 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _728_
timestamp 1698431365
transform 1 0 20832 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _729_
timestamp 1698431365
transform 1 0 22848 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _730_
timestamp 1698431365
transform 1 0 19600 0 -1 15680
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _731_
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _732_
timestamp 1698431365
transform 1 0 24640 0 1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _733_
timestamp 1698431365
transform 1 0 26768 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _734_
timestamp 1698431365
transform -1 0 26320 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _735_
timestamp 1698431365
transform -1 0 4368 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _736_
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _737_
timestamp 1698431365
transform 1 0 19040 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _738_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _739_
timestamp 1698431365
transform -1 0 15120 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _740_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 25088
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _741_
timestamp 1698431365
transform -1 0 22736 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _742_
timestamp 1698431365
transform 1 0 21280 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _743_
timestamp 1698431365
transform -1 0 24416 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _744_
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _745_
timestamp 1698431365
transform -1 0 19936 0 1 18816
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _746_
timestamp 1698431365
transform 1 0 3584 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _747_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _748_
timestamp 1698431365
transform -1 0 27104 0 1 25088
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _749_
timestamp 1698431365
transform -1 0 28560 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _750_
timestamp 1698431365
transform -1 0 8848 0 -1 21952
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _751_
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _752_
timestamp 1698431365
transform 1 0 11760 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _753_
timestamp 1698431365
transform 1 0 10640 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _754_
timestamp 1698431365
transform 1 0 21168 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _755_
timestamp 1698431365
transform 1 0 20944 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _756_
timestamp 1698431365
transform 1 0 8512 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _757_
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _758_
timestamp 1698431365
transform 1 0 7168 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _759_
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _760_
timestamp 1698431365
transform -1 0 10304 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _761_
timestamp 1698431365
transform -1 0 9184 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _762_
timestamp 1698431365
transform -1 0 12768 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _763_
timestamp 1698431365
transform 1 0 11424 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _764_
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _765_
timestamp 1698431365
transform 1 0 10528 0 -1 25088
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _766_
timestamp 1698431365
transform -1 0 28224 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _767_
timestamp 1698431365
transform 1 0 23632 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _768_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6944 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _769_
timestamp 1698431365
transform 1 0 23408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _770_
timestamp 1698431365
transform 1 0 23856 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _771_
timestamp 1698431365
transform 1 0 23856 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _772_
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _773_
timestamp 1698431365
transform 1 0 2576 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _774_
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _775_
timestamp 1698431365
transform 1 0 5152 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _776_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _777_
timestamp 1698431365
transform 1 0 12992 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _778_
timestamp 1698431365
transform 1 0 14784 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _779_
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__A1 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__A2
timestamp 1698431365
transform 1 0 20496 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__I
timestamp 1698431365
transform 1 0 12880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__A1
timestamp 1698431365
transform -1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__A1
timestamp 1698431365
transform 1 0 18032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__I
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__I
timestamp 1698431365
transform -1 0 19488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__I
timestamp 1698431365
transform -1 0 13328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__I
timestamp 1698431365
transform 1 0 15680 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__I
timestamp 1698431365
transform 1 0 11648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__I
timestamp 1698431365
transform -1 0 16352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__I
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__I
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__A1
timestamp 1698431365
transform 1 0 12768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__A2
timestamp 1698431365
transform 1 0 10640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__B2
timestamp 1698431365
transform -1 0 12992 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__A2
timestamp 1698431365
transform -1 0 6160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__501__I
timestamp 1698431365
transform -1 0 9408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__I
timestamp 1698431365
transform -1 0 19040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__A2
timestamp 1698431365
transform 1 0 6944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__C2
timestamp 1698431365
transform -1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__A1
timestamp 1698431365
transform 1 0 15344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__I
timestamp 1698431365
transform -1 0 11760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__I
timestamp 1698431365
transform -1 0 12656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__I
timestamp 1698431365
transform 1 0 12320 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__I
timestamp 1698431365
transform 1 0 22064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__I
timestamp 1698431365
transform -1 0 7280 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__A1
timestamp 1698431365
transform 1 0 18032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__B1
timestamp 1698431365
transform 1 0 18928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__A2
timestamp 1698431365
transform 1 0 19376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__A3
timestamp 1698431365
transform 1 0 18928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__A3
timestamp 1698431365
transform -1 0 11536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__A1
timestamp 1698431365
transform 1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__A2
timestamp 1698431365
transform -1 0 10080 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__B1
timestamp 1698431365
transform 1 0 14672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__C2
timestamp 1698431365
transform 1 0 15120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__552__I
timestamp 1698431365
transform 1 0 13552 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__B2
timestamp 1698431365
transform 1 0 17920 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__C2
timestamp 1698431365
transform -1 0 15232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__559__A2
timestamp 1698431365
transform 1 0 14672 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__560__A2
timestamp 1698431365
transform 1 0 12768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__A2
timestamp 1698431365
transform 1 0 18592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__572__B1
timestamp 1698431365
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__C2
timestamp 1698431365
transform -1 0 14448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__583__A1
timestamp 1698431365
transform 1 0 10192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__I
timestamp 1698431365
transform -1 0 10416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__A2
timestamp 1698431365
transform -1 0 10864 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__B
timestamp 1698431365
transform -1 0 12320 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__587__A2
timestamp 1698431365
transform 1 0 22400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__A1
timestamp 1698431365
transform 1 0 23072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__A2
timestamp 1698431365
transform 1 0 22288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__595__A1
timestamp 1698431365
transform 1 0 21616 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__598__I
timestamp 1698431365
transform -1 0 12880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__A2
timestamp 1698431365
transform 1 0 22512 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__A2
timestamp 1698431365
transform 1 0 23296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__603__A2
timestamp 1698431365
transform 1 0 21616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__A2
timestamp 1698431365
transform 1 0 22400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__B
timestamp 1698431365
transform -1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__605__A1
timestamp 1698431365
transform 1 0 17808 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__614__I
timestamp 1698431365
transform 1 0 23408 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__615__A1
timestamp 1698431365
transform 1 0 24864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__616__C1
timestamp 1698431365
transform 1 0 9968 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__616__C2
timestamp 1698431365
transform 1 0 8400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__A2
timestamp 1698431365
transform 1 0 14560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__629__A1
timestamp 1698431365
transform -1 0 11312 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__629__B2
timestamp 1698431365
transform -1 0 11312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__633__A1
timestamp 1698431365
transform 1 0 14448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__634__A1
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__635__A1
timestamp 1698431365
transform 1 0 14000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__635__B1
timestamp 1698431365
transform -1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__641__A1
timestamp 1698431365
transform -1 0 15680 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__642__A1
timestamp 1698431365
transform -1 0 17472 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__645__I
timestamp 1698431365
transform 1 0 20720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__A1
timestamp 1698431365
transform 1 0 8064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__653__B1
timestamp 1698431365
transform 1 0 18480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__I
timestamp 1698431365
transform 1 0 22736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__659__I
timestamp 1698431365
transform -1 0 18704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__660__C
timestamp 1698431365
transform -1 0 23296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__662__B
timestamp 1698431365
transform -1 0 18032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__663__A1
timestamp 1698431365
transform 1 0 15456 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__665__A1
timestamp 1698431365
transform 1 0 16016 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__665__B
timestamp 1698431365
transform 1 0 16464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__671__I
timestamp 1698431365
transform -1 0 9408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__672__B1
timestamp 1698431365
transform -1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__673__A2
timestamp 1698431365
transform 1 0 19488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__B1
timestamp 1698431365
transform -1 0 15792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__B2
timestamp 1698431365
transform 1 0 16128 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__679__B2
timestamp 1698431365
transform -1 0 12320 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__682__A2
timestamp 1698431365
transform -1 0 8960 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__A3
timestamp 1698431365
transform -1 0 9968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__A4
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__692__A3
timestamp 1698431365
transform 1 0 20272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__694__A2
timestamp 1698431365
transform 1 0 22176 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__696__I
timestamp 1698431365
transform -1 0 11088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__B
timestamp 1698431365
transform 1 0 19152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__705__A4
timestamp 1698431365
transform -1 0 21168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__B2
timestamp 1698431365
transform 1 0 6832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__709__A2
timestamp 1698431365
transform -1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__709__B1
timestamp 1698431365
transform 1 0 21392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__A2
timestamp 1698431365
transform -1 0 20048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__A1
timestamp 1698431365
transform -1 0 22624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__A2
timestamp 1698431365
transform -1 0 23072 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__717__A1
timestamp 1698431365
transform 1 0 24528 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__720__A1
timestamp 1698431365
transform 1 0 24976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__732__A3
timestamp 1698431365
transform 1 0 24416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__734__A1
timestamp 1698431365
transform 1 0 26544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__A1
timestamp 1698431365
transform -1 0 19376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__747__A2
timestamp 1698431365
transform -1 0 19824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__750__C1
timestamp 1698431365
transform 1 0 7392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__751__A1
timestamp 1698431365
transform 1 0 22736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__751__A4
timestamp 1698431365
transform -1 0 23408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__753__A1
timestamp 1698431365
transform 1 0 10640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__756__A2
timestamp 1698431365
transform -1 0 7504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__761__A1
timestamp 1698431365
transform -1 0 8064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__769__A2
timestamp 1698431365
transform 1 0 23184 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__770__A2
timestamp 1698431365
transform 1 0 24304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 7280 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 15008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 7280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 3136 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 6832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 3584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 8064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 4480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 8176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 7728 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 4592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 1792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 2912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 2800 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 1792 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 1792 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 2016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 5712 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 3808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 6384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 3136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 2688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 2016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 2912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 2912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 2912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 2464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 2464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output44_I
timestamp 1698431365
transform 1 0 19936 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output50_I
timestamp 1698431365
transform 1 0 35952 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output51_I
timestamp 1698431365
transform -1 0 37520 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_8 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_12 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_28 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4480 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_32
timestamp 1698431365
transform 1 0 4928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698431365
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_8
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_12
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_28
timestamp 1698431365
transform 1 0 4480 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_32
timestamp 1698431365
transform 1 0 4928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_8
timestamp 1698431365
transform 1 0 2240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_12
timestamp 1698431365
transform 1 0 2688 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_44
timestamp 1698431365
transform 1 0 6272 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_60 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8064 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_68
timestamp 1698431365
transform 1 0 8960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698431365
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_8
timestamp 1698431365
transform 1 0 2240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_12
timestamp 1698431365
transform 1 0 2688 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_28
timestamp 1698431365
transform 1 0 4480 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698431365
transform 1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_8
timestamp 1698431365
transform 1 0 2240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_12
timestamp 1698431365
transform 1 0 2688 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_44
timestamp 1698431365
transform 1 0 6272 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_60
timestamp 1698431365
transform 1 0 8064 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698431365
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_8
timestamp 1698431365
transform 1 0 2240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_12
timestamp 1698431365
transform 1 0 2688 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_28
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_8
timestamp 1698431365
transform 1 0 2240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_12
timestamp 1698431365
transform 1 0 2688 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_44
timestamp 1698431365
transform 1 0 6272 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_60
timestamp 1698431365
transform 1 0 8064 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_68
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698431365
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1698431365
transform 1 0 2240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_12
timestamp 1698431365
transform 1 0 2688 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1698431365
transform 1 0 4480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698431365
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1698431365
transform 1 0 2240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_12
timestamp 1698431365
transform 1 0 2688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1698431365
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698431365
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_8
timestamp 1698431365
transform 1 0 2240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_12
timestamp 1698431365
transform 1 0 2688 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_44
timestamp 1698431365
transform 1 0 6272 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_60
timestamp 1698431365
transform 1 0 8064 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698431365
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_12
timestamp 1698431365
transform 1 0 2688 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1698431365
transform 1 0 4480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_8
timestamp 1698431365
transform 1 0 2240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_12
timestamp 1698431365
transform 1 0 2688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_16
timestamp 1698431365
transform 1 0 3136 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_48
timestamp 1698431365
transform 1 0 6720 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_64
timestamp 1698431365
transform 1 0 8512 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698431365
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_76
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_78
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_81
timestamp 1698431365
transform 1 0 10416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_87
timestamp 1698431365
transform 1 0 11088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_95
timestamp 1698431365
transform 1 0 11984 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_99
timestamp 1698431365
transform 1 0 12432 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_103
timestamp 1698431365
transform 1 0 12880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_107
timestamp 1698431365
transform 1 0 13328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_115
timestamp 1698431365
transform 1 0 14224 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_125
timestamp 1698431365
transform 1 0 15344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_129
timestamp 1698431365
transform 1 0 15792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_131
timestamp 1698431365
transform 1 0 16016 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_134
timestamp 1698431365
transform 1 0 16352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_146
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_154
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_158
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_190
timestamp 1698431365
transform 1 0 22624 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698431365
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698431365
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_8
timestamp 1698431365
transform 1 0 2240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_12
timestamp 1698431365
transform 1 0 2688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_16
timestamp 1698431365
transform 1 0 3136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_25
timestamp 1698431365
transform 1 0 4144 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_33
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_69
timestamp 1698431365
transform 1 0 9072 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_72
timestamp 1698431365
transform 1 0 9408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_74
timestamp 1698431365
transform 1 0 9632 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_77
timestamp 1698431365
transform 1 0 9968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_81
timestamp 1698431365
transform 1 0 10416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_85
timestamp 1698431365
transform 1 0 10864 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_89
timestamp 1698431365
transform 1 0 11312 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_93
timestamp 1698431365
transform 1 0 11760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_95
timestamp 1698431365
transform 1 0 11984 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_98
timestamp 1698431365
transform 1 0 12320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_102
timestamp 1698431365
transform 1 0 12768 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_129
timestamp 1698431365
transform 1 0 15792 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_131
timestamp 1698431365
transform 1 0 16016 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_142
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_160
timestamp 1698431365
transform 1 0 19264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_164
timestamp 1698431365
transform 1 0 19712 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_181
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_187
timestamp 1698431365
transform 1 0 22288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_191
timestamp 1698431365
transform 1 0 22736 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_223
timestamp 1698431365
transform 1 0 26320 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_14
timestamp 1698431365
transform 1 0 2912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_60
timestamp 1698431365
transform 1 0 8064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_95
timestamp 1698431365
transform 1 0 11984 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_101
timestamp 1698431365
transform 1 0 12656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_127
timestamp 1698431365
transform 1 0 15568 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_158
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_162
timestamp 1698431365
transform 1 0 19488 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_188
timestamp 1698431365
transform 1 0 22400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_192
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_196
timestamp 1698431365
transform 1 0 23296 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698431365
transform 1 0 24192 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698431365
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698431365
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_8
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_10
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_43
timestamp 1698431365
transform 1 0 6160 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_51
timestamp 1698431365
transform 1 0 7056 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_55
timestamp 1698431365
transform 1 0 7504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_115
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_117
timestamp 1698431365
transform 1 0 14448 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_136
timestamp 1698431365
transform 1 0 16576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_138
timestamp 1698431365
transform 1 0 16800 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_227
timestamp 1698431365
transform 1 0 26768 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_36
timestamp 1698431365
transform 1 0 5376 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_44
timestamp 1698431365
transform 1 0 6272 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_48
timestamp 1698431365
transform 1 0 6720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_50
timestamp 1698431365
transform 1 0 6944 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_85
timestamp 1698431365
transform 1 0 10864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_87
timestamp 1698431365
transform 1 0 11088 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_151
timestamp 1698431365
transform 1 0 18256 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_27
timestamp 1698431365
transform 1 0 4368 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_31
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_45
timestamp 1698431365
transform 1 0 6384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_47
timestamp 1698431365
transform 1 0 6608 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_80
timestamp 1698431365
transform 1 0 10304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_82
timestamp 1698431365
transform 1 0 10528 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_85
timestamp 1698431365
transform 1 0 10864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_115
timestamp 1698431365
transform 1 0 14224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_117
timestamp 1698431365
transform 1 0 14448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_129
timestamp 1698431365
transform 1 0 15792 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_140
timestamp 1698431365
transform 1 0 17024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_144
timestamp 1698431365
transform 1 0 17472 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_148
timestamp 1698431365
transform 1 0 17920 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_151
timestamp 1698431365
transform 1 0 18256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_179
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_224
timestamp 1698431365
transform 1 0 26432 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_10
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_20
timestamp 1698431365
transform 1 0 3584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_24
timestamp 1698431365
transform 1 0 4032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_26
timestamp 1698431365
transform 1 0 4256 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_43
timestamp 1698431365
transform 1 0 6160 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_51
timestamp 1698431365
transform 1 0 7056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_58
timestamp 1698431365
transform 1 0 7840 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_80
timestamp 1698431365
transform 1 0 10304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_122
timestamp 1698431365
transform 1 0 15008 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_154
timestamp 1698431365
transform 1 0 18592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_158
timestamp 1698431365
transform 1 0 19040 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_177
timestamp 1698431365
transform 1 0 21168 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_196
timestamp 1698431365
transform 1 0 23296 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_205
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_41
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_57
timestamp 1698431365
transform 1 0 7728 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_65
timestamp 1698431365
transform 1 0 8624 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_68
timestamp 1698431365
transform 1 0 8960 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_96
timestamp 1698431365
transform 1 0 12096 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_100
timestamp 1698431365
transform 1 0 12544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698431365
transform 1 0 15120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_127
timestamp 1698431365
transform 1 0 15568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_129
timestamp 1698431365
transform 1 0 15792 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_186
timestamp 1698431365
transform 1 0 22176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_190
timestamp 1698431365
transform 1 0 22624 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_194
timestamp 1698431365
transform 1 0 23072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_197
timestamp 1698431365
transform 1 0 23408 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_206
timestamp 1698431365
transform 1 0 24416 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_218
timestamp 1698431365
transform 1 0 25760 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_234
timestamp 1698431365
transform 1 0 27552 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698431365
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_14
timestamp 1698431365
transform 1 0 2912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_39
timestamp 1698431365
transform 1 0 5712 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_43
timestamp 1698431365
transform 1 0 6160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_47
timestamp 1698431365
transform 1 0 6608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_49
timestamp 1698431365
transform 1 0 6832 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_63
timestamp 1698431365
transform 1 0 8400 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_87
timestamp 1698431365
transform 1 0 11088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_100
timestamp 1698431365
transform 1 0 12544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_130
timestamp 1698431365
transform 1 0 15904 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_160
timestamp 1698431365
transform 1 0 19264 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_164
timestamp 1698431365
transform 1 0 19712 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_166
timestamp 1698431365
transform 1 0 19936 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_171
timestamp 1698431365
transform 1 0 20496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_186
timestamp 1698431365
transform 1 0 22176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_190
timestamp 1698431365
transform 1 0 22624 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_194
timestamp 1698431365
transform 1 0 23072 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_196
timestamp 1698431365
transform 1 0 23296 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_252
timestamp 1698431365
transform 1 0 29568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_268
timestamp 1698431365
transform 1 0 31360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698431365
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698431365
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_10
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698431365
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_53
timestamp 1698431365
transform 1 0 7280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_77
timestamp 1698431365
transform 1 0 9968 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_87
timestamp 1698431365
transform 1 0 11088 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_94
timestamp 1698431365
transform 1 0 11872 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_98
timestamp 1698431365
transform 1 0 12320 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_100
timestamp 1698431365
transform 1 0 12544 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_103
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_147
timestamp 1698431365
transform 1 0 17808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_151
timestamp 1698431365
transform 1 0 18256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_155
timestamp 1698431365
transform 1 0 18704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_164
timestamp 1698431365
transform 1 0 19712 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_188
timestamp 1698431365
transform 1 0 22400 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_194
timestamp 1698431365
transform 1 0 23072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_198
timestamp 1698431365
transform 1 0 23520 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_4
timestamp 1698431365
transform 1 0 1792 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_67
timestamp 1698431365
transform 1 0 8848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_88
timestamp 1698431365
transform 1 0 11200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_111
timestamp 1698431365
transform 1 0 13776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_115
timestamp 1698431365
transform 1 0 14224 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_131
timestamp 1698431365
transform 1 0 16016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_135
timestamp 1698431365
transform 1 0 16464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_137
timestamp 1698431365
transform 1 0 16688 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_194
timestamp 1698431365
transform 1 0 23072 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_198
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_214
timestamp 1698431365
transform 1 0 25312 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_259
timestamp 1698431365
transform 1 0 30352 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_275
timestamp 1698431365
transform 1 0 32144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698431365
transform 1 0 40096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_8
timestamp 1698431365
transform 1 0 2240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_10
timestamp 1698431365
transform 1 0 2464 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_49
timestamp 1698431365
transform 1 0 6832 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_53
timestamp 1698431365
transform 1 0 7280 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_56
timestamp 1698431365
transform 1 0 7616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_95
timestamp 1698431365
transform 1 0 11984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_102
timestamp 1698431365
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698431365
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_127
timestamp 1698431365
transform 1 0 15568 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_167
timestamp 1698431365
transform 1 0 20048 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_179
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_193
timestamp 1698431365
transform 1 0 22960 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_197
timestamp 1698431365
transform 1 0 23408 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_205
timestamp 1698431365
transform 1 0 24304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_209
timestamp 1698431365
transform 1 0 24752 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_6
timestamp 1698431365
transform 1 0 2016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_10
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_14
timestamp 1698431365
transform 1 0 2912 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_18
timestamp 1698431365
transform 1 0 3360 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_45
timestamp 1698431365
transform 1 0 6384 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_51
timestamp 1698431365
transform 1 0 7056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_74
timestamp 1698431365
transform 1 0 9632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_90
timestamp 1698431365
transform 1 0 11424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_92
timestamp 1698431365
transform 1 0 11648 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_151
timestamp 1698431365
transform 1 0 18256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_194
timestamp 1698431365
transform 1 0 23072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_196
timestamp 1698431365
transform 1 0 23296 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_248
timestamp 1698431365
transform 1 0 29120 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_8
timestamp 1698431365
transform 1 0 2240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_12
timestamp 1698431365
transform 1 0 2688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_16
timestamp 1698431365
transform 1 0 3136 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_20
timestamp 1698431365
transform 1 0 3584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_22
timestamp 1698431365
transform 1 0 3808 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_50
timestamp 1698431365
transform 1 0 6944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_111
timestamp 1698431365
transform 1 0 13776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_161
timestamp 1698431365
transform 1 0 19376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698431365
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_219
timestamp 1698431365
transform 1 0 25872 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_240
timestamp 1698431365
transform 1 0 28224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_14
timestamp 1698431365
transform 1 0 2912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_62
timestamp 1698431365
transform 1 0 8288 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_81
timestamp 1698431365
transform 1 0 10416 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_119
timestamp 1698431365
transform 1 0 14672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698431365
transform 1 0 16688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_179
timestamp 1698431365
transform 1 0 21392 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_183
timestamp 1698431365
transform 1 0 21840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_187
timestamp 1698431365
transform 1 0 22288 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_193
timestamp 1698431365
transform 1 0 22960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_197
timestamp 1698431365
transform 1 0 23408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_244
timestamp 1698431365
transform 1 0 28672 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698431365
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_8
timestamp 1698431365
transform 1 0 2240 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_59
timestamp 1698431365
transform 1 0 7952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_61
timestamp 1698431365
transform 1 0 8176 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_115
timestamp 1698431365
transform 1 0 14224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_168
timestamp 1698431365
transform 1 0 20160 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_235
timestamp 1698431365
transform 1 0 27664 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698431365
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_4
timestamp 1698431365
transform 1 0 1792 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_27
timestamp 1698431365
transform 1 0 4368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_61
timestamp 1698431365
transform 1 0 8176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_76
timestamp 1698431365
transform 1 0 9856 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_163
timestamp 1698431365
transform 1 0 19600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_182
timestamp 1698431365
transform 1 0 21728 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_186
timestamp 1698431365
transform 1 0 22176 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_243
timestamp 1698431365
transform 1 0 28560 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_275
timestamp 1698431365
transform 1 0 32144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_60
timestamp 1698431365
transform 1 0 8064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_117
timestamp 1698431365
transform 1 0 14448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_157
timestamp 1698431365
transform 1 0 18928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_161
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_167
timestamp 1698431365
transform 1 0 20048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_184
timestamp 1698431365
transform 1 0 21952 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_190
timestamp 1698431365
transform 1 0 22624 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_196
timestamp 1698431365
transform 1 0 23296 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698431365
transform 1 0 27104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698431365
transform 1 0 28000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_59
timestamp 1698431365
transform 1 0 7952 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_104
timestamp 1698431365
transform 1 0 12992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_106
timestamp 1698431365
transform 1 0 13216 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_123
timestamp 1698431365
transform 1 0 15120 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_125
timestamp 1698431365
transform 1 0 15344 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_137
timestamp 1698431365
transform 1 0 16688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_160
timestamp 1698431365
transform 1 0 19264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_162
timestamp 1698431365
transform 1 0 19488 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_171
timestamp 1698431365
transform 1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_175
timestamp 1698431365
transform 1 0 20944 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_183
timestamp 1698431365
transform 1 0 21840 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_187
timestamp 1698431365
transform 1 0 22288 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_190
timestamp 1698431365
transform 1 0 22624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_205
timestamp 1698431365
transform 1 0 24304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_223
timestamp 1698431365
transform 1 0 26320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_227
timestamp 1698431365
transform 1 0 26768 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_259
timestamp 1698431365
transform 1 0 30352 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_275
timestamp 1698431365
transform 1 0 32144 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698431365
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_8
timestamp 1698431365
transform 1 0 2240 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_12
timestamp 1698431365
transform 1 0 2688 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_29
timestamp 1698431365
transform 1 0 4592 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_58
timestamp 1698431365
transform 1 0 7840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_126
timestamp 1698431365
transform 1 0 15456 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_138
timestamp 1698431365
transform 1 0 16800 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_145
timestamp 1698431365
transform 1 0 17584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_149
timestamp 1698431365
transform 1 0 18032 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_156
timestamp 1698431365
transform 1 0 18816 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_189
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_224
timestamp 1698431365
transform 1 0 26432 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_240
timestamp 1698431365
transform 1 0 28224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_24
timestamp 1698431365
transform 1 0 4032 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_63
timestamp 1698431365
transform 1 0 8400 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_82
timestamp 1698431365
transform 1 0 10528 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_101
timestamp 1698431365
transform 1 0 12656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_103
timestamp 1698431365
transform 1 0 12880 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_129
timestamp 1698431365
transform 1 0 15792 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_133
timestamp 1698431365
transform 1 0 16240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_137
timestamp 1698431365
transform 1 0 16688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_146
timestamp 1698431365
transform 1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_163
timestamp 1698431365
transform 1 0 19600 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_171
timestamp 1698431365
transform 1 0 20496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_188
timestamp 1698431365
transform 1 0 22400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_192
timestamp 1698431365
transform 1 0 22848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_194
timestamp 1698431365
transform 1 0 23072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_200
timestamp 1698431365
transform 1 0 23744 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_208
timestamp 1698431365
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_8
timestamp 1698431365
transform 1 0 2240 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_26
timestamp 1698431365
transform 1 0 4256 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_81
timestamp 1698431365
transform 1 0 10416 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_85
timestamp 1698431365
transform 1 0 10864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_87
timestamp 1698431365
transform 1 0 11088 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_102
timestamp 1698431365
transform 1 0 12768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_158
timestamp 1698431365
transform 1 0 19040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_168
timestamp 1698431365
transform 1 0 20160 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_172
timestamp 1698431365
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_189
timestamp 1698431365
transform 1 0 22512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_191
timestamp 1698431365
transform 1 0 22736 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_197
timestamp 1698431365
transform 1 0 23408 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_209
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_18
timestamp 1698431365
transform 1 0 3360 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_50
timestamp 1698431365
transform 1 0 6944 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_54
timestamp 1698431365
transform 1 0 7392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_56
timestamp 1698431365
transform 1 0 7616 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_65
timestamp 1698431365
transform 1 0 8624 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_113
timestamp 1698431365
transform 1 0 14000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_117
timestamp 1698431365
transform 1 0 14448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_121
timestamp 1698431365
transform 1 0 14896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_125
timestamp 1698431365
transform 1 0 15344 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_132
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_159
timestamp 1698431365
transform 1 0 19152 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_167
timestamp 1698431365
transform 1 0 20048 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_173
timestamp 1698431365
transform 1 0 20720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_192
timestamp 1698431365
transform 1 0 22848 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_218
timestamp 1698431365
transform 1 0 25760 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_250
timestamp 1698431365
transform 1 0 29344 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_266
timestamp 1698431365
transform 1 0 31136 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_274
timestamp 1698431365
transform 1 0 32032 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_278
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698431365
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698431365
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_4
timestamp 1698431365
transform 1 0 1792 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_90
timestamp 1698431365
transform 1 0 11424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_100
timestamp 1698431365
transform 1 0 12544 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_117
timestamp 1698431365
transform 1 0 14448 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_121
timestamp 1698431365
transform 1 0 14896 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_146
timestamp 1698431365
transform 1 0 17696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_150
timestamp 1698431365
transform 1 0 18144 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_166
timestamp 1698431365
transform 1 0 19936 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_185
timestamp 1698431365
transform 1 0 22064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_208
timestamp 1698431365
transform 1 0 24640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_212
timestamp 1698431365
transform 1 0 25088 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_65
timestamp 1698431365
transform 1 0 8624 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_74
timestamp 1698431365
transform 1 0 9632 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_100
timestamp 1698431365
transform 1 0 12544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_104
timestamp 1698431365
transform 1 0 12992 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_116
timestamp 1698431365
transform 1 0 14336 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_120
timestamp 1698431365
transform 1 0 14784 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_122
timestamp 1698431365
transform 1 0 15008 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_129
timestamp 1698431365
transform 1 0 15792 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_150
timestamp 1698431365
transform 1 0 18144 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_154
timestamp 1698431365
transform 1 0 18592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_156
timestamp 1698431365
transform 1 0 18816 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_159
timestamp 1698431365
transform 1 0 19152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_184
timestamp 1698431365
transform 1 0 21952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_188
timestamp 1698431365
transform 1 0 22400 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_190
timestamp 1698431365
transform 1 0 22624 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_203
timestamp 1698431365
transform 1 0 24080 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_207
timestamp 1698431365
transform 1 0 24528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698431365
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698431365
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_43
timestamp 1698431365
transform 1 0 6160 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_58
timestamp 1698431365
transform 1 0 7840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_60
timestamp 1698431365
transform 1 0 8064 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_87
timestamp 1698431365
transform 1 0 11088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_97
timestamp 1698431365
transform 1 0 12208 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_115
timestamp 1698431365
transform 1 0 14224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_193
timestamp 1698431365
transform 1 0 22960 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_199
timestamp 1698431365
transform 1 0 23632 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_231
timestamp 1698431365
transform 1 0 27216 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_239
timestamp 1698431365
transform 1 0 28112 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_243
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_80
timestamp 1698431365
transform 1 0 10304 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_88
timestamp 1698431365
transform 1 0 11200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_90
timestamp 1698431365
transform 1 0 11424 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_101
timestamp 1698431365
transform 1 0 12656 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_105
timestamp 1698431365
transform 1 0 13104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_107
timestamp 1698431365
transform 1 0 13328 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_116
timestamp 1698431365
transform 1 0 14336 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_146
timestamp 1698431365
transform 1 0 17696 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_152
timestamp 1698431365
transform 1 0 18368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_156
timestamp 1698431365
transform 1 0 18816 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_168
timestamp 1698431365
transform 1 0 20160 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_200
timestamp 1698431365
transform 1 0 23744 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_6
timestamp 1698431365
transform 1 0 2016 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_51
timestamp 1698431365
transform 1 0 7056 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_55
timestamp 1698431365
transform 1 0 7504 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_57
timestamp 1698431365
transform 1 0 7728 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_141
timestamp 1698431365
transform 1 0 17136 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_14
timestamp 1698431365
transform 1 0 2912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_18
timestamp 1698431365
transform 1 0 3360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_22
timestamp 1698431365
transform 1 0 3808 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_28
timestamp 1698431365
transform 1 0 4480 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_47
timestamp 1698431365
transform 1 0 6608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_51
timestamp 1698431365
transform 1 0 7056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_55
timestamp 1698431365
transform 1 0 7504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_63
timestamp 1698431365
transform 1 0 8400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_67
timestamp 1698431365
transform 1 0 8848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_135
timestamp 1698431365
transform 1 0 16464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_150
timestamp 1698431365
transform 1 0 18144 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_182
timestamp 1698431365
transform 1 0 21728 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_198
timestamp 1698431365
transform 1 0 23520 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698431365
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_8
timestamp 1698431365
transform 1 0 2240 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_27
timestamp 1698431365
transform 1 0 4368 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_47
timestamp 1698431365
transform 1 0 6608 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_58
timestamp 1698431365
transform 1 0 7840 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_130
timestamp 1698431365
transform 1 0 15904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_146
timestamp 1698431365
transform 1 0 17696 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_162
timestamp 1698431365
transform 1 0 19488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_170
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_22
timestamp 1698431365
transform 1 0 3808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_24
timestamp 1698431365
transform 1 0 4032 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_67
timestamp 1698431365
transform 1 0 8848 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_69
timestamp 1698431365
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_126
timestamp 1698431365
transform 1 0 15456 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_134
timestamp 1698431365
transform 1 0 16352 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_138
timestamp 1698431365
transform 1 0 16800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_158
timestamp 1698431365
transform 1 0 19040 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_160
timestamp 1698431365
transform 1 0 19264 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_187
timestamp 1698431365
transform 1 0 22288 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698431365
transform 1 0 23856 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698431365
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_214
timestamp 1698431365
transform 1 0 25312 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_247
timestamp 1698431365
transform 1 0 29008 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_298
timestamp 1698431365
transform 1 0 34720 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_306
timestamp 1698431365
transform 1 0 35616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_308
timestamp 1698431365
transform 1 0 35840 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_311
timestamp 1698431365
transform 1 0 36176 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_319
timestamp 1698431365
transform 1 0 37072 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_14
timestamp 1698431365
transform 1 0 2912 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_36
timestamp 1698431365
transform 1 0 5376 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_38
timestamp 1698431365
transform 1 0 5600 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_51
timestamp 1698431365
transform 1 0 7056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_55
timestamp 1698431365
transform 1 0 7504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_59
timestamp 1698431365
transform 1 0 7952 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_63
timestamp 1698431365
transform 1 0 8400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_65
timestamp 1698431365
transform 1 0 8624 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_70
timestamp 1698431365
transform 1 0 9184 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_79
timestamp 1698431365
transform 1 0 10192 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_120
timestamp 1698431365
transform 1 0 14784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_124
timestamp 1698431365
transform 1 0 15232 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_132
timestamp 1698431365
transform 1 0 16128 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_164
timestamp 1698431365
transform 1 0 19712 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_168
timestamp 1698431365
transform 1 0 20160 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698431365
transform 1 0 20608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_180
timestamp 1698431365
transform 1 0 21504 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_196
timestamp 1698431365
transform 1 0 23296 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698431365
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698431365
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_240
timestamp 1698431365
transform 1 0 28224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_274
timestamp 1698431365
transform 1 0 32032 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_278
timestamp 1698431365
transform 1 0 32480 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_308
timestamp 1698431365
transform 1 0 35840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_310
timestamp 1698431365
transform 1 0 36064 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_337
timestamp 1698431365
transform 1 0 39088 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_339
timestamp 1698431365
transform 1 0 39312 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698431365
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698431365
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698431365
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2
timestamp 1698431365
transform 1 0 9296 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 14112 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform 1 0 2128 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input6
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698431365
transform -1 0 2912 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 5152 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 2240 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 4480 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 3136 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input17
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 2240 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 2240 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 2240 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input29
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 2240 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input36
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input40
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform -1 0 2240 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output44 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19712 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output45
timestamp 1698431365
transform -1 0 22288 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output46
timestamp 1698431365
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output47
timestamp 1698431365
transform 1 0 26096 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output48
timestamp 1698431365
transform 1 0 28896 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output49
timestamp 1698431365
transform 1 0 32704 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output50
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51
timestamp 1698431365
transform 1 0 37520 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698431365
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698431365
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698431365
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698431365
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698431365
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698431365
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698431365
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698431365
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698431365
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal2 s 15904 41200 16016 42000 0 FreeSans 448 90 0 0 bus_out[0]
port 0 nsew signal tristate
flabel metal2 s 19264 41200 19376 42000 0 FreeSans 448 90 0 0 bus_out[1]
port 1 nsew signal tristate
flabel metal2 s 22624 41200 22736 42000 0 FreeSans 448 90 0 0 bus_out[2]
port 2 nsew signal tristate
flabel metal2 s 25984 41200 26096 42000 0 FreeSans 448 90 0 0 bus_out[3]
port 3 nsew signal tristate
flabel metal2 s 29344 41200 29456 42000 0 FreeSans 448 90 0 0 bus_out[4]
port 4 nsew signal tristate
flabel metal2 s 32704 41200 32816 42000 0 FreeSans 448 90 0 0 bus_out[5]
port 5 nsew signal tristate
flabel metal2 s 36064 41200 36176 42000 0 FreeSans 448 90 0 0 bus_out[6]
port 6 nsew signal tristate
flabel metal2 s 39424 41200 39536 42000 0 FreeSans 448 90 0 0 bus_out[7]
port 7 nsew signal tristate
flabel metal2 s 5824 41200 5936 42000 0 FreeSans 448 90 0 0 cs_port[0]
port 8 nsew signal input
flabel metal2 s 9184 41200 9296 42000 0 FreeSans 448 90 0 0 cs_port[1]
port 9 nsew signal input
flabel metal2 s 12544 41200 12656 42000 0 FreeSans 448 90 0 0 cs_port[2]
port 10 nsew signal input
flabel metal3 s 0 32032 800 32144 0 FreeSans 448 0 0 0 last_addr[0]
port 11 nsew signal input
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 last_addr[1]
port 12 nsew signal input
flabel metal3 s 0 33824 800 33936 0 FreeSans 448 0 0 0 last_addr[2]
port 13 nsew signal input
flabel metal3 s 0 34720 800 34832 0 FreeSans 448 0 0 0 last_addr[3]
port 14 nsew signal input
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 last_addr[4]
port 15 nsew signal input
flabel metal3 s 0 36512 800 36624 0 FreeSans 448 0 0 0 last_addr[5]
port 16 nsew signal input
flabel metal3 s 0 37408 800 37520 0 FreeSans 448 0 0 0 last_addr[6]
port 17 nsew signal input
flabel metal3 s 0 38304 800 38416 0 FreeSans 448 0 0 0 last_addr[7]
port 18 nsew signal input
flabel metal3 s 0 17696 800 17808 0 FreeSans 448 0 0 0 ram_end[0]
port 19 nsew signal input
flabel metal3 s 0 26656 800 26768 0 FreeSans 448 0 0 0 ram_end[10]
port 20 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 ram_end[11]
port 21 nsew signal input
flabel metal3 s 0 28448 800 28560 0 FreeSans 448 0 0 0 ram_end[12]
port 22 nsew signal input
flabel metal3 s 0 29344 800 29456 0 FreeSans 448 0 0 0 ram_end[13]
port 23 nsew signal input
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 ram_end[14]
port 24 nsew signal input
flabel metal3 s 0 31136 800 31248 0 FreeSans 448 0 0 0 ram_end[15]
port 25 nsew signal input
flabel metal3 s 0 18592 800 18704 0 FreeSans 448 0 0 0 ram_end[1]
port 26 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 ram_end[2]
port 27 nsew signal input
flabel metal3 s 0 20384 800 20496 0 FreeSans 448 0 0 0 ram_end[3]
port 28 nsew signal input
flabel metal3 s 0 21280 800 21392 0 FreeSans 448 0 0 0 ram_end[4]
port 29 nsew signal input
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 ram_end[5]
port 30 nsew signal input
flabel metal3 s 0 23072 800 23184 0 FreeSans 448 0 0 0 ram_end[6]
port 31 nsew signal input
flabel metal3 s 0 23968 800 24080 0 FreeSans 448 0 0 0 ram_end[7]
port 32 nsew signal input
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 ram_end[8]
port 33 nsew signal input
flabel metal3 s 0 25760 800 25872 0 FreeSans 448 0 0 0 ram_end[9]
port 34 nsew signal input
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 ram_start[0]
port 35 nsew signal input
flabel metal3 s 0 12320 800 12432 0 FreeSans 448 0 0 0 ram_start[10]
port 36 nsew signal input
flabel metal3 s 0 13216 800 13328 0 FreeSans 448 0 0 0 ram_start[11]
port 37 nsew signal input
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 ram_start[12]
port 38 nsew signal input
flabel metal3 s 0 15008 800 15120 0 FreeSans 448 0 0 0 ram_start[13]
port 39 nsew signal input
flabel metal3 s 0 15904 800 16016 0 FreeSans 448 0 0 0 ram_start[14]
port 40 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 ram_start[15]
port 41 nsew signal input
flabel metal3 s 0 4256 800 4368 0 FreeSans 448 0 0 0 ram_start[1]
port 42 nsew signal input
flabel metal3 s 0 5152 800 5264 0 FreeSans 448 0 0 0 ram_start[2]
port 43 nsew signal input
flabel metal3 s 0 6048 800 6160 0 FreeSans 448 0 0 0 ram_start[3]
port 44 nsew signal input
flabel metal3 s 0 6944 800 7056 0 FreeSans 448 0 0 0 ram_start[4]
port 45 nsew signal input
flabel metal3 s 0 7840 800 7952 0 FreeSans 448 0 0 0 ram_start[5]
port 46 nsew signal input
flabel metal3 s 0 8736 800 8848 0 FreeSans 448 0 0 0 ram_start[6]
port 47 nsew signal input
flabel metal3 s 0 9632 800 9744 0 FreeSans 448 0 0 0 ram_start[7]
port 48 nsew signal input
flabel metal3 s 0 10528 800 10640 0 FreeSans 448 0 0 0 ram_start[8]
port 49 nsew signal input
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 ram_start[9]
port 50 nsew signal input
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 51 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 51 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 52 nsew ground bidirectional
flabel metal2 s 2464 41200 2576 42000 0 FreeSans 448 90 0 0 wb_clk_i
port 53 nsew signal input
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal3 21056 25256 21056 25256 0 _000_
rlabel metal2 7448 31584 7448 31584 0 _001_
rlabel metal2 5656 31248 5656 31248 0 _002_
rlabel metal3 9240 30296 9240 30296 0 _003_
rlabel metal2 11032 19992 11032 19992 0 _004_
rlabel metal3 18928 23576 18928 23576 0 _005_
rlabel metal3 13048 13832 13048 13832 0 _006_
rlabel metal2 15176 14224 15176 14224 0 _007_
rlabel metal2 14728 13944 14728 13944 0 _008_
rlabel metal2 19376 16184 19376 16184 0 _009_
rlabel metal2 20720 17752 20720 17752 0 _010_
rlabel metal3 5768 24808 5768 24808 0 _011_
rlabel metal2 4536 24696 4536 24696 0 _012_
rlabel metal2 5992 25088 5992 25088 0 _013_
rlabel metal2 5096 25536 5096 25536 0 _014_
rlabel metal2 10248 23184 10248 23184 0 _015_
rlabel metal2 10136 24080 10136 24080 0 _016_
rlabel metal2 18424 25424 18424 25424 0 _017_
rlabel via2 10024 37128 10024 37128 0 _018_
rlabel metal2 13160 38080 13160 38080 0 _019_
rlabel metal2 16128 35784 16128 35784 0 _020_
rlabel metal2 16296 33432 16296 33432 0 _021_
rlabel metal2 14840 27440 14840 27440 0 _022_
rlabel metal2 16632 31528 16632 31528 0 _023_
rlabel metal3 12936 23128 12936 23128 0 _024_
rlabel metal2 19544 23184 19544 23184 0 _025_
rlabel metal3 15512 11592 15512 11592 0 _026_
rlabel metal2 7784 36008 7784 36008 0 _027_
rlabel metal2 9352 14868 9352 14868 0 _028_
rlabel metal3 13888 29400 13888 29400 0 _029_
rlabel metal3 9408 21448 9408 21448 0 _030_
rlabel metal2 4536 29904 4536 29904 0 _031_
rlabel metal3 5936 30184 5936 30184 0 _032_
rlabel metal3 5320 33432 5320 33432 0 _033_
rlabel metal3 13328 13944 13328 13944 0 _034_
rlabel metal2 16408 15568 16408 15568 0 _035_
rlabel metal3 8568 30968 8568 30968 0 _036_
rlabel metal3 15344 26824 15344 26824 0 _037_
rlabel metal2 13832 23968 13832 23968 0 _038_
rlabel metal2 18536 19264 18536 19264 0 _039_
rlabel metal2 8344 17080 8344 17080 0 _040_
rlabel metal2 23800 17136 23800 17136 0 _041_
rlabel metal3 13048 33992 13048 33992 0 _042_
rlabel metal2 15792 13944 15792 13944 0 _043_
rlabel metal2 15848 22350 15848 22350 0 _044_
rlabel metal2 8120 17360 8120 17360 0 _045_
rlabel metal2 6440 22736 6440 22736 0 _046_
rlabel metal3 2968 26488 2968 26488 0 _047_
rlabel metal3 5040 25368 5040 25368 0 _048_
rlabel metal2 8568 24248 8568 24248 0 _049_
rlabel metal2 5152 16072 5152 16072 0 _050_
rlabel metal2 3584 14504 3584 14504 0 _051_
rlabel metal2 3696 15400 3696 15400 0 _052_
rlabel metal2 11312 14616 11312 14616 0 _053_
rlabel metal2 15176 16800 15176 16800 0 _054_
rlabel metal2 10472 27832 10472 27832 0 _055_
rlabel metal2 9464 19208 9464 19208 0 _056_
rlabel metal2 9016 16408 9016 16408 0 _057_
rlabel metal2 7336 17920 7336 17920 0 _058_
rlabel metal2 5768 27776 5768 27776 0 _059_
rlabel metal2 22568 27608 22568 27608 0 _060_
rlabel metal2 3752 20888 3752 20888 0 _061_
rlabel metal2 4312 21280 4312 21280 0 _062_
rlabel metal2 5992 23016 5992 23016 0 _063_
rlabel metal2 5880 21896 5880 21896 0 _064_
rlabel metal2 2968 22064 2968 22064 0 _065_
rlabel metal2 3304 21168 3304 21168 0 _066_
rlabel metal2 9912 19992 9912 19992 0 _067_
rlabel metal2 16576 32312 16576 32312 0 _068_
rlabel metal2 17360 25928 17360 25928 0 _069_
rlabel metal2 18648 14840 18648 14840 0 _070_
rlabel metal2 5880 24248 5880 24248 0 _071_
rlabel metal3 5152 23800 5152 23800 0 _072_
rlabel metal2 6216 21280 6216 21280 0 _073_
rlabel metal3 7504 29512 7504 29512 0 _074_
rlabel metal2 1960 17136 1960 17136 0 _075_
rlabel metal2 7224 20272 7224 20272 0 _076_
rlabel metal2 21896 22456 21896 22456 0 _077_
rlabel metal2 18368 18648 18368 18648 0 _078_
rlabel metal2 10472 30464 10472 30464 0 _079_
rlabel metal2 11704 14672 11704 14672 0 _080_
rlabel metal2 11032 16800 11032 16800 0 _081_
rlabel metal3 13048 15288 13048 15288 0 _082_
rlabel metal2 16408 16408 16408 16408 0 _083_
rlabel metal3 17976 18536 17976 18536 0 _084_
rlabel metal2 18200 19936 18200 19936 0 _085_
rlabel metal2 20384 20216 20384 20216 0 _086_
rlabel metal2 11032 18704 11032 18704 0 _087_
rlabel metal2 10584 20888 10584 20888 0 _088_
rlabel metal2 20216 19488 20216 19488 0 _089_
rlabel metal2 18648 24640 18648 24640 0 _090_
rlabel metal2 16408 35672 16408 35672 0 _091_
rlabel metal3 17024 22344 17024 22344 0 _092_
rlabel metal3 9128 29400 9128 29400 0 _093_
rlabel metal2 18648 29120 18648 29120 0 _094_
rlabel metal2 19992 24640 19992 24640 0 _095_
rlabel metal2 15288 36624 15288 36624 0 _096_
rlabel metal2 15400 32228 15400 32228 0 _097_
rlabel metal2 16296 31920 16296 31920 0 _098_
rlabel metal2 19432 26264 19432 26264 0 _099_
rlabel metal2 15400 31696 15400 31696 0 _100_
rlabel metal2 11592 17248 11592 17248 0 _101_
rlabel metal2 10024 19152 10024 19152 0 _102_
rlabel metal2 20272 21000 20272 21000 0 _103_
rlabel metal2 20664 21616 20664 21616 0 _104_
rlabel metal3 17248 33208 17248 33208 0 _105_
rlabel metal2 22120 14784 22120 14784 0 _106_
rlabel metal3 20720 31864 20720 31864 0 _107_
rlabel metal2 20888 14448 20888 14448 0 _108_
rlabel metal2 12152 31640 12152 31640 0 _109_
rlabel metal2 18088 25648 18088 25648 0 _110_
rlabel metal3 7224 25256 7224 25256 0 _111_
rlabel metal2 7336 25424 7336 25424 0 _112_
rlabel metal2 7672 25760 7672 25760 0 _113_
rlabel metal2 13048 31472 13048 31472 0 _114_
rlabel metal2 25368 29176 25368 29176 0 _115_
rlabel metal2 28728 21280 28728 21280 0 _116_
rlabel metal2 22344 21616 22344 21616 0 _117_
rlabel metal2 15624 25480 15624 25480 0 _118_
rlabel metal2 16520 30632 16520 30632 0 _119_
rlabel metal2 13888 34104 13888 34104 0 _120_
rlabel metal2 15736 32704 15736 32704 0 _121_
rlabel metal2 16464 33320 16464 33320 0 _122_
rlabel metal2 16520 31332 16520 31332 0 _123_
rlabel metal3 19768 30856 19768 30856 0 _124_
rlabel metal2 17080 33376 17080 33376 0 _125_
rlabel metal2 17304 32984 17304 32984 0 _126_
rlabel metal3 16968 33096 16968 33096 0 _127_
rlabel metal2 17808 33320 17808 33320 0 _128_
rlabel metal3 18144 30968 18144 30968 0 _129_
rlabel metal2 21672 25424 21672 25424 0 _130_
rlabel metal3 20496 17080 20496 17080 0 _131_
rlabel metal2 16632 28784 16632 28784 0 _132_
rlabel metal2 16968 22904 16968 22904 0 _133_
rlabel metal2 16856 21392 16856 21392 0 _134_
rlabel metal2 9576 22400 9576 22400 0 _135_
rlabel metal2 9912 15624 9912 15624 0 _136_
rlabel metal2 17864 20384 17864 20384 0 _137_
rlabel metal2 23800 22736 23800 22736 0 _138_
rlabel metal2 15344 28616 15344 28616 0 _139_
rlabel metal3 15764 23800 15764 23800 0 _140_
rlabel metal2 17416 24136 17416 24136 0 _141_
rlabel metal3 15960 25592 15960 25592 0 _142_
rlabel metal2 11592 19544 11592 19544 0 _143_
rlabel metal2 27048 24024 27048 24024 0 _144_
rlabel metal2 15176 33432 15176 33432 0 _145_
rlabel metal2 24136 27888 24136 27888 0 _146_
rlabel metal2 28392 23072 28392 23072 0 _147_
rlabel metal2 23688 23632 23688 23632 0 _148_
rlabel metal2 12264 16016 12264 16016 0 _149_
rlabel metal2 11704 15680 11704 15680 0 _150_
rlabel metal3 12152 16072 12152 16072 0 _151_
rlabel metal2 12824 15456 12824 15456 0 _152_
rlabel metal3 24024 18816 24024 18816 0 _153_
rlabel metal2 24080 22344 24080 22344 0 _154_
rlabel metal2 11480 29288 11480 29288 0 _155_
rlabel metal2 23576 27384 23576 27384 0 _156_
rlabel metal2 16968 21280 16968 21280 0 _157_
rlabel metal2 12824 27328 12824 27328 0 _158_
rlabel metal2 28392 25872 28392 25872 0 _159_
rlabel metal2 23912 24976 23912 24976 0 _160_
rlabel metal2 22680 23016 22680 23016 0 _161_
rlabel metal2 22904 22064 22904 22064 0 _162_
rlabel metal3 22344 14392 22344 14392 0 _163_
rlabel metal2 22008 14784 22008 14784 0 _164_
rlabel metal2 22680 21672 22680 21672 0 _165_
rlabel metal2 8792 26628 8792 26628 0 _166_
rlabel metal2 24472 17752 24472 17752 0 _167_
rlabel metal2 24136 18032 24136 18032 0 _168_
rlabel metal3 24248 24696 24248 24696 0 _169_
rlabel metal2 20328 28560 20328 28560 0 _170_
rlabel metal3 19824 28504 19824 28504 0 _171_
rlabel metal3 21056 26824 21056 26824 0 _172_
rlabel metal2 21336 33320 21336 33320 0 _173_
rlabel metal2 20216 24920 20216 24920 0 _174_
rlabel metal3 19768 25424 19768 25424 0 _175_
rlabel metal2 19656 26264 19656 26264 0 _176_
rlabel metal2 21448 27944 21448 27944 0 _177_
rlabel metal2 21560 26656 21560 26656 0 _178_
rlabel metal3 24360 31080 24360 31080 0 _179_
rlabel metal2 23800 29736 23800 29736 0 _180_
rlabel metal2 23352 27440 23352 27440 0 _181_
rlabel metal2 23184 27384 23184 27384 0 _182_
rlabel metal2 22512 21560 22512 21560 0 _183_
rlabel metal2 18648 25760 18648 25760 0 _184_
rlabel metal2 12824 26180 12824 26180 0 _185_
rlabel metal2 17304 24472 17304 24472 0 _186_
rlabel metal3 11424 24024 11424 24024 0 _187_
rlabel metal2 4368 19096 4368 19096 0 _188_
rlabel metal3 6160 16744 6160 16744 0 _189_
rlabel metal3 11816 18200 11816 18200 0 _190_
rlabel metal2 16856 18256 16856 18256 0 _191_
rlabel metal3 24696 15008 24696 15008 0 _192_
rlabel metal3 15680 16856 15680 16856 0 _193_
rlabel metal2 12600 17192 12600 17192 0 _194_
rlabel metal2 15288 16352 15288 16352 0 _195_
rlabel metal2 16296 17416 16296 17416 0 _196_
rlabel metal2 6552 25312 6552 25312 0 _197_
rlabel metal2 17752 25088 17752 25088 0 _198_
rlabel metal3 13608 20888 13608 20888 0 _199_
rlabel metal2 15960 21000 15960 21000 0 _200_
rlabel metal2 3080 19544 3080 19544 0 _201_
rlabel metal2 4144 17416 4144 17416 0 _202_
rlabel metal2 2912 15176 2912 15176 0 _203_
rlabel metal2 15904 24696 15904 24696 0 _204_
rlabel metal2 14616 22456 14616 22456 0 _205_
rlabel metal2 16520 18032 16520 18032 0 _206_
rlabel metal2 16968 19600 16968 19600 0 _207_
rlabel metal3 21560 37912 21560 37912 0 _208_
rlabel metal3 18256 23912 18256 23912 0 _209_
rlabel metal2 14952 22120 14952 22120 0 _210_
rlabel metal2 9576 25816 9576 25816 0 _211_
rlabel metal4 17192 21840 17192 21840 0 _212_
rlabel metal2 15400 21840 15400 21840 0 _213_
rlabel metal2 16744 23072 16744 23072 0 _214_
rlabel metal2 18256 22120 18256 22120 0 _215_
rlabel metal2 9016 24304 9016 24304 0 _216_
rlabel metal3 20552 22344 20552 22344 0 _217_
rlabel metal2 24304 28504 24304 28504 0 _218_
rlabel metal2 27272 25088 27272 25088 0 _219_
rlabel metal2 24472 31360 24472 31360 0 _220_
rlabel metal2 23352 29624 23352 29624 0 _221_
rlabel metal2 24920 29008 24920 29008 0 _222_
rlabel metal2 19880 16912 19880 16912 0 _223_
rlabel metal2 24360 20496 24360 20496 0 _224_
rlabel metal2 24808 28728 24808 28728 0 _225_
rlabel metal2 19992 18536 19992 18536 0 _226_
rlabel metal2 18872 27776 18872 27776 0 _227_
rlabel metal2 14728 35756 14728 35756 0 _228_
rlabel metal2 18648 28168 18648 28168 0 _229_
rlabel metal2 18424 27608 18424 27608 0 _230_
rlabel metal3 20328 28728 20328 28728 0 _231_
rlabel metal2 21728 26488 21728 26488 0 _232_
rlabel metal3 25172 26376 25172 26376 0 _233_
rlabel metal3 23184 28616 23184 28616 0 _234_
rlabel metal2 17360 14392 17360 14392 0 _235_
rlabel metal2 17528 15456 17528 15456 0 _236_
rlabel metal3 20104 16856 20104 16856 0 _237_
rlabel metal2 17416 15344 17416 15344 0 _238_
rlabel metal3 17416 15288 17416 15288 0 _239_
rlabel metal2 18760 17696 18760 17696 0 _240_
rlabel metal3 17752 19936 17752 19936 0 _241_
rlabel metal3 5656 20776 5656 20776 0 _242_
rlabel metal2 16408 19040 16408 19040 0 _243_
rlabel metal2 13384 26768 13384 26768 0 _244_
rlabel metal2 9016 19936 9016 19936 0 _245_
rlabel metal2 8960 20216 8960 20216 0 _246_
rlabel metal2 3192 16408 3192 16408 0 _247_
rlabel metal2 20552 16240 20552 16240 0 _248_
rlabel metal3 8736 15960 8736 15960 0 _249_
rlabel metal2 6104 15568 6104 15568 0 _250_
rlabel metal2 7672 20496 7672 20496 0 _251_
rlabel metal2 23016 28840 23016 28840 0 _252_
rlabel metal2 23240 33040 23240 33040 0 _253_
rlabel metal2 27664 23128 27664 23128 0 _254_
rlabel metal2 27440 23128 27440 23128 0 _255_
rlabel metal2 26488 23184 26488 23184 0 _256_
rlabel metal4 22008 29344 22008 29344 0 _257_
rlabel metal3 19880 16744 19880 16744 0 _258_
rlabel metal2 19768 15288 19768 15288 0 _259_
rlabel metal2 20440 16520 20440 16520 0 _260_
rlabel metal2 20552 17640 20552 17640 0 _261_
rlabel metal2 19656 18536 19656 18536 0 _262_
rlabel metal2 21224 17864 21224 17864 0 _263_
rlabel metal2 11704 20328 11704 20328 0 _264_
rlabel metal3 4592 14728 4592 14728 0 _265_
rlabel metal3 17024 20104 17024 20104 0 _266_
rlabel metal3 15008 11480 15008 11480 0 _267_
rlabel metal2 26320 22904 26320 22904 0 _268_
rlabel metal2 10304 17080 10304 17080 0 _269_
rlabel metal3 6216 23912 6216 23912 0 _270_
rlabel metal2 27720 22176 27720 22176 0 _271_
rlabel metal2 21672 16688 21672 16688 0 _272_
rlabel metal3 19376 17752 19376 17752 0 _273_
rlabel metal2 25816 20888 25816 20888 0 _274_
rlabel metal2 19376 21000 19376 21000 0 _275_
rlabel metal2 18704 23800 18704 23800 0 _276_
rlabel metal2 26488 22568 26488 22568 0 _277_
rlabel metal2 26936 29792 26936 29792 0 _278_
rlabel metal2 27384 21112 27384 21112 0 _279_
rlabel metal2 26712 22288 26712 22288 0 _280_
rlabel metal2 25760 23352 25760 23352 0 _281_
rlabel metal2 28280 22008 28280 22008 0 _282_
rlabel metal3 28560 22904 28560 22904 0 _283_
rlabel metal2 24136 23744 24136 23744 0 _284_
rlabel metal3 26264 20776 26264 20776 0 _285_
rlabel metal2 3864 16352 3864 16352 0 _286_
rlabel metal2 3864 17528 3864 17528 0 _287_
rlabel metal2 9464 18088 9464 18088 0 _288_
rlabel metal2 24472 20384 24472 20384 0 _289_
rlabel metal2 21336 31192 21336 31192 0 _290_
rlabel metal2 30408 24976 30408 24976 0 _291_
rlabel metal2 23576 19320 23576 19320 0 _292_
rlabel metal2 24808 20216 24808 20216 0 _293_
rlabel metal2 27496 21280 27496 21280 0 _294_
rlabel metal2 25816 27048 25816 27048 0 _295_
rlabel metal3 11592 13160 11592 13160 0 _296_
rlabel metal2 17528 25032 17528 25032 0 _297_
rlabel metal2 19544 26208 19544 26208 0 _298_
rlabel metal2 27608 26432 27608 26432 0 _299_
rlabel metal2 11032 23968 11032 23968 0 _300_
rlabel metal2 23800 25592 23800 25592 0 _301_
rlabel metal2 22456 16576 22456 16576 0 _302_
rlabel metal2 30296 21112 30296 21112 0 _303_
rlabel metal2 26208 27496 26208 27496 0 _304_
rlabel metal2 25368 25032 25368 25032 0 _305_
rlabel metal2 21504 20440 21504 20440 0 _306_
rlabel metal3 5600 22456 5600 22456 0 _307_
rlabel metal2 21448 24752 21448 24752 0 _308_
rlabel metal2 27048 25760 27048 25760 0 _309_
rlabel metal3 13216 11368 13216 11368 0 _310_
rlabel metal2 27272 24136 27272 24136 0 _311_
rlabel metal3 11648 29288 11648 29288 0 _312_
rlabel metal2 21896 29400 21896 29400 0 _313_
rlabel metal2 21336 30744 21336 30744 0 _314_
rlabel metal2 15960 28224 15960 28224 0 _315_
rlabel metal2 7448 24192 7448 24192 0 _316_
rlabel metal2 2296 17808 2296 17808 0 _317_
rlabel metal2 7672 24192 7672 24192 0 _318_
rlabel metal3 6384 23128 6384 23128 0 _319_
rlabel metal2 10024 22456 10024 22456 0 _320_
rlabel metal2 8344 23968 8344 23968 0 _321_
rlabel metal2 12264 23128 12264 23128 0 _322_
rlabel metal2 11760 21336 11760 21336 0 _323_
rlabel metal2 11816 24472 11816 24472 0 _324_
rlabel metal2 26936 24080 26936 24080 0 _325_
rlabel metal2 25032 20664 25032 20664 0 _326_
rlabel metal3 22568 19320 22568 19320 0 _327_
rlabel metal2 23856 18648 23856 18648 0 _328_
rlabel metal2 24192 30408 24192 30408 0 _329_
rlabel metal2 25256 21112 25256 21112 0 _330_
rlabel metal2 25704 19712 25704 19712 0 _331_
rlabel metal2 2856 20664 2856 20664 0 _332_
rlabel metal2 2072 17360 2072 17360 0 _333_
rlabel metal3 10416 19992 10416 19992 0 _334_
rlabel metal2 17640 22176 17640 22176 0 _335_
rlabel metal2 14840 19992 14840 19992 0 _336_
rlabel metal2 15736 19824 15736 19824 0 _337_
rlabel metal2 19880 33600 19880 33600 0 _338_
rlabel metal2 5992 36512 5992 36512 0 _339_
rlabel metal2 9576 36008 9576 36008 0 _340_
rlabel metal2 6776 38248 6776 38248 0 _341_
rlabel metal3 3052 37128 3052 37128 0 _342_
rlabel metal2 8232 36848 8232 36848 0 _343_
rlabel metal2 8400 34888 8400 34888 0 _344_
rlabel metal2 10080 32536 10080 32536 0 _345_
rlabel metal2 12040 32760 12040 32760 0 _346_
rlabel metal2 7000 31864 7000 31864 0 _347_
rlabel metal2 2296 33768 2296 33768 0 _348_
rlabel metal2 2968 34608 2968 34608 0 _349_
rlabel metal2 3192 26572 3192 26572 0 _350_
rlabel metal2 6776 33040 6776 33040 0 _351_
rlabel metal2 7840 32648 7840 32648 0 _352_
rlabel metal3 16296 34104 16296 34104 0 _353_
rlabel metal2 16800 33320 16800 33320 0 _354_
rlabel metal3 22960 23240 22960 23240 0 _355_
rlabel metal3 22680 23128 22680 23128 0 _356_
rlabel metal2 3416 29344 3416 29344 0 _357_
rlabel metal2 2968 29736 2968 29736 0 _358_
rlabel metal3 2884 29400 2884 29400 0 _359_
rlabel metal2 6664 31808 6664 31808 0 _360_
rlabel metal2 16072 32592 16072 32592 0 _361_
rlabel metal3 17360 14616 17360 14616 0 _362_
rlabel metal2 3192 37184 3192 37184 0 _363_
rlabel metal2 13720 36120 13720 36120 0 _364_
rlabel metal2 15176 36624 15176 36624 0 _365_
rlabel metal2 12824 35280 12824 35280 0 _366_
rlabel metal2 10808 34944 10808 34944 0 _367_
rlabel metal2 4312 36624 4312 36624 0 _368_
rlabel metal2 10248 34048 10248 34048 0 _369_
rlabel metal2 15512 28168 15512 28168 0 _370_
rlabel metal2 15456 23912 15456 23912 0 _371_
rlabel metal3 19320 17528 19320 17528 0 _372_
rlabel metal2 4928 33432 4928 33432 0 _373_
rlabel metal2 10808 32872 10808 32872 0 _374_
rlabel metal3 18536 17416 18536 17416 0 _375_
rlabel metal2 12264 35560 12264 35560 0 _376_
rlabel metal2 17416 35616 17416 35616 0 _377_
rlabel metal2 21112 25088 21112 25088 0 _378_
rlabel metal2 20888 23968 20888 23968 0 _379_
rlabel metal2 19656 17752 19656 17752 0 _380_
rlabel metal2 6552 27496 6552 27496 0 _381_
rlabel metal2 6552 30912 6552 30912 0 _382_
rlabel metal2 3640 29064 3640 29064 0 _383_
rlabel metal2 12936 26880 12936 26880 0 _384_
rlabel metal2 19544 15680 19544 15680 0 _385_
rlabel metal3 16576 38248 16576 38248 0 bus_out[0]
rlabel metal2 19544 37128 19544 37128 0 bus_out[1]
rlabel metal3 24136 38248 24136 38248 0 bus_out[2]
rlabel metal2 26040 39354 26040 39354 0 bus_out[3]
rlabel metal2 29400 41146 29400 41146 0 bus_out[4]
rlabel metal2 32760 39746 32760 39746 0 bus_out[5]
rlabel metal2 36120 39746 36120 39746 0 bus_out[6]
rlabel metal2 39480 39298 39480 39298 0 bus_out[7]
rlabel metal2 5880 39942 5880 39942 0 cs_port[0]
rlabel metal2 9072 38920 9072 38920 0 cs_port[1]
rlabel metal3 13440 38024 13440 38024 0 cs_port[2]
rlabel metal2 1848 35728 1848 35728 0 last_addr[0]
rlabel metal2 2240 34664 2240 34664 0 last_addr[1]
rlabel metal2 1736 36176 1736 36176 0 last_addr[2]
rlabel metal3 1960 35168 1960 35168 0 last_addr[3]
rlabel metal3 952 35896 952 35896 0 last_addr[4]
rlabel metal3 1246 36568 1246 36568 0 last_addr[5]
rlabel metal2 2408 37688 2408 37688 0 last_addr[6]
rlabel metal3 2058 38360 2058 38360 0 last_addr[7]
rlabel metal3 20328 31192 20328 31192 0 net1
rlabel metal2 2744 37576 2744 37576 0 net10
rlabel metal2 2296 37520 2296 37520 0 net11
rlabel metal2 2016 18648 2016 18648 0 net12
rlabel metal2 2576 24248 2576 24248 0 net13
rlabel metal3 4368 18984 4368 18984 0 net14
rlabel metal3 1736 29512 1736 29512 0 net15
rlabel metal2 2072 30240 2072 30240 0 net16
rlabel metal2 3696 24248 3696 24248 0 net17
rlabel metal2 3136 22344 3136 22344 0 net18
rlabel metal2 3192 18592 3192 18592 0 net19
rlabel metal2 20552 30800 20552 30800 0 net2
rlabel metal2 2744 20440 2744 20440 0 net20
rlabel metal2 2128 20104 2128 20104 0 net21
rlabel metal2 2072 20440 2072 20440 0 net22
rlabel metal3 3136 22120 3136 22120 0 net23
rlabel metal2 1848 19264 1848 19264 0 net24
rlabel metal2 2128 24808 2128 24808 0 net25
rlabel metal2 3248 21784 3248 21784 0 net26
rlabel metal3 3192 23352 3192 23352 0 net27
rlabel metal3 1848 20776 1848 20776 0 net28
rlabel metal3 5180 13720 5180 13720 0 net29
rlabel metal2 19992 34272 19992 34272 0 net3
rlabel metal2 3864 14112 3864 14112 0 net30
rlabel metal2 2800 15288 2800 15288 0 net31
rlabel metal2 2744 15848 2744 15848 0 net32
rlabel metal2 2128 15512 2128 15512 0 net33
rlabel metal2 2128 15960 2128 15960 0 net34
rlabel metal2 2688 18424 2688 18424 0 net35
rlabel metal2 3752 7364 3752 7364 0 net36
rlabel metal2 4088 7924 4088 7924 0 net37
rlabel metal3 3472 7672 3472 7672 0 net38
rlabel metal3 2912 8120 2912 8120 0 net39
rlabel metal3 2576 34104 2576 34104 0 net4
rlabel metal3 4200 9240 4200 9240 0 net40
rlabel metal2 1792 9688 1792 9688 0 net41
rlabel metal2 3192 15512 3192 15512 0 net42
rlabel metal2 2128 12376 2128 12376 0 net43
rlabel metal2 28728 30688 28728 30688 0 net44
rlabel metal3 21336 37800 21336 37800 0 net45
rlabel metal2 23688 37744 23688 37744 0 net46
rlabel metal2 25928 37296 25928 37296 0 net47
rlabel metal2 28840 26684 28840 26684 0 net48
rlabel metal3 30688 26376 30688 26376 0 net49
rlabel metal2 2632 34384 2632 34384 0 net5
rlabel metal3 31304 24024 31304 24024 0 net50
rlabel metal3 33600 19880 33600 19880 0 net51
rlabel metal2 2296 32816 2296 32816 0 net6
rlabel metal2 2856 34048 2856 34048 0 net7
rlabel metal2 2968 36680 2968 36680 0 net8
rlabel metal2 3640 37520 3640 37520 0 net9
rlabel metal2 1736 18088 1736 18088 0 ram_end[0]
rlabel metal3 1246 26712 1246 26712 0 ram_end[10]
rlabel metal2 3304 27888 3304 27888 0 ram_end[11]
rlabel metal2 1848 28952 1848 28952 0 ram_end[12]
rlabel metal2 1736 30464 1736 30464 0 ram_end[13]
rlabel metal3 1848 30968 1848 30968 0 ram_end[14]
rlabel metal2 2520 31584 2520 31584 0 ram_end[15]
rlabel metal2 1736 18872 1736 18872 0 ram_end[1]
rlabel metal2 2408 19768 2408 19768 0 ram_end[2]
rlabel metal2 1736 20272 1736 20272 0 ram_end[3]
rlabel metal2 1736 20720 1736 20720 0 ram_end[4]
rlabel metal2 1848 22624 1848 22624 0 ram_end[5]
rlabel metal3 1358 23128 1358 23128 0 ram_end[6]
rlabel metal2 1736 24360 1736 24360 0 ram_end[7]
rlabel metal2 1848 25256 1848 25256 0 ram_end[8]
rlabel metal2 2408 25312 2408 25312 0 ram_end[9]
rlabel metal3 1246 3416 1246 3416 0 ram_start[0]
rlabel metal2 1736 12544 1736 12544 0 ram_start[10]
rlabel metal2 1736 13496 1736 13496 0 ram_start[11]
rlabel metal2 3416 14224 3416 14224 0 ram_start[12]
rlabel metal3 1582 15064 1582 15064 0 ram_start[13]
rlabel metal2 1680 15400 1680 15400 0 ram_start[14]
rlabel metal2 1736 16464 1736 16464 0 ram_start[15]
rlabel metal2 1736 4648 1736 4648 0 ram_start[1]
rlabel metal2 1736 5544 1736 5544 0 ram_start[2]
rlabel metal2 1736 6328 1736 6328 0 ram_start[3]
rlabel metal2 1736 7224 1736 7224 0 ram_start[4]
rlabel metal2 1736 8008 1736 8008 0 ram_start[5]
rlabel metal2 1736 8904 1736 8904 0 ram_start[6]
rlabel metal2 1960 9744 1960 9744 0 ram_start[7]
rlabel metal2 1736 10920 1736 10920 0 ram_start[8]
rlabel metal2 1736 11816 1736 11816 0 ram_start[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
