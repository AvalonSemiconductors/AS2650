* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

.subckt wrapped_as2650 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vdd vss wb_clk_i wb_rst_i
XFILLER_67_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7406__A1 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7963_ _0082_ clknet_leaf_45_wb_clk_i as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6914_ _2464_ _2567_ _2575_ _2475_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6425__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7894_ _0013_ clknet_leaf_58_wb_clk_i as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7709__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ as2650.stack\[3\]\[4\] _2507_ _2508_ as2650.stack\[0\]\[4\] _2509_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6776_ _2434_ _2439_ _2440_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3988_ _3523_ _3495_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5727_ _1525_ _1527_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4943__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6160__I _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ _1244_ _1234_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4609_ _0452_ _0460_ _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _1384_ _1393_ _1394_ _1396_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8037__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7328_ _2970_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7645__A1 _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7259_ _2828_ _0491_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5656__B1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3959__I _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6335__I _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4631__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4934__A2 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6136__A1 _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6687__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7636__A1 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6439__A2 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6611__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4960_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7785__B _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4891_ _0435_ _0718_ _0735_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6630_ _2241_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6561_ _0312_ _1796_ _2228_ _3511_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5512_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6127__A1 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6492_ _3611_ _3576_ _1915_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5443_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7875__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4689__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5374_ _0967_ as2650.r123_2\[1\]\[3\] _1187_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7113_ _2579_ _2768_ _2769_ _2581_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4325_ _3859_ _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8093_ _0212_ clknet_leaf_31_wb_clk_i as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _2001_ _2698_ _2700_ _2702_ _2378_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_59_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ as2650.holding_reg\[0\] _3784_ _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__I0 as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6850__A2 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4187_ _3722_ _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6602__A2 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7946_ _0065_ clknet_leaf_49_wb_clk_i as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7877_ _1414_ _2214_ _3455_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6828_ _2488_ _2438_ _2491_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4831__C _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6759_ _2362_ _2423_ _2375_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7866__A1 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6669__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7714__I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6758__C _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4852__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A1 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5409__I _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6949__B _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7857__A1 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4110_ _3480_ as2650.r123_2\[0\]\[7\] _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ _0859_ _0927_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4041_ _3489_ _3567_ _3576_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4843__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7800_ _0265_ _0353_ _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6596__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5992_ _1731_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7731_ _3336_ _3061_ _3347_ _3352_ _1986_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4943_ _0369_ _0774_ _0792_ _3746_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4071__A2 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7662_ _3031_ _3281_ _3286_ _2099_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4874_ _0705_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6613_ _1540_ _1649_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7593_ net34 net51 net32 _3149_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_127_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5020__A1 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6544_ _2212_ _1196_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _1920_ _2153_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5426_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6520__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5357_ _1177_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5054__I _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _3842_ _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8076_ _0195_ clknet_leaf_28_wb_clk_i as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ _0790_ _0882_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5087__A1 _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7027_ _2661_ _2675_ _2686_ _2293_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6823__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4239_ _3625_ _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7929_ _0048_ clknet_leaf_50_wb_clk_i as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4062__A2 _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6339__A1 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5937__I1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5011__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4445__S0 _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4133__I _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7872__C _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7839__A1 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5314__A2 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5078__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4509__S _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4825__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__I0 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4308__I _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6523__I _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5139__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5002__A1 _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6750__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ as2650.holding_reg\[4\] _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5553__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7354__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _1318_ _1241_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5305__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5211_ _1032_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7892__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6191_ _1361_ _1232_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _0494_ _0892_ _0893_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5069__A1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5069__B2 _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _3833_ _0830_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4816__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4024_ _3557_ _3558_ _3559_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_37_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6569__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7230__A2 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5975_ _1721_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7529__I _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4044__A2 _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7781__A3 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7714_ net40 _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4926_ _3643_ _3691_ _3663_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_100_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7645_ _2721_ _2657_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4857_ _0700_ _0706_ _0547_ _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5049__I _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7576_ _1848_ _1023_ _2826_ _3203_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4788_ _0599_ _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6527_ _2180_ _0561_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6458_ _2072_ _2136_ _2139_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5409_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6389_ _0940_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8128_ _0247_ clknet_leaf_59_wb_clk_i as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4837__B _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8059_ _0178_ clknet_leaf_18_wb_clk_i as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5512__I _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4807__A1 _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3967__I _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7439__I _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5232__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4035__A2 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6343__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6980__A1 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4291__C _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6980__B2 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5535__A2 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7288__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6799__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__I _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4649__I1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5066__A4 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4274__A2 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4026__A2 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _3585_ _3626_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6971__A1 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4711_ _3649_ as2650.r123_2\[1\]\[6\] _3493_ _3863_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _1372_ _1496_ _1497_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7430_ _1990_ _2832_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4642_ net9 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5526__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7361_ _2994_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4573_ _0413_ _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _1267_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7279__A2 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7292_ _1485_ _2876_ _2052_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6243_ _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6174_ _1872_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5125_ _0838_ _0962_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5332__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5056_ _3881_ _0892_ _0893_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4265__A2 _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4007_ _3542_ _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7754__A3 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6962__A1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5765__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5958_ _1625_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _0755_ _0757_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5889_ _1653_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7628_ _2253_ _3253_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5517__A2 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7559_ _1593_ _3001_ _3187_ _2529_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6493__A3 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6338__I _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7878__B _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4256__A2 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6705__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_14_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8093__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4334__I3 as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5692__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4495__B3 _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7930__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6930_ _2588_ _2590_ _2591_ _2555_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5995__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7300__C _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6861_ _1688_ _2523_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7197__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5812_ as2650.stack\[2\]\[7\] _1584_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6792_ _2408_ _2415_ _2455_ _2456_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6944__A1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ _1542_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6711__I _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5674_ as2650.psu\[7\] _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7413_ _1415_ _3040_ _3043_ _3045_ _2069_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4625_ _0424_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4231__I as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7344_ _2978_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4556_ _0316_ _0380_ _0409_ _3909_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_117_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7275_ _2825_ _0553_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4487_ _0339_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6226_ _1911_ _1912_ _1916_ _1923_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_103_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5683__A1 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ _1299_ _1855_ _1857_ _1804_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_112_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _3713_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6088_ _3848_ _1796_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5039_ _0859_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5986__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7188__A1 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6935__A1 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7360__A1 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput20 net20 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput31 net31 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7953__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5901__S _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3988__A1 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7179__A1 _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4316__I _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6926__A1 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4401__A2 _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7351__A1 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6154__A2 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7351__B2 _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4051__I as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4165__A1 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4410_ _3938_ _0263_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5390_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4341_ _3557_ _3626_ _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7060_ _1614_ _2244_ _2718_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4272_ _3557_ _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6011_ _1744_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7406__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5610__I _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7962_ _0081_ clknet_leaf_43_wb_clk_i as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6913_ _2306_ _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7893_ _0012_ clknet_leaf_58_wb_clk_i as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6844_ _2287_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7590__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3987_ _3522_ _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6775_ _1420_ _1969_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5726_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5657_ _3767_ _1453_ _1456_ _1388_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_108_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4608_ _3937_ _0442_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5588_ _1395_ _3664_ _0656_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4539_ as2650.r123\[0\]\[4\] _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7327_ _1685_ as2650.stack\[7\]\[4\] _2969_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7645__A2 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7258_ _2899_ _2909_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5656__A1 _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5006__B _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5656__B2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6209_ _1236_ _1905_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7189_ _3556_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4136__I _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6908__A1 as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4395__A1 _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6136__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4147__A1 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__A1 as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4698__A2 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4739__C _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8131__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7785__C _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4890_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7021__B1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4386__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7999__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _1197_ _1222_ _2082_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5511_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6491_ _0831_ _1913_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5442_ _3672_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5373_ _1181_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_114_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__I _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7112_ _2579_ _2754_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4324_ as2650.r0\[2\] _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8092_ _0211_ clknet_leaf_25_wb_clk_i as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7043_ _1613_ _2701_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4255_ _3774_ _3790_ _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4310__A1 _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4186_ _3621_ _3721_ _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7041__B _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4861__A2 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7945_ _0064_ clknet_leaf_37_wb_clk_i as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7876_ _3472_ _3473_ _2688_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7012__B1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6827_ _2490_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5169__A3 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6171__I _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8004__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6758_ _2364_ _2415_ _2421_ _2422_ _2373_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_108_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5709_ _1510_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6118__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6689_ _1572_ _2298_ _2355_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7866__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5515__I _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7618__A2 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5629__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6054__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A1 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4604__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__A1 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7177__I _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7306__A1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6949__C _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7857__A2 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5425__I _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5096__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6293__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4040_ _3573_ _3575_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4843__A2 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6256__I _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5991_ _1610_ as2650.stack\[5\]\[8\] _1726_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6596__A2 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7730_ _1625_ _3002_ _3351_ _2459_ _3013_ _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8027__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4942_ _0787_ _0791_ _3909_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7661_ _3283_ _3285_ _3047_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4873_ _3775_ _0699_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_60_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4504__I _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ _2271_ _2276_ _2279_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7592_ net35 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5020__A2 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6543_ net4 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6474_ _2133_ _2152_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5859__A1 as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5425_ _3593_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4531__A1 _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5356_ as2650.r123\[3\]\[4\] _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ _3836_ _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8075_ _0194_ clknet_leaf_28_wb_clk_i as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5287_ _1114_ _0841_ _0881_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6594__C _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7026_ _2599_ _2660_ _2685_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4238_ _3766_ _3769_ _3773_ _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ _3701_ _3704_ _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6587__A2 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7784__A1 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7928_ _0047_ clknet_leaf_4_wb_clk_i as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4062__A3 _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7859_ _3454_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4445__S1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7839__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4522__A1 _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7460__I _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_39_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6275__A1 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4825__A2 _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7775__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7527__A1 _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6735__C1 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5002__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6889__I0 as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__I as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _1040_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_124_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6190_ _1887_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4994__I _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5141_ _0976_ _0977_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6266__A1 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4116__I1 as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _0830_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7303__C _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4023_ as2650.ins_reg\[7\] _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4943__B _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6569__A2 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6714__I _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _1573_ as2650.stack\[5\]\[1\] _1720_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4044__A3 _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7713_ _3018_ _3334_ _3335_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ _0699_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4234__I _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7644_ _3246_ _3247_ _2939_ _3269_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4856_ _3578_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7575_ _3198_ _3201_ _3202_ _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4787_ _0601_ _0602_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6526_ _2199_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4752__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__I _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6457_ _0973_ _2137_ _2138_ _2071_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5408_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6388_ _3526_ _1886_ _2072_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8127_ _0246_ clknet_leaf_44_wb_clk_i as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _1013_ _0992_ _1164_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6257__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8058_ _0177_ clknet_leaf_15_wb_clk_i as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7009_ _2667_ _2668_ _1255_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__B _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7757__A1 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5232__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7509__A1 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6980__A2 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4991__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3983__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__A3 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6496__A1 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7404__B _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6248__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6799__A2 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4649__I2 as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4319__I _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7748__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5759__B1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4026__A3 _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__A1 _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _0396_ as2650.r123\[1\]\[6\] _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A1 as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5690_ as2650.psl\[7\] _1372_ _1431_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4989__I _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _0440_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5526__A3 _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4734__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5782__I0 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4572_ _0424_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7360_ _1352_ _2304_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6311_ _2004_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7291_ _2866_ _1055_ _2937_ _2938_ _2939_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_143_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6487__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6242_ _3675_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6709__I _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6173_ _1358_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5613__I _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5124_ _0407_ _0840_ _0959_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_111_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4229__I _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5055_ _0894_ _0846_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4006_ _3541_ _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7739__A1 _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6411__A1 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5957_ _1706_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6962__A2 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _0661_ _3839_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5888_ _1659_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7627_ _3249_ _3251_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4839_ _0687_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7558_ _1689_ _3024_ _3184_ _3186_ _2338_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ net41 _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7489_ _2418_ _3119_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6478__A1 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5523__I _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5453__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4964__A1 _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4716__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_wb_clk_i clknet_opt_1_1_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6469__A1 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7666__B1 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7130__A2 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A3 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5692__A2 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6973__B _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4049__I _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5819__I1 as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5589__B _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6860_ as2650.pc\[4\] _2465_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_90_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ _1603_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6791_ _1854_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4955__A1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5742_ as2650.stack_ptr\[1\] _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5673_ _1479_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6213__B _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__I _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7412_ _3041_ _3042_ _3044_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _0475_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7343_ _1707_ as2650.stack\[7\]\[12\] _2969_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4555_ _3637_ _0405_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7274_ _2828_ _0559_ _2886_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7121__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4486_ _0303_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6225_ _1522_ _1917_ _1918_ _1922_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_132_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6880__A1 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _1856_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5107_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ _1793_ _1795_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_57_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6632__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _0828_ _0874_ _0878_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6174__I _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5199__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6989_ as2650.pc\[8\] _0668_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7360__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5371__A1 as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4174__A2 _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7733__I _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput21 net21 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7112__A2 _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput43 net43 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5123__A1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6623__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7179__A2 _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6926__A2 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8060__CLK clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4937__A1 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5428__I _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6687__C _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4340_ _3668_ _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5114__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4271_ _3754_ _3805_ _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6010_ _1679_ as2650.stack\[0\]\[1\] _1743_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7961_ _0080_ clknet_leaf_39_wb_clk_i as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7311__C _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6912_ _2569_ _2573_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7892_ _0011_ clknet_leaf_61_wb_clk_i as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6843_ _2283_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6774_ _2384_ _2437_ _2438_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5976__I0 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3986_ _3521_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ _1386_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5656_ _3644_ _1420_ _0580_ _1457_ _1462_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4607_ _0453_ _0455_ _0459_ _3939_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4156__A2 _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5587_ _3597_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7326_ _2960_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4538_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7257_ _2020_ _2885_ _2908_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4469_ _3723_ _0277_ _0323_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__A2 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6853__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6208_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7188_ _1370_ _2842_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6139_ as2650.addr_buff\[4\] _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5022__B _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6081__A2 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8083__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A1 _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4631__A3 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4919__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4395__A2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7333__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3991__I _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6079__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7412__B _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7021__B2 as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7572__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4386__A2 _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5583__A1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5510_ _1308_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6490_ _1793_ _1890_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7324__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5335__A1 _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5441_ _1249_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7875__A3 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5372_ _0933_ _1182_ _1186_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7111_ _2763_ _2767_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7088__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4323_ as2650.r123\[1\]\[2\] as2650.r123_2\[1\]\[2\] _3647_ _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8091_ _0210_ clknet_leaf_39_wb_clk_i as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6835__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7042_ _1607_ _1693_ _2623_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4254_ _3772_ _3777_ _3778_ _3781_ _3789_ _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6717__I as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4185_ _3592_ _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6063__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7260__A1 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7944_ _0063_ clknet_leaf_38_wb_clk_i as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7875_ _2013_ _3456_ _3459_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7012__A1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7012__B2 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ net9 _2489_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5949__I0 as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7943__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6757_ _2267_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5068__I _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3969_ as2650.ins_reg\[6\] _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5708_ _1414_ _1512_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _1898_ _2336_ _2354_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6118__A3 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5639_ _1267_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7309_ _2914_ _0780_ _2859_ _1401_ _2956_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_137_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6826__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5629__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output42_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7251__A1 _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A1 as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5687__B _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5907__S _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5706__I _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6965__C _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6817__A1 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7490__A1 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5441__I _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4057__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7242__A1 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _1604_ _1718_ _1730_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4056__A1 _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7966__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4941_ _3719_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7368__I _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6272__I _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7660_ _1836_ _3252_ _3284_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4872_ as2650.holding_reg\[6\] _3775_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6611_ as2650.stack\[5\]\[0\] _2277_ _2278_ as2650.stack\[7\]\[0\] _2279_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5556__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7591_ _3020_ _3216_ _3218_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5020__A3 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6542_ _2185_ _2210_ _2211_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_119_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6473_ _3587_ _2145_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5616__I _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5859__A2 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4516__C1 _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__C _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5355_ _1176_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4531__A2 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6808__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4306_ _3539_ _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8074_ _0193_ clknet_leaf_26_wb_clk_i as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5286_ _0841_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7481__A1 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7025_ _2684_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4237_ _3753_ _3772_ _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4295__A1 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4168_ _3520_ _3703_ _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4047__A1 _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4099_ _3519_ _3634_ _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7784__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7927_ _0046_ clknet_leaf_6_wb_clk_i as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4598__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7858_ _0662_ _1529_ _3459_ _1848_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5547__A1 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6809_ _2053_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8121__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7789_ _2068_ _3388_ _3389_ _3396_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4430__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7472__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6275__A2 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7472__B2 _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5261__I _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7989__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7775__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7527__A2 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A1 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6735__B1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4340__I _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6889__I1 as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5710__A1 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _0845_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4496__B _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7463__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6266__A2 _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5071_ _0902_ _0904_ _0906_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4022_ as2650.ins_reg\[6\] _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7600__B _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4943__C _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6569__A3 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5973_ _1715_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7098__I _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__B _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7712_ net39 _3017_ _1883_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4515__I _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4924_ _0773_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7643_ _2167_ _3264_ _3268_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5529__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _0570_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7574_ _3198_ _3201_ _0314_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4201__A1 _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4786_ _0636_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6525_ _2198_ net44 _2178_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _1448_ _2077_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6387_ _1886_ _2071_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8126_ _0245_ clknet_leaf_44_wb_clk_i as2650.stack_ptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5338_ _1167_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6257__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7454__B2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8057_ _0176_ clknet_leaf_15_wb_clk_i as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5269_ _0662_ _0880_ _0881_ _1103_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7008_ _1833_ _2059_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7757__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4425__I _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4991__A2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6193__A1 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5535__A4 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8017__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7445__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6248__A2 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4259__A1 _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5920__S _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4649__I3 as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6815__I _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5759__A1 _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5759__B2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4982__A2 _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4640_ _0382_ _0381_ _0340_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7381__B1 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5526__A4 _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4571_ _0328_ _0414_ _0423_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6310_ _1997_ _1998_ _2003_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_116_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7290_ _2867_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7684__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6487__A2 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6241_ _1938_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4498__A1 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5123_ _0960_ _0885_ _0839_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _3883_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5998__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4005_ _3540_ _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__A1 as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4670__B2 _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5956_ as2650.stack\[1\]\[11\] _1705_ _1697_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ _0628_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5887_ _1579_ as2650.stack\[4\]\[2\] _1657_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7626_ _1833_ _3249_ _3251_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4838_ _3821_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6175__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7557_ _2545_ _3185_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4769_ _0593_ _0611_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6508_ _2177_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5009__C _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7488_ _2419_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7124__B1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7675__A1 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6478__A2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6439_ _2121_ _2119_ _2048_ _1554_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7427__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8109_ _0228_ clknet_leaf_19_wb_clk_i net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__A2 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4964__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3994__I _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6166__A1 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7363__B1 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7415__B _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7666__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7666__B2 _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6545__I _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _1602_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6790_ _1218_ _2450_ _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4404__A1 _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4955__A2 _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5672_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6157__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6213__C _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7411_ _0313_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4623_ _0418_ _0422_ _0421_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5904__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7342_ _2977_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _0407_ _3632_ _3850_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7657__A1 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7273_ _2830_ _0588_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4485_ as2650.holding_reg\[3\] _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6224_ _1920_ _1407_ _1888_ _1921_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7409__A1 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6880__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6155_ _1376_ _1246_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4891__A1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5106_ as2650.r123_2\[0\]\[3\] _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6086_ _3586_ _1794_ _1238_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6455__I _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6632__A2 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5037_ as2650.r123_2\[2\]\[0\] _0875_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4643__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6396__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6988_ _1609_ _2359_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5939_ as2650.pc\[7\] _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6190__I _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7219__C _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7609_ _2617_ _3235_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7648__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput11 net11 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5534__I _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput33 net33 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput44 net44 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6320__A1 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4882__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6623__A2 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7820__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4634__A1 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5709__I _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7145__B _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5444__I _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7103__A3 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _3625_ _3705_ _3804_ _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6984__B _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6862__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5380__S _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4873__A1 _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7811__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7960_ _0079_ clknet_leaf_39_wb_clk_i as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6911_ _2468_ _2470_ _2525_ _2572_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_35_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7891_ _0010_ clknet_leaf_61_wb_clk_i as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6842_ _2282_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6378__A1 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6773_ _2390_ _2394_ _2436_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3985_ _3520_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6224__B _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5724_ _1526_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7039__C _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7878__A1 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5655_ as2650.psl\[1\] _1460_ _0288_ as2650.overflow _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6925__I0 as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4606_ _3916_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5586_ _3597_ _0775_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6550__A1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7325_ _1723_ _2961_ _2968_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4537_ _0390_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4398__C _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7256_ _2857_ _2902_ _2907_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4468_ _3722_ _0310_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6207_ _1342_ _1362_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6853__A2 _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7187_ _3553_ _3584_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4399_ _3815_ _3928_ _3932_ _3773_ _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6138_ _1480_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6185__I _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7802__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _3848_ _1558_ _1341_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4616__A1 _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A1 _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7030__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4919__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7869__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7744__I _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6541__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4607__A1 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4083__A2 _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7021__A2 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5032__A1 _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5439__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5583__A2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5440_ _3527_ _3589_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6532__A1 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7895__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ as2650.r123_2\[1\]\[2\] _1183_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7110_ _2764_ _2766_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4322_ _3856_ _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8090_ _0209_ clknet_leaf_3_wb_clk_i as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7041_ _2330_ _2699_ _1255_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6835__A2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4253_ _3782_ _3786_ _3788_ _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4184_ _3637_ _3710_ _3717_ _3719_ _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_1_1_wb_clk_i clknet_opt_1_0_wb_clk_i clknet_opt_1_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5123__B _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4518__I _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6599__A1 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7943_ _0062_ clknet_leaf_38_wb_clk_i as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4074__A2 _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7874_ as2650.psu\[1\] _3471_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6825_ as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\] _3481_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5949__I1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6756_ _2418_ _2420_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6771__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3968_ _3500_ _3503_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5707_ _1340_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6687_ _2338_ _2300_ _2352_ _2353_ _2242_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5638_ _1444_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ _1355_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7079__A2 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7308_ _2216_ _2875_ _2955_ _1938_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6826__A2 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7239_ _1482_ _2876_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5885__I0 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7251__A2 _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A2 _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5014__A1 _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4163__I _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7711__B1 _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5923__S _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6817__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6818__I as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5722__I _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4338__I _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4056__A2 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4940_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ as2650.holding_reg\[7\] _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6610_ _1650_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7590_ net34 _3217_ _3125_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5556__A2 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6541_ net21 _2178_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6472_ _1320_ _1871_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4516__B1 _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5423_ _3490_ _1209_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4516__C2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5354_ as2650.r123\[3\]\[3\] _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4305_ _3836_ _3714_ _3744_ _3839_ _3840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8073_ _0192_ clknet_leaf_35_wb_clk_i as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6808__A2 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5285_ _0775_ _0886_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5632__I _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7024_ _2408_ _2660_ _2683_ _1243_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4236_ _3771_ _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5492__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ as2650.r123\[0\]\[1\] _3702_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\]
+ _3477_ _3492_ _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__7910__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4098_ _3524_ _3633_ _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4047__A2 _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7926_ _0045_ clknet_leaf_59_wb_clk_i as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7857_ _2023_ _3458_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6808_ _2306_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6744__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5547__A2 _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7788_ _3390_ _3391_ _3395_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6739_ _2282_ _2404_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7472__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4286__A2 _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6680__B1 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5235__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3997__I _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A1 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_48_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8096__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5849__I0 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7933__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7463__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5070_ _0907_ _0909_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4277__A2 _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5474__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4021_ as2650.ins_reg\[5\] _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4029__A2 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6974__A1 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5972_ _1709_ _1717_ _1719_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7711_ _1621_ _3021_ _3328_ _1991_ _3333_ _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_80_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4923_ _3659_ _0514_ _0770_ _0372_ _0772_ _3903_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_52_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7642_ _2986_ _3267_ _3116_ _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6726__A1 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4854_ _0684_ _0570_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5529__A2 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7573_ _3199_ _3172_ _3200_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4785_ _0626_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5627__I _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ _2197_ _2020_ _2180_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6455_ _2078_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6886__C _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5406_ _1205_ _1197_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6386_ _3876_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5337_ _0967_ _0945_ _1164_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8125_ _0244_ clknet_leaf_45_wb_clk_i as2650.stack_ptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7454__A2 _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5268_ _1096_ _0886_ _1100_ _1102_ _0898_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6257__A3 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8056_ _0175_ clknet_leaf_21_wb_clk_i as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5465__A1 _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7007_ _1412_ _0940_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4219_ _3754_ _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ as2650.r0\[5\] as2650.r123_2\[0\]\[0\] _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6965__A1 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7909_ _0028_ clknet_leaf_62_wb_clk_i as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6921__I _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4991__A3 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7238__B _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6193__A2 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7390__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8060__D _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4441__I _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7142__A1 _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7956__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6368__I _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7445__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5208__A1 _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5759__A2 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7381__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7381__B2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__I _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4570_ _0328_ _0414_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6240_ _1237_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7684__A2 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6487__A3 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4498__A2 _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6171_ _1342_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5122_ _3930_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8111__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5053_ _0888_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5998__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4004_ as2650.ins_reg\[4\] _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4526__I _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6947__A1 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ _1621_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4906_ _0627_ _0628_ _0630_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5886_ _1658_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7625_ _0313_ _3250_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4837_ _0533_ _0686_ _0685_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6175__A2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7372__A1 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4186__A1 _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7979__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7556_ _2074_ _3162_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4768_ _0619_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6507_ _0865_ _2181_ _2183_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7487_ _2368_ _3083_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4699_ _3937_ _0550_ _0434_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6438_ _1811_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5686__A1 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ _2051_ _1223_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8108_ _0227_ clknet_leaf_26_wb_clk_i net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8039_ _0158_ clknet_leaf_19_wb_clk_i net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4110__A1 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7240__C _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6938__A1 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4880__B _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4413__A2 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7363__A1 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6166__A2 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7666__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6874__B1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A1 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6929__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__S _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ as2650.stack_ptr\[2\] _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5671_ _1477_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6157__A2 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4081__I _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7410_ _3041_ _3042_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4168__A1 _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4622_ _0468_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5904__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7606__B _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4553_ _0406_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7341_ _1705_ as2650.stack\[7\]\[11\] _2969_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7106__A1 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4484_ _0262_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7272_ _2885_ _2921_ _2922_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6223_ _1890_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7409__A2 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _1854_ _1263_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6617__B1 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__I _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5105_ _0868_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6085_ _3601_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6093__A1 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7593__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6987_ _2298_ _2646_ _2647_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8007__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5938_ _1692_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ as2650.stack\[6\]\[10\] _1634_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7608_ _2569_ _3196_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7539_ _3032_ _3166_ _3167_ _2984_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput12 net12 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput23 net23 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6856__B1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput45 net45 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6320__A2 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6608__B1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4882__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7820__A2 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6387__A2 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4398__A1 _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5926__S _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5898__A1 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7426__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__I _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__B1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6984__C _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4873__A2 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6075__A1 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7811__A2 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6910_ as2650.pc\[5\] _0577_ _2571_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7890_ _0009_ clknet_leaf_61_wb_clk_i as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6841_ _2112_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7575__A1 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6378__A2 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6291__I _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6772_ _2390_ _2394_ _2436_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3984_ as2650.ins_reg\[0\] _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6224__C _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5723_ _1507_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5654_ _1219_ _0782_ _0495_ _3650_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7878__A2 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6925__I1 as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ _0456_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5635__I _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5585_ _1386_ _1390_ _1392_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6550__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7324_ as2650.stack\[7\]\[3\] _2967_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4561__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4536_ as2650.r0\[4\] _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7255_ _2858_ _0384_ _2161_ _2197_ _2906_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _0316_ _0321_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6206_ _1895_ _1899_ _1903_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6853__A3 _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4398_ _3776_ _3930_ _3931_ _3814_ _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_98_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7186_ _1453_ _1410_ _2838_ _2840_ _1939_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4864__A2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6137_ _1840_ _1832_ _1842_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _1777_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5813__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5019_ _0823_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__B1 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__A1 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A2 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5280__I _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7254__B1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4083__A3 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7000__I _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7309__A1 _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7309__B2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5455__I _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _0913_ _1182_ _1185_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4321_ _3619_ _3855_ _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6296__A1 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7040_ _1836_ _2059_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5343__I0 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4252_ _3787_ _3578_ _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4846__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4183_ _3718_ _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6599__A2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ _0061_ clknet_leaf_41_wb_clk_i as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5271__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7548__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7873_ _1416_ _3450_ _3456_ _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4534__I _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6824_ _0386_ _2435_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7012__A3 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6220__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6755_ _2419_ _2370_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3967_ _3502_ _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6771__A2 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4782__A1 _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5706_ _1253_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6686_ _1243_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5637_ _1377_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5365__I _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5568_ _3595_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7307_ _1399_ _2954_ _1409_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4519_ _0269_ _0304_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_105_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5499_ _1299_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6287__A1 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7238_ _2872_ _0266_ _2868_ _2890_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4709__I _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7169_ _2823_ _2824_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7787__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7539__A1 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7711__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7711__B2 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4525__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7778__A1 _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6825__I0 as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6834__I _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4056__A3 _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4870_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4764__A1 _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6540_ _2187_ _1101_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6471_ _1920_ _1884_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7702__A1 _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5422_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4516__B2 _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8141_ _0260_ clknet_leaf_13_wb_clk_i as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5353_ _1175_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6269__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6010__S _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4304_ _3838_ _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8072_ _0191_ clknet_leaf_26_wb_clk_i as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5284_ _0776_ _0893_ _0885_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7023_ _1218_ _2678_ _2682_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4235_ _3770_ _3595_ _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5492__A2 _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4166_ as2650.r123_2\[0\]\[1\] _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7769__A1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4097_ _3539_ _3563_ _3622_ _3632_ _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6441__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7925_ _0044_ clknet_leaf_7_wb_clk_i as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6992__A2 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4264__I _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7856_ _1274_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6807_ _2468_ _2470_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7787_ _1357_ _3394_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6744__A2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5547__A3 _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ as2650.stack\[1\]\[2\] _2286_ _1713_ as2650.stack\[0\]\[2\] _2404_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6669_ _2266_ _2300_ _2303_ _2306_ _2335_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_137_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4507__A1 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6919__I _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5180__A1 as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5823__I _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7243__C _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4439__I as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7472__A3 _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5483__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4883__B _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6432__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7885__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7485__I _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6735__A2 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A3 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4746__A1 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5934__S _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_17_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6499__A1 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6829__I _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4349__I _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4020_ _3554_ _3555_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5474__A2 _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4029__A3 _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ as2650.stack\[5\]\[0\] _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7710_ _2775_ _3330_ _3331_ _3332_ _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_64_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4084__I _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4922_ _3659_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7641_ _3266_ _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4853_ _0690_ _0703_ _3916_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6726__A2 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4812__I _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4737__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7572_ _0579_ _0587_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4784_ _0631_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _0307_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _2133_ _2135_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7151__A2 _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _0547_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8124_ _0243_ clknet_leaf_57_wb_clk_i as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5336_ _0933_ _1162_ _1166_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8055_ _0174_ clknet_leaf_21_wb_clk_i as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5267_ _1101_ _0890_ _0891_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7006_ _2380_ _2657_ _2665_ _1953_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6662__A1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5465__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4218_ _3753_ _3574_ _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5198_ _3859_ as2650.r123_2\[0\]\[3\] _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4149_ as2650.r123\[0\]\[0\] _3684_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\]
+ as2650.psl\[4\] _3531_ _3685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5217__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6414__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7908_ _0027_ clknet_leaf_62_wb_clk_i as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4976__A1 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7839_ _2022_ _2214_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5818__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5776__I0 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6193__A3 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7390__A2 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7142__A2 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__A1 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6384__I _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6405__A1 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5208__A2 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6956__A2 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8063__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6708__A2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__A1 _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7900__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__A1 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7164__B _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6487__A4 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__I _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5695__A2 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6170_ net23 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5121_ _0402_ _0844_ _0957_ _0958_ _0842_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6644__A1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5052_ _0845_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4003_ _3537_ _3538_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6294__I _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__S _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5954_ _1704_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4905_ _0406_ _0394_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5638__I _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ _1573_ as2650.stack\[4\]\[1\] _1657_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4542__I _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7624_ _1981_ _0789_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4836_ _0533_ _0685_ _0686_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7372__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7555_ _3091_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5383__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4186__A2 _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ _0524_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7853__I _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _2182_ _0883_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7486_ _2986_ _3099_ _3116_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4698_ as2650.holding_reg\[5\] _0532_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7124__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7074__B _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6437_ _2094_ _2119_ _1974_ _1945_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5373__I _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6883__A1 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6368_ _3611_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8107_ _0226_ clknet_leaf_26_wb_clk_i net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5319_ _1124_ _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6299_ _3554_ _1989_ _1992_ _3605_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6635__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__A2 _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8038_ _0157_ clknet_leaf_13_wb_clk_i net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6418__B _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4110__A2 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4717__I _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8086__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7060__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4880__C _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8071__D _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4452__I _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7923__CLK clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6166__A3 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7363__A2 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7763__I _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5126__A1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6874__B2 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7712__B _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6626__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6929__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6842__I _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7051__A1 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5458__I _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_32_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5670_ net9 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6157__A3 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4621_ _0472_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _1734_ _2962_ _2976_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4552_ _0296_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7106__A2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7271_ _2028_ _2862_ _2751_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4483_ _3518_ _0337_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6222_ _1919_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6153_ _1235_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5104_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7814__B1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6084_ as2650.cycle\[6\] _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__I _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5142__B _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _0862_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7848__I _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7042__A1 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _1694_ _2357_ _2461_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7946__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7069__B _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5937_ as2650.stack\[1\]\[6\] _1691_ _1686_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4272__I _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _1614_ _1632_ _1645_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7345__A2 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7607_ _3031_ _3221_ _3233_ _3049_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4819_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5799_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7538_ _1269_ _3071_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5108__A1 _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7469_ _2327_ _3099_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput13 net49 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6856__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5659__A2 _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput35 net35 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6927__I _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7281__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7033__A1 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4398__A2 _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5595__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8101__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__B2 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7442__B _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7272__A1 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7811__A3 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7969__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7024__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6840_ _2478_ _2467_ _2502_ _2503_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ net8 _2435_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5586__A1 _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3983_ net10 _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _1408_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5653_ _1459_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5916__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _0358_ _0440_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5584_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7323_ _2960_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4535_ _0388_ _3669_ _3694_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6838__A1 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7254_ _1840_ _2875_ _2904_ _2905_ _1938_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4466_ _0317_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6205_ _1502_ _1897_ _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5651__I _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7185_ _1379_ _2188_ _3664_ _2839_ _1941_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4397_ _3917_ _3775_ _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6136_ _1841_ _1837_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4267__I _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6067_ _1707_ as2650.stack\[3\]\[12\] _1768_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4077__A1 _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5813__A2 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5018_ _3721_ _0858_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7015__A1 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__A2 _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8124__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _2588_ _2593_ _2629_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5826__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4001__A1 _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7262__B _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4177__I _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__A1 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__A1 _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7006__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5937__S _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7309__A2 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ _3577_ _3582_ _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7493__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6296__A2 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4251_ _3505_ _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5343__I1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5471__I _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4182_ _3693_ _3609_ _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7245__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7941_ _0060_ clknet_leaf_38_wb_clk_i as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7398__I _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7872_ _1482_ _3468_ _3470_ _2132_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6823_ _2378_ _2481_ _2486_ _2006_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5559__A1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6754_ _1576_ _0285_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3966_ _3501_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5705_ _1510_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6685_ _2350_ _2351_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5646__I _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5636_ _1442_ _1411_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5731__A1 _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ _0707_ _1246_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5731__B2 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7306_ _1394_ _2953_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4518_ _3737_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_137_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _1055_ _1305_ _1154_ _0572_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7082__B _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7237_ _2886_ _2888_ _2889_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4449_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7168_ _1625_ _2357_ _2159_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7236__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7810__B _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6119_ _1820_ _1822_ _1824_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_112_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7099_ _1702_ _2733_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7787__A2 _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A1 _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6161__B _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4460__I _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7711__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7475__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4289__A1 _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7778__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6825__I1 as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5789__A1 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4461__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6738__B1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4764__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _1987_ _2149_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5421_ _1228_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__A1 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8140_ _0259_ clknet_leaf_12_wb_clk_i as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5352_ as2650.r123\[3\]\[2\] _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7614__C _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4303_ _3837_ _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8071_ _0190_ clknet_leaf_28_wb_clk_i as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7466__B2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5283_ _0780_ _0977_ _0889_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5477__B1 _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7022_ _2679_ _2680_ _2681_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4234_ _3505_ _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5492__A3 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4165_ _3532_ _3697_ _3700_ _3550_ _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6977__B1 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4096_ _3631_ _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7924_ _0043_ clknet_leaf_59_wb_clk_i as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7855_ _1425_ _3450_ _3456_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7856__I _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6806_ _2469_ _2420_ _2417_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4998_ _0799_ _0835_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7786_ _1354_ _1860_ _3392_ _3393_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5547__A4 _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3949_ as2650.cycle\[1\] _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6737_ as2650.stack\[5\]\[2\] _2402_ _2346_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4280__I _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _2322_ _2334_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5619_ _1410_ _1422_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6599_ _1438_ _1782_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7457__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7209__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6680__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4691__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8074__D _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6432__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6196__A1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A4 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4746__A2 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7696__A1 _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6499__A2 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_57_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7620__A1 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5970_ _1716_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4921_ _0653_ _0654_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4985__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6580__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7640_ net50 _3265_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4852_ _0691_ _0697_ _0702_ _0453_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7571_ _0579_ _0587_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4783_ _0632_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4737__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _2179_ _2195_ _2196_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6453_ _1555_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ _1204_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6384_ _0315_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8123_ _0242_ clknet_leaf_57_wb_clk_i as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5335_ _3868_ _1164_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8054_ _0173_ clknet_leaf_18_wb_clk_i as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ _0720_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6111__A1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7005_ _2248_ _2659_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6662__A2 _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4217_ _3752_ _3753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5197_ _3699_ _0944_ _1004_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4148_ as2650.r123_2\[0\]\[0\] _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7611__A1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6414__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4079_ _3520_ _3614_ _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7907_ _0026_ clknet_leaf_62_wb_clk_i as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7838_ _3439_ _3441_ _3442_ _2132_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7769_ _2506_ _3376_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6193__A4 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7678__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3951__A3 as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5153__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__C _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6350__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8069__D _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7850__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6653__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6405__A2 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4416__A1 _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A1 _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4719__A2 _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__S _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7669__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5144__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _0388_ _0846_ _0843_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6575__I _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6644__A2 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5051_ _0884_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7841__A1 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7841__B2 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4655__A1 _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4002_ _3482_ _3514_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4095__I _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4407__A1 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ as2650.stack\[1\]\[10\] _1703_ _1697_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5919__I _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4904_ _0631_ _0634_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5884_ _1652_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7623_ _3198_ _3201_ _3248_ _3222_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4835_ _0444_ _0530_ _0543_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7372__A3 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7554_ _3062_ _3178_ _3182_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4766_ _0525_ _0616_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6505_ _0974_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7485_ _2077_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4697_ _0542_ _0546_ _0548_ _3829_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_101_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6436_ _2118_ _2110_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6883__A2 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6367_ _3581_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8106_ _0225_ clknet_leaf_19_wb_clk_i net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5318_ _0907_ _1151_ _0829_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6298_ _1987_ _1993_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7090__B _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6635__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7832__A1 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5249_ _1081_ _1082_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8037_ _0156_ clknet_3_6_0_wb_clk_i net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_2_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6418__C _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7249__C _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6571__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6874__A2 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4885__A1 _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5513__B _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6626__A2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7823__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6344__B _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5739__I _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4620_ _3860_ _3865_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6562__A1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7898__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4551_ _3642_ _3874_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7270_ _2913_ _2920_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4482_ as2650.r123\[2\]\[2\] _3636_ _0336_ _3800_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6314__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ _1793_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _1852_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _0937_ _0940_ _3561_ _0833_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__4818__I _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6617__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7814__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ _1382_ _1782_ _1791_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7814__B2 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A1 _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _0827_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6985_ _2622_ _2636_ _2637_ _2645_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7593__A3 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4553__I _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _1597_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7069__C _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__A1 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5867_ as2650.stack\[6\]\[9\] _1634_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7606_ _3227_ _3232_ _3047_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4818_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6553__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5798_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7537_ _1846_ _0559_ _3165_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4749_ _0599_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5384__I as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5108__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6305__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7468_ net31 _3098_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4167__I0 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput14 net14 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7813__B _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput25 net25 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6419_ _1273_ _2089_ _2055_ _1320_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput36 net36 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__8053__CLK clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7399_ _2844_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6608__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7281__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4714__S1 _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7033__A2 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5044__A1 _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6792__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5595__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A2 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4858__A1 _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__I _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6075__A3 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4086__A2 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__A1 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7024__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3982_ _3517_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6770_ as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\] _3481_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5586__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5721_ _1524_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7617__C _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _1458_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6535__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4603_ as2650.holding_reg\[4\] _3625_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5583_ _0707_ _1377_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7322_ _2966_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4534_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4149__I0 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6838__A2 _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4465_ _0318_ _3873_ _0274_ _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7253_ _2839_ _0887_ _0449_ _1398_ _1940_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5932__I as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ _1309_ _1901_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7184_ _1391_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4396_ _3929_ _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6249__B _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6135_ as2650.addr_buff\[3\] _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4548__I _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6066_ _1776_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4077__A2 _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7859__I _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _0836_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6968_ net3 _3652_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5919_ _1572_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6899_ _2524_ _2534_ _2561_ _2293_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4001__A2 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6159__B _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5265__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4068__A2 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6673__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7006__A2 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6622__B _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8099__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__A1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__A3 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5953__S _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7190__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4250_ _3624_ _3784_ _3785_ _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7936__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6069__B _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4181_ _3715_ _3716_ _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7245__A2 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7940_ _0059_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7871_ _2016_ _2214_ _3469_ _3468_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5008__A1 _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6822_ _2482_ _1852_ _2484_ _2381_ _2485_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5559__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _2416_ _2417_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3965_ as2650.ins_reg\[2\] as2650.ins_reg\[3\] _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_108_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5704_ _1502_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6684_ _1204_ _2300_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5148__B _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5635_ _1373_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5566_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7305_ _1481_ _2876_ _2952_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4517_ _0370_ _0303_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5497_ _0465_ _0553_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7082__C _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7236_ _2070_ _0277_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4448_ _0302_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5495__A1 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4379_ _3913_ _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7167_ _2599_ _2791_ _2810_ _2822_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6118_ _1783_ _1825_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7236__A2 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7098_ _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7589__I _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6049_ _1723_ _1760_ _1767_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4227__B _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6747__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5837__I _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6161__C _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6770__I1 as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5572__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7475__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5486__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__I _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5238__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A2 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6986__A1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A2 _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5747__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3972__A1 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _1198_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6910__A1 as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5351_ _1174_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6578__I _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4302_ as2650.r123\[0\]\[1\] _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7466__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8070_ _0189_ clknet_leaf_35_wb_clk_i as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5282_ _1115_ _0846_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8114__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__B2 _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4233_ _3768_ _3764_ _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7021_ as2650.stack\[3\]\[8\] _2278_ _2275_ as2650.stack\[2\]\[8\] _2681_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6674__B1 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4164_ _3699_ _3492_ _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4095_ _3630_ _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7202__I _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6977__B2 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout52_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7923_ _0042_ clknet_leaf_4_wb_clk_i as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6729__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7854_ _3455_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6805_ _2416_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7785_ _3772_ _1780_ _1252_ _1226_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4997_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6736_ _2286_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3948_ _3483_ _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7154__A1 _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6667_ _2323_ _2300_ _2332_ _2333_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5618_ _1423_ _1271_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6598_ _1438_ _2245_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4510__B _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5549_ _1355_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5392__I _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5468__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7219_ _2828_ _3908_ _2871_ _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7209__A2 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6437__B _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4691__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4736__I _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5060__C _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__A2 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7393__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8090__D _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4404__C _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6900__B _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8137__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_69_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5459__A1 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6120__A2 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4646__I _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_26_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6959__A1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4920_ _0719_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4851_ _0698_ _0699_ _0701_ _0691_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7570_ _1456_ _0678_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4782_ _3698_ as2650.r123\[0\]\[5\] _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ net43 _2192_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _1556_ _2109_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5403_ _0822_ _1208_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6383_ _1373_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4370__A1 _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8122_ _0241_ clknet_leaf_57_wb_clk_i as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ _0913_ _1162_ _1165_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8053_ _0172_ clknet_leaf_18_wb_clk_i as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5265_ _1098_ _0892_ _0844_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6111__A2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7004_ _2253_ _2663_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4122__A1 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4122__B2 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4216_ _3500_ _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5196_ _0996_ _1030_ _1031_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5870__A1 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4147_ _3532_ _3680_ _3682_ _3550_ _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4078_ _3531_ _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7906_ _0025_ clknet_leaf_4_wb_clk_i as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7837_ _3484_ _3439_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7375__A1 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7768_ _3375_ _3378_ _3379_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6719_ _1549_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7127__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7699_ _2758_ _3299_ _3300_ _3301_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5689__B2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6350__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7850__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5861__A1 as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8085__D _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7777__I _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7366__A1 _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A2 _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A3 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7118__A1 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6877__B1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4104__A1 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7841__A2 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ _3530_ _3536_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4655__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4407__A2 _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _1702_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4903_ _0644_ _0647_ _0650_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5883_ _1539_ _1654_ _1656_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7357__A1 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7622_ _1115_ _0789_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4834_ _0684_ _0664_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7553_ _3051_ _3181_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ as2650.r123\[2\]\[5\] _0433_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _2180_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6032__S _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7484_ _3108_ _3113_ _3114_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4696_ _0547_ _0530_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6435_ _1968_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5871__S _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__A1 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6366_ _1217_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8105_ _0224_ clknet_leaf_26_wb_clk_i net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4894__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7371__B _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _1125_ _1144_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5670__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6297_ _3555_ _1989_ _1992_ _3606_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7090__C _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8036_ _0155_ clknet_leaf_22_wb_clk_i as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5248_ _1081_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7832__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ _1014_ _1015_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7596__A1 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7348__A1 _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6006__I _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7546__B _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6571__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4889__C _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__I as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6087__A1 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5513__C _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7823__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7036__B1 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7587__A1 _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4924__I _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5956__S _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6360__B _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5755__I as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4550_ _0385_ _0389_ _0402_ _3695_ _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7511__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4481_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6314__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ _1216_ _1907_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6151_ _1210_ _1549_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_41_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A1 _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _1783_ _1786_ _1788_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7814__A2 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5825__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7578__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6984_ _2505_ _2615_ _2644_ _2353_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7210__I _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6254__C _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6250__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5935_ _1690_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4800__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5866_ _1644_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7605_ _1449_ _3032_ _3034_ _3231_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4817_ net2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5797_ as2650.pc\[5\] _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7750__A1 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6553__A2 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7536_ _3140_ _3163_ _3141_ _3164_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4748_ _3860_ _0298_ _0394_ _3698_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7467_ net30 net52 net28 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7502__A1 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6305__A2 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ as2650.holding_reg\[5\] _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7992__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4167__I1 _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6418_ _2079_ _2101_ _2082_ _1433_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput15 net15 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7813__C _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput26 net26 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7398_ _1800_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput37 net37 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6349_ _1425_ _1967_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6069__A1 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7805__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8019_ _0138_ clknet_leaf_36_wb_clk_i as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7321__S _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6164__C _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6792__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5776__S _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7276__B _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7741__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4555__A1 _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5807__A1 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4086__A3 _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6480__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4654__I _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6232__A1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3981_ _3516_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5720_ _1521_ _1511_ _1523_ _1419_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5651_ _3882_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7732__A1 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4546__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _0445_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4546__B2 _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5582_ _3534_ _1387_ _1257_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7321_ _1681_ as2650.stack\[7\]\[2\] _2964_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _0386_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6299__B2 _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4149__I1 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7252_ as2650.psu\[3\] _2836_ _2903_ _1444_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4464_ _3727_ _3606_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_132_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6203_ _1365_ _1900_ _1335_ _0359_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7183_ as2650.psu\[0\] _2836_ _2837_ _1445_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4395_ _3864_ _3870_ _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6249__C _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6134_ _1472_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6065_ _1705_ as2650.stack\[3\]\[11\] _1768_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6471__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5274__A2 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5016_ _3731_ _0838_ _0854_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6265__B _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _2250_ _2624_ _2626_ _2627_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5918_ _1678_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6898_ _2542_ _2560_ _2532_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__I _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5849_ _1573_ as2650.stack\[6\]\[1\] _1634_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7723__A1 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8020__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7519_ _3148_ _3098_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_120_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7824__B _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5337__I0 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6954__I _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__A1 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6462__B2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6175__B _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7888__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6214__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4776__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__B2 _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7190__A2 _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__A1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4180_ _3631_ _3716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5256__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7870_ _1967_ _3458_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5008__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _1423_ _1810_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6752_ _1581_ _1471_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8043__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4767__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3964_ as2650.ins_reg\[5\] _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5703_ _1383_ _1503_ _1506_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6683_ _2339_ _2345_ _2349_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7705__A1 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4519__A1 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5634_ _1114_ _1311_ _1312_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7644__B _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5192__A1 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5565_ _0937_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5943__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7304_ as2650.psl\[7\] _1230_ _1377_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4516_ _3757_ _3758_ _3701_ _3704_ _3864_ _3870_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_117_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5496_ _3796_ _0936_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7235_ _2887_ _0321_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4447_ _0292_ _0293_ _0297_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6692__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5495__A2 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7166_ _2297_ _2821_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4378_ _3802_ _3833_ _3912_ _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6117_ _1789_ _1785_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7097_ _1619_ _2753_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5247__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6048_ as2650.stack\[3\]\[3\] _1766_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4508__B _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4294__I _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7999_ _0118_ clknet_leaf_44_wb_clk_i as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__I _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5183__A1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8088__D _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7475__A3 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6683__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5238__A2 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6986__A2 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8066__CLK clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A3 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6738__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7903__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6910__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5350_ as2650.r123\[3\]\[1\] _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7183__C _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4301_ _3835_ _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4379__I _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5281_ _0781_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ as2650.stack\[1\]\[8\] _2277_ _2272_ as2650.stack\[0\]\[8\] _2680_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ as2650.psl\[3\] _3767_ _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ _3698_ _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4094_ _3620_ _3629_ _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6977__A2 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7922_ _0041_ clknet_leaf_4_wb_clk_i as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5003__I _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7853_ _3454_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6804_ as2650.pc\[4\] _1477_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7784_ _1507_ _1208_ _2222_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4996_ _0832_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6735_ as2650.stack\[7\]\[2\] _2342_ _2400_ as2650.stack\[6\]\[2\] _1714_ as2650.stack\[4\]\[2\]
+ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3947_ _3482_ _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6666_ _2245_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6769__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5165__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5673__I _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6597_ _1538_ _2247_ _2249_ _2251_ _2264_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6901__A2 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5548_ _1235_ _1323_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5479_ _0344_ _1283_ _1285_ _1286_ _0446_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6665__A1 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7218_ _2074_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7149_ _1619_ _1702_ _2733_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4140__A2 _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8089__CLK clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6417__A1 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6437__C _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7614__B1 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__A2 _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7090__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A2 _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7549__B _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5848__I _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7268__C _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7926__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7393__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout50 net36 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7145__A2 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5156__A1 _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7284__B _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6656__A1 _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7731__C _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6408__A1 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5959__S _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4850_ _0700_ _0539_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4781_ _3711_ as2650.r123\[0\]\[6\] _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6520_ _2016_ _2181_ _2194_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5147__A1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ as2650.cycle\[3\] _1556_ _2109_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6895__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ _1210_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6382_ _1320_ _2066_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8121_ _0240_ clknet_leaf_57_wb_clk_i as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5333_ _0905_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4370__A2 _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8052_ _0171_ clknet_3_3_0_wb_clk_i as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5264_ _0667_ _0977_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7003_ _2662_ _2631_ _0938_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4215_ _3538_ _3562_ _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4122__A2 _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5195_ _0988_ _1005_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5870__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4146_ _3681_ _3531_ _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7072__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4077_ _3579_ _3612_ _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7949__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7905_ _0024_ clknet_leaf_63_wb_clk_i as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7836_ _2028_ _2036_ _3440_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4979_ _3551_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7767_ _1674_ _3375_ _1883_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6718_ _2056_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7698_ _1914_ _3299_ _3301_ _3320_ _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_137_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5138__A1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6649_ _2314_ _2056_ _2315_ _1352_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6886__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5689__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7832__B _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4361__A2 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6638__A1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5861__A2 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8104__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5129__A1 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6877__A1 as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6877__B2 as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4352__A2 _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4104__A2 _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4000_ _3534_ _3535_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7054__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6872__I _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6801__A1 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ as2650.pc\[10\] _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4902_ _0744_ _0745_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_80_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5882_ as2650.stack\[4\]\[0\] _1655_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7621_ _2649_ _3245_ _3085_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5368__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4833_ as2650.holding_reg\[6\] _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7552_ _2525_ _3180_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4764_ _3751_ _0553_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4040__A1 _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6503_ _0974_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7483_ _3047_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4591__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4695_ _3753_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6868__A1 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6434_ _1527_ _2049_ _2110_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5540__A1 _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__A2 _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ _2047_ _1382_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5951__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8104_ _0223_ clknet_leaf_26_wb_clk_i net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5316_ _1147_ _1148_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6296_ _1991_ _1989_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8035_ _0154_ clknet_leaf_14_wb_clk_i as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6096__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _3835_ _0501_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ as2650.r123_2\[2\]\[4\] _0969_ _0970_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__A1 as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ net5 _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8127__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7348__A2 _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7819_ _3424_ _3425_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6020__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7319__S _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4031__A1 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6571__A3 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6859__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5531__A1 _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7284__A1 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4098__A1 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5101__I _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__A2 _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4270__A1 _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4940__I _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5770__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4480_ _3802_ _0266_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7511__A2 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5522__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5771__I as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _1851_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7275__A1 _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6078__A2 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5101_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _1789_ _1340_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5825__A2 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _3796_ _0830_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_10_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7578__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5589__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _2113_ _2640_ _2643_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6250__A2 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__I _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5934_ as2650.stack\[1\]\[5\] _1689_ _1686_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4261__A1 _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5865_ _1610_ as2650.stack\[6\]\[8\] _1639_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6551__B _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7604_ _3071_ _3230_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4816_ _0664_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6043__S _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5796_ _1591_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7535_ _1478_ _0516_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4747_ _3860_ _3698_ _0298_ _0393_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5761__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7466_ _3060_ _3061_ _3088_ _3097_ _2131_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4678_ as2650.holding_reg\[5\] _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7502__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6417_ _2099_ _2100_ _2091_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6777__I _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7397_ _1571_ _3024_ _3029_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4167__I2 as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput16 net16 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput27 net27 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput38 net38 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6348_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6069__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7266__A1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6279_ _1810_ _1975_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8018_ _0137_ clknet_leaf_31_wb_clk_i as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7018__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7401__I _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7569__A2 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6445__C _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__I _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A1 _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5752__A1 _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7292__B _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5504__A1 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7257__A1 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5807__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6768__B1 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6232__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3980_ _3484_ _3511_ _3515_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7186__C _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ as2650.psl\[5\] _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7732__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4601_ _0342_ _0349_ _0345_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4546__A2 _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ _1388_ _1387_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6940__B1 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7320_ _2965_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4532_ net8 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7496__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6299__A2 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7251_ _3644_ _2878_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4463_ _3729_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5346__I1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__I2 as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6202_ _3627_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7182_ _3767_ _1231_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4394_ _3921_ _3927_ _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7248__A1 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6133_ _0289_ _1832_ _1839_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6064_ _1734_ _1761_ _1775_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5015_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6471__A2 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7221__I _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4482__B2 _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6265__C _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6966_ _2216_ _2057_ _1853_ _1850_ _2032_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_81_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5917_ as2650.stack\[1\]\[0\] _1673_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6897_ _1855_ _2524_ _2531_ _2559_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_139_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5848_ _1629_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7723__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5779_ _1576_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7518_ net31 _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7449_ _1418_ _1024_ _2827_ _3080_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5337__I1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7840__B as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7239__A1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4473__A1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6922__B1 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7190__A3 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6525__I0 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7650__A1 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7402__A1 _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6820_ _2380_ _2471_ _2483_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6751_ as2650.pc\[3\] net8 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3963_ _3498_ _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ _1448_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6682_ _2346_ _2347_ _2348_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5633_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4519__A2 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6321__S _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7644__C _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5564_ _1347_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5192__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7469__A1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4515_ _3901_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7303_ _2866_ _1436_ _2949_ _2950_ _2939_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_117_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5495_ _3833_ _0266_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7216__I _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7234_ _2826_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6141__A1 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4446_ _3520_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6692__A2 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7165_ _2505_ _2791_ _2817_ _2820_ _2353_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4377_ _3749_ _3911_ _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _3547_ _1250_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7096_ _1616_ _2719_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6047_ _1759_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4455__A1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7998_ _0117_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6949_ _2505_ _2567_ _2610_ _2353_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5707__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7327__S _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6380__A1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6132__A1 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7880__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4694__A1 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7632__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4446__A1 _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6914__B _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4461__A4 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6199__A1 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7148__B1 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7699__A1 _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5265__B _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4921__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4300_ _3834_ _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_114_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4231_ as2650.carry _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7871__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6674__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4162_ as2650.r0\[1\] _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7623__A1 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4093_ _3529_ _3628_ _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8010__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7921_ _0040_ clknet_leaf_4_wb_clk_i as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7852_ _1202_ _1866_ _3453_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6803_ _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7783_ _1995_ _1343_ _2174_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4995_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _2274_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3946_ _3481_ _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6665_ _2326_ _2329_ _2330_ _2331_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__S _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5616_ _1387_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6596_ _1386_ _2263_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6901__A3 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5175__B _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5547_ _3569_ _3934_ _3585_ _3787_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__A1 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5478_ _3921_ _0346_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7390__B _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4429_ _3873_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7217_ _2870_ _3900_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7862__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7148_ _2121_ _2802_ _2803_ _1826_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7614__A1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7614__B2 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7079_ _2663_ _2736_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4428__A1 _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7090__A2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7549__C _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout51 net33 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7284__C _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5156__A2 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6353__A1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5085__B _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__A1 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__A2 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8033__CLK clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7605__A1 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5104__I _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4419__A1 _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4780_ _0629_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6592__A1 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_35_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5774__I _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6344__A1 _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _1279_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5401_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6895__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6381_ _2047_ _2049_ _1865_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _1160_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8120_ _0239_ clknet_leaf_61_wb_clk_i as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8051_ _0170_ clknet_leaf_10_wb_clk_i as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7844__A1 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4658__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7002_ _0782_ _3652_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4214_ _3517_ _3741_ _3747_ _3749_ _3750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5194_ _0988_ _1005_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4145_ as2650.r0\[0\] _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7072__A2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4076_ _3611_ _3491_ _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5083__A1 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7904_ _0023_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4830__A1 _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7835_ _2035_ _3385_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5885__S _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6583__A1 _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7766_ _3376_ _3377_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_127_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4978_ _0795_ _0814_ _0819_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7385__B _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6717_ as2650.addr_buff\[2\] _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7697_ _1801_ _2736_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5138__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6648_ _0894_ _1549_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6886__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5689__A3 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6579_ _1872_ _1944_ _2062_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4897__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8056__CLK clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7835__A1 _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6638__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5074__A1 as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7279__C _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5795__S _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__A1 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6877__A2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4888__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7826__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7314__I _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4673__I _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5950_ _1701_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _0746_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5881_ _1653_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7620_ _2649_ _3245_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4832_ _0649_ _0651_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6565__A1 _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4576__B1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7551_ _2570_ _3179_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4763_ _0591_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4040__A2 _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8079__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _2178_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7482_ _3066_ _3111_ _3112_ _3034_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4694_ _0453_ _0545_ _3824_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6868__A2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6433_ _2106_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6364_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5540__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6549__B _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8103_ _0222_ clknet_leaf_47_wb_clk_i as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5315_ _0661_ _0905_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4848__I _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6295_ _1990_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7224__I _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7916__CLK clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8034_ _0153_ clknet_leaf_14_wb_clk_i as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6096__A3 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5246_ _1078_ _1079_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5177_ _0935_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4128_ _3644_ _3661_ _3663_ _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_84_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5056__A1 _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__I _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4059_ _3559_ _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4803__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5851__I0 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7818_ _3767_ _3419_ _3159_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7749_ _0616_ _3361_ _3364_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4031__A2 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6308__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6859__A2 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7843__B _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7335__S _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5531__A2 _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6459__B _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7808__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7284__A2 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4098__A2 _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__A2 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4493__I _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6795__A1 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6795__B2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4270__A2 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5770__A2 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7939__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6369__B _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ _3548_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7275__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6080_ _1209_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _0864_ _0870_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _2346_ _2641_ _2642_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5933_ _1688_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_50_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4261__A2 _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5864_ _1604_ _1632_ _1643_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7647__C _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7603_ _1115_ _0774_ _3229_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4815_ _0573_ _0656_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5795_ _1589_ as2650.stack\[2\]\[4\] _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6123__I _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7534_ _1477_ _0516_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4746_ _3711_ _0500_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7663__B _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7465_ _1578_ _3002_ _3096_ _2127_ _3014_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4677_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6010__I0 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6416_ _2072_ _2076_ _2089_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ _2992_ _3028_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4167__I3 as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput17 net17 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput28 net28 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5183__B _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput39 net39 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6347_ _2032_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7266__A2 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6278_ _1943_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5277__A1 as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8017_ _0136_ clknet_leaf_45_wb_clk_i as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5229_ _1062_ _1045_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5029__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4252__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5752__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6001__I0 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5504__A2 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7257__A2 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5268__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7009__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6768__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6768__B2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6232__A3 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7193__A1 _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5983__S _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7732__A3 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4600_ _3821_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5580_ as2650.psl\[6\] _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6940__B2 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _3678_ _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7496__A2 _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7250_ _2872_ _0368_ _2868_ _2901_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4462_ _3896_ _0268_ _0269_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4149__I3 as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8117__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6201_ _1253_ _1896_ _1898_ _1272_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4393_ _3805_ _3926_ _3922_ _3819_ _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7181_ _2835_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6132_ as2650.addr_buff\[2\] _1837_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7248__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6063_ as2650.stack\[3\]\[10\] _1763_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__C _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5014_ _3721_ _0836_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4482__A2 _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _1521_ _2620_ _2625_ _2581_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6562__B _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5431__A1 _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _2121_ _2550_ _2558_ _2442_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6281__C _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3993__A1 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ _1539_ _1631_ _1633_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5893__S _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5778_ as2650.pc\[2\] _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7517_ net32 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4729_ _0580_ _3884_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7448_ _3075_ _3078_ _3079_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7379_ _3004_ _3012_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7613__S _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4101__I _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6737__B _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3940__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6998__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__A2 _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6922__A1 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6922__B2 _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6698__I _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6525__I1 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5489__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5107__I _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4464__A2 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6750_ _1683_ _2414_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3962_ as2650.ins_reg\[4\] _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5964__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3975__A1 _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5701_ _1351_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6681_ as2650.stack\[3\]\[1\] _2342_ _2343_ as2650.stack\[2\]\[1\] _2348_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5632_ _1438_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6913__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ _1354_ _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7302_ _2830_ _0790_ _2886_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7469__A2 _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4514_ _0338_ _0344_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_89_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5494_ _1298_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6677__B1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7233_ _2118_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4445_ _0299_ as2650.r123_2\[0\]\[3\] as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\]
+ _3478_ _3492_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6141__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7164_ _2271_ _2818_ _2819_ _2339_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4376_ _3840_ _3845_ _3910_ _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6557__B _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4856__I _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6115_ _1025_ _1823_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7095_ _1617_ _2244_ _2752_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6046_ _1765_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6292__B _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7997_ _0116_ clknet_leaf_38_wb_clk_i as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5404__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _2113_ _2606_ _2609_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6879_ _2538_ _2541_ _2116_ _1264_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7157__B2 as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7407__I _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6380__A2 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6311__I _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6132__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7343__S _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4143__A1 _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5891__A1 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6186__C _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7632__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__A1 as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6840__B1 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7298__B _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7396__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6199__A2 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7148__A1 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7148__B2 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4006__I _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6221__I _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__I0 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4134__A1 _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4230_ _3761_ _3763_ as2650.psl\[3\] as2650.carry _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_99_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7871__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4685__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4161_ as2650.r123\[1\]\[1\] as2650.r123_2\[1\]\[1\] _3477_ _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7084__B1 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ _3625_ _3627_ _3628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5634__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7920_ _0039_ clknet_leaf_52_wb_clk_i as2650.r123\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7851_ _3536_ _1872_ _3451_ _3452_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _1586_ _2465_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7782_ _3855_ _3639_ _3644_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4994_ _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6733_ _2377_ _2388_ _2398_ _2049_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7139__A1 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3945_ _3480_ _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6664_ _1358_ _1811_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ _0976_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6595_ _1975_ _2258_ _2262_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5175__C _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5546_ _3537_ _1350_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_117_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5477_ _1284_ _3813_ _3818_ _3761_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7311__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6114__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7216_ _2075_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4428_ _3877_ _3690_ _3706_ _0282_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_120_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6287__B _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5191__B _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7147_ _2482_ _2760_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4359_ _3893_ _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7614__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7078_ _2252_ _2313_ _2383_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5625__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6029_ _1732_ _1741_ _1754_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_74_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4535__B _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7378__A1 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6306__I _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout52 net29 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6353__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__A1 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6105__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7972__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5864__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7369__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6216__I _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_90 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_60_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6041__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6592__A2 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7541__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6344__A2 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__S _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5400_ _3565_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6380_ _2050_ _2055_ _2058_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5331_ _0874_ _1162_ _1163_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5790__I as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8050_ _0169_ clknet_leaf_10_wb_clk_i as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5262_ _0669_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7844__A2 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5855__A1 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7001_ _2422_ _2657_ _2660_ _2464_ _2475_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4658__A2 _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _3748_ _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _0987_ _1008_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4144_ as2650.r123\[1\]\[0\] as2650.r123_2\[1\]\[0\] as2650.psl\[4\] _3680_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6327__S _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4075_ _3594_ _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6280__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout50_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7903_ _0022_ clknet_leaf_5_wb_clk_i as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7834_ _1843_ _2023_ _3438_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5030__I _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7765_ _2108_ _2507_ _2510_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4977_ as2650.r123\[1\]\[7\] _0815_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6583__A2 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6716_ _2380_ _2361_ _2371_ _2381_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7696_ _2987_ _3318_ _2137_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6647_ _2313_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4346__A1 _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7995__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4897__A2 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6796__I _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5529_ _1332_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7835__A2 _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4821__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7771__A1 _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6326__A2 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7523__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8000__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4888__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7826__A2 _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4954__I _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6262__A1 _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ _0747_ _0748_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_74_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ _1653_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7486__B _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _3723_ _0660_ _0681_ _0412_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__I _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__B _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7762__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7550_ _3127_ _3129_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4762_ _0524_ _0613_ _0333_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6501_ _2177_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7481_ _1472_ _3066_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7514__A1 _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6317__A2 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4693_ _0535_ _0544_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5376__I0 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6432_ _1527_ _1857_ _2111_ _2114_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4879__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6363_ _1782_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8102_ _0221_ clknet_leaf_48_wb_clk_i as2650.stack\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5314_ _0406_ _0992_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6294_ _1241_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8033_ _0152_ clknet_leaf_21_wb_clk_i as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5245_ _1000_ _1036_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__I _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ _0972_ _0942_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4500__B2 _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ _3662_ _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_110_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6253__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4058_ _3593_ _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7817_ _3416_ _3417_ _3423_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7753__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6556__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8023__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4567__A1 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7748_ _0500_ _3362_ _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7679_ _1914_ _3299_ _3301_ _3302_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6308__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3943__I _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7269__B1 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7808__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5295__A2 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6492__A1 _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6922__C _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5030_ _0829_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5038__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6981_ as2650.stack\[3\]\[7\] _2604_ _2535_ as2650.stack\[0\]\[7\] _2642_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5932_ as2650.pc\[5\] _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8046__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ as2650.stack\[6\]\[7\] _1637_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6538__A2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4633__B _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7602_ _3205_ _3208_ _3228_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4814_ _0529_ _0571_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5794_ _1566_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7533_ net51 _3161_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _0466_ _0467_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7663__C _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7464_ _2372_ _3093_ _3095_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4676_ _0503_ _0504_ _0526_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_107_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6415_ _1796_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7395_ _2048_ _2303_ _3027_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6710__A2 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput18 net18 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput29 net29 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4721__A1 _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6346_ _2034_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6277_ _1973_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8016_ _0135_ clknet_leaf_36_wb_clk_i as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5228_ _1033_ _1039_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5159_ _0994_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7838__C _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7726__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6465__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8069__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6217__A1 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6768__A2 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4779__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5440__A2 _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7717__A1 _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7906__CLK clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7193__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7732__A4 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7764__B _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6940__A2 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4530_ _0305_ _0383_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4679__I as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4461_ _0312_ _3693_ _0314_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_102_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6200_ _1897_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4703__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7180_ _0802_ _1229_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4392_ _3803_ _3816_ _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6131_ _1460_ _1832_ _1838_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A1 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _1732_ _1761_ _1774_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _0841_ _0851_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6759__A2 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6964_ _2579_ _2614_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5431__A2 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1674_ _1675_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7708__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6895_ _1270_ _2493_ _2497_ _2557_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6134__I _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3993__A2 _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5846_ as2650.stack\[6\]\[0\] _1632_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5973__I _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5777_ _1575_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_3_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7516_ _2827_ _3137_ _3145_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4728_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7447_ _3075_ _3078_ _3044_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4659_ _0281_ _0491_ _0511_ _3722_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6695__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5498__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7378_ _1894_ _3007_ _3011_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6329_ _0407_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6447__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4473__A3 _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7849__B _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7929__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7584__B _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__A1 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6922__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4528__A4 _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4933__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5110__A1 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _3496_ _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5700_ _1253_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3975__A2 _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ as2650.stack\[1\]\[1\] _1547_ _1714_ as2650.stack\[0\]\[1\] _2347_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5631_ _1324_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5793__I _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6913__A2 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ _1357_ _1363_ _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_129_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ _2870_ _0774_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4513_ _0365_ _0366_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5493_ _3764_ _1286_ _1291_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7232_ _2857_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4444_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7163_ as2650.stack\[1\]\[12\] _2811_ _2814_ as2650.stack\[0\]\[12\] _2819_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4375_ _3892_ _3902_ _3908_ _3909_ _3516_ _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_113_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6557__C _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6114_ _0311_ _1324_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7094_ _2243_ _2750_ _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _1681_ as2650.stack\[3\]\[2\] _1763_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6129__I _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7669__B _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5968__I _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6065__S _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7996_ _0115_ clknet_leaf_38_wb_clk_i as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6292__C _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6601__A1 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5404__A2 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6601__B2 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6947_ _2513_ _2607_ _2608_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6878_ _2513_ _2539_ _2540_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _1617_ _1568_ _1618_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4143__A2 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7423__I _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6039__I _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6840__A1 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5643__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6840__B2 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7396__A2 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8107__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6659__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4509__I1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4957__I _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5331__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5882__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4160_ _3678_ _3692_ _3695_ _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4091_ _3500_ _3541_ _3626_ _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_110_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5634__A2 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7850_ _1217_ _1226_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6801_ _1581_ _2414_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5398__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4445__I0 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4993_ _3618_ _0833_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7781_ _1270_ _1299_ _2221_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6732_ _2393_ _2395_ _2397_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3944_ _3479_ _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7139__A2 _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6663_ _1415_ _1875_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5614_ _1414_ _1416_ _1419_ _1421_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6594_ _1412_ _2260_ _2261_ _1826_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5545_ _1228_ _1352_ _1207_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5570__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5476_ _3805_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7311__A2 _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4427_ _3689_ _3706_ _3878_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7215_ _2868_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7146_ _2548_ _2799_ _2800_ _2801_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4358_ _3687_ _3705_ _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7075__A1 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7077_ _2001_ _2730_ _2732_ _2308_ _2734_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_58_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4289_ _3752_ _3809_ _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6822__A1 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6028_ as2650.stack\[0\]\[9\] _1743_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6822__B2 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5698__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7378__A2 _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__A1 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7979_ _0098_ clknet_leaf_31_wb_clk_i as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4107__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7418__I _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5561__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7302__A2 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5864__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7066__A1 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6813__A1 _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5401__I _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7369__A2 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7613__I0 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_80 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_91 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__4017__I _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7541__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5330_ _0867_ _1162_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4687__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _0507_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7063__I _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7000_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5855__A2 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4212_ _3563_ _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5192_ _0559_ _0903_ _0943_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_44_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7057__A1 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4143_ _3498_ _3505_ _3506_ _3679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6804__A1 as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4074_ _3599_ _3609_ _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7902_ _0021_ clknet_leaf_7_wb_clk_i as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6280__A2 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4291__A1 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7833_ _1204_ _1254_ _1873_ _3437_ _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_52_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7666__C _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4043__A1 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7764_ _2812_ _2815_ _2409_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4976_ _0713_ _0814_ _0818_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5467__B _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6715_ _1877_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7695_ net39 _3317_ _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_138_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6142__I _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6646_ as2650.addr_buff\[1\] _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7682__B _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6591__I0 as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6740__B1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6577_ _1821_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5528_ _1333_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7296__A1 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5459_ _1017_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5846__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7048__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7129_ _2375_ _2785_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6023__A2 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7220__A1 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4034__A1 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__I0 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7523__A2 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7287__A1 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4300__I _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7039__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6262__A2 _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5131__I _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_2_0_wb_clk_i clknet_3_5_0_wb_clk_i clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7767__B _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4830_ _3722_ _0676_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4025__A1 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6565__A3 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _0592_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4576__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6500_ _2171_ _2173_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7480_ _1420_ _0376_ _3110_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _0444_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6431_ _3672_ _2109_ _2113_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5376__I1 as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7933__D _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6362_ as2650.cycle\[0\] _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8101_ _0220_ clknet_leaf_39_wb_clk_i as2650.stack\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5313_ _1061_ _1145_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7278__A1 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6293_ _1338_ _1891_ _1988_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_88_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5828__A2 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__I _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8032_ _0151_ clknet_leaf_17_wb_clk_i as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5244_ _1000_ _1036_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _0984_ _0985_ _1011_ _0941_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4500__A2 _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _3643_ as2650.carry _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_84_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ as2650.ins_reg\[3\] _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7677__B _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7816_ _3419_ _3422_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7962__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6556__A3 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7747_ _0521_ _3361_ _3363_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5764__A1 _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _0807_ _0805_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7678_ _1833_ as2650.addr_buff\[1\] _1801_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6308__A3 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _1986_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7269__A1 _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7269__B2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6492__A2 _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6047__I _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6180__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4730__A2 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4030__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7680__B2 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6980_ as2650.stack\[1\]\[7\] _2603_ _2601_ as2650.stack\[2\]\[7\] _2641_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7985__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _1687_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ _1600_ _1631_ _1642_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7196__B1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7601_ _1097_ _0660_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4813_ _0653_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6943__B1 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5793_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7532_ _3147_ _3149_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4744_ _0406_ _3838_ _0416_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7463_ _1577_ _3094_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4675_ _3522_ _0502_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6414_ _1338_ _1342_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7394_ _2315_ _3026_ _2994_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput19 net19 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_143_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4721__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6345_ _2033_ _0531_ _2026_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5036__I _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6276_ _3846_ _1548_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7671__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5227_ _1040_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8015_ _0134_ clknet_leaf_45_wb_clk_i as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6474__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5682__B1 _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5158_ _0991_ _0993_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109_ as2650.r0\[7\] _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5029__A3 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6226__A2 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5089_ _0321_ _0837_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7726__A2 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8140__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3954__I _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6162__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4173__B1 _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7662__A1 _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7414__A1 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6217__A2 _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4228__A1 _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6505__I _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7717__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7193__A3 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4951__A2 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6240__I _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4460_ _3603_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5900__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4391_ _3921_ _3924_ _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ _1836_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7653__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6061_ as2650.stack\[3\]\[9\] _1763_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6456__A2 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8013__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _3715_ _0840_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _1602_ _2623_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5967__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6415__I _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5914_ _1541_ _1544_ _1564_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6894_ _2554_ _2556_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7708__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__A1 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5845_ _1630_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6351__S _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7674__C _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__A1 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5195__A2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5776_ _1573_ as2650.stack\[2\]\[1\] _1574_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7515_ _1480_ _3032_ _3033_ _3144_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4727_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6144__A1 _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7446_ _3076_ _3077_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4658_ _0492_ _3632_ _3850_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7377_ _1918_ _1908_ _2225_ _3010_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_104_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6328_ _2019_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7644__A1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6447__A2 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6259_ _1944_ _1952_ _1954_ _1332_ _1955_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4458__A1 _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5655__B1 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__A4 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4554__B _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4630__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4697__B2 _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7635__A1 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A2 _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3960_ _3495_ _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5630_ _3560_ _1436_ _1298_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5177__A2 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5561_ _0727_ _1364_ _1366_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7300_ _1380_ _2865_ _2947_ _2948_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6126__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4512_ _3937_ _0345_ _3755_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5492_ _1299_ _3818_ _1288_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7231_ _2189_ _2865_ _2874_ _2884_ _2131_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6677__A2 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7874__A1 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4443_ as2650.r123\[0\]\[3\] _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4374_ _3901_ _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7162_ as2650.stack\[3\]\[12\] _2812_ _2815_ as2650.stack\[2\]\[12\] _2818_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_99_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7626__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6113_ _1498_ _1821_ _1554_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7093_ _0807_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6044_ _1764_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6854__B _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7995_ _0114_ clknet_leaf_40_wb_clk_i as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6145__I _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ as2650.stack\[5\]\[6\] _2603_ _2604_ as2650.stack\[7\]\[6\] _2608_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4612__A1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6877_ as2650.stack\[4\]\[5\] _2535_ _2400_ as2650.stack\[6\]\[5\] _2540_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5828_ as2650.stack\[2\]\[10\] _1574_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6365__A1 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5759_ _3600_ _0938_ _1558_ _1551_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8059__CLK clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6117__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7865__A1 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7429_ _3013_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4143__A3 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4851__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4603__A1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4303__I _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6659__A2 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7084__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _3558_ _3559_ _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5095__A1 as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4842__A1 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6800_ _2363_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7780_ _2927_ _2931_ _3387_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6595__A1 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4992_ _3483_ _0823_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4445__I1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6731_ _2331_ _2396_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3943_ _3478_ _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6662_ _2327_ _2328_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _3667_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4213__I _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5544_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5570__A2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5475_ _0261_ _0353_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7919__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7214_ _2867_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4426_ _3718_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5472__C _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7145_ _1520_ _2797_ _1211_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4357_ _3843_ _3716_ _3851_ _3891_ _3892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7075__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7076_ _1703_ _2733_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4288_ _3818_ _3822_ _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5086__A1 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6822__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ _1753_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5389__A2 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6586__A1 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7978_ _0097_ clknet_leaf_45_wb_clk_i as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _0578_ _2552_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4832__B _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__A1 _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4123__I _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6759__B _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3962__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7434__I _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7066__A2 _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A1 _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6813__A2 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4824__A1 _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7613__I1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_70 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_81 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_92 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6513__I _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4033__I _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7829__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5260_ _1058_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4211_ _3742_ _3745_ _3746_ _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5191_ _1022_ _1026_ _0903_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7057__A2 _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4142_ _3620_ _3677_ _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5799__I _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6804__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4073_ _3604_ _3608_ _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7901_ _0020_ clknet_leaf_6_wb_clk_i as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4291__A2 _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_13_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7832_ _2006_ _1348_ _3436_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6568__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7763_ _3373_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4975_ as2650.r123\[1\]\[6\] _0815_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6714_ _1942_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4144__S as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6423__I _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7694_ _3316_ _3295_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6645_ _2310_ _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5039__I _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6576_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6591__I1 as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6579__B _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5527_ _3529_ _1334_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7296__A2 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5458_ _1266_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7891__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4409_ _3755_ _3921_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5389_ _3496_ _3504_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7128_ _2408_ _2755_ _2784_ _2456_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5059__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7059_ _2243_ _2717_ _2461_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4806__A1 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4282__A2 _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7220__A2 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7429__I _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5231__A1 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3957__I _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4034__A2 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6731__A1 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6489__B _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7039__A2 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6508__I _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6798__A1 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4025__A2 _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6565__A4 _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4760_ _0593_ _0611_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4691_ _0342_ _0349_ _0442_ _0345_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6722__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5525__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6361_ _1248_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8100_ _0219_ clknet_leaf_32_wb_clk_i as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _1064_ _1088_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7278__A2 _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6292_ _1373_ _1805_ _1824_ _1865_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5289__A1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8031_ _0150_ clknet_leaf_17_wb_clk_i as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ _1035_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5174_ _0986_ _1007_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4125_ _3660_ _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6789__A1 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4056_ _3585_ _3591_ _3556_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_83_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7815_ _3420_ _3421_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4016__A2 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6153__I _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7746_ _0394_ _3362_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4958_ _3513_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5764__A2 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7677_ _3249_ _3251_ _2069_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4889_ _3939_ _0736_ _0738_ _0262_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_6628_ _1539_ _2244_ _2295_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6713__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _1958_ _2226_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7269__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4557__B _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5452__A1 _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4292__B _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6952__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5407__I _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5343__S _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5691__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5930_ as2650.stack\[1\]\[4\] _1685_ _1686_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5994__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ as2650.stack\[6\]\[6\] _1637_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7196__A1 _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7196__B2 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7600_ _1449_ _3040_ _2069_ _3226_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_61_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4812_ _0532_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5792_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6943__A1 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7531_ _3158_ _3160_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4743_ _0468_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7462_ _3023_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4674_ _0499_ _3616_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6413_ _2088_ _2093_ _2096_ _1896_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4706__B1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7393_ _0940_ _3025_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4221__I _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4182__A1 _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6344_ _1846_ _2032_ _1268_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5761__B _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7120__A1 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6275_ _1969_ _1971_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7120__B2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8014_ _0133_ clknet_leaf_48_wb_clk_i as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5226_ _1059_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7671__A2 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5682__A1 as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6148__I _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5682__B2 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5157_ _0991_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5052__I _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4108_ _3643_ _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6226__A3 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5088_ _0280_ _0898_ _0881_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4237__A2 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4039_ _3540_ _3574_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7187__A1 _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6934__A1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7729_ _2798_ _3350_ _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6162__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4131__I _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7662__A2 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7414__A2 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6217__A3 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5728__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4951__A3 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4164__A1 _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4390_ _3813_ _3923_ _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5900__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7102__A1 _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7952__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7653__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6060_ _1773_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input8_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5011_ _0832_ _0836_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6962_ _1598_ _2577_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5967__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__I _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3978__A1 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5913_ as2650.stack_ptr\[1\] _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6893_ _2059_ _2555_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7708__A3 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4216__I _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5844_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3993__A4 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4660__B _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5775_ _1565_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7514_ _3071_ _3143_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4726_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7445_ _1417_ _0321_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6144__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4657_ _3890_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__I _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7376_ _1266_ _1201_ _3003_ _1933_ _3009_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4588_ as2650.holding_reg\[4\] _0440_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6327_ _2018_ _3917_ _2005_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6258_ _1386_ _1348_ _1878_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4458__A2 _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _1043_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5655__B2 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _3543_ _1240_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5510__I _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4630__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5666__B _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7332__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4146__A1 _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7975__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7105__C _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6516__I _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5420__I _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7020__B1 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _3595_ _3491_ _1367_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_38_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4511_ _0351_ _0362_ _0364_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7791__B _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6126__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5491_ _1267_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7230_ _2188_ _2162_ _2883_ _1442_ _2864_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4137__A1 _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4442_ _0296_ _3615_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4688__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7161_ _2346_ _2813_ _2816_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4373_ _3906_ _3907_ _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7087__B1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6112_ _3569_ _1784_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7092_ _2720_ _2728_ _2749_ _2459_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6043_ _1679_ as2650.stack\[3\]\[1\] _1763_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6426__I _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7994_ _0113_ clknet_leaf_41_wb_clk_i as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6062__A1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ as2650.stack\[4\]\[6\] _2508_ _2601_ as2650.stack\[6\]\[6\] _2607_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ as2650.stack\[5\]\[5\] _1547_ _1651_ as2650.stack\[7\]\[5\] _2539_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5827_ _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6365__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _1249_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4915__A3 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4709_ _0402_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6117__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5689_ _1434_ _1437_ _1441_ _1443_ _1495_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_108_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4128__A1 _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7428_ net30 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7865__A2 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7359_ _2581_ _2333_ _2992_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7617__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5628__A1 _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4851__A2 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7876__B _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4603__A2 _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6071__I _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8003__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4367__A1 _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7305__A1 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4119__A1 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7608__A2 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6292__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4842__A2 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7241__B1 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4991_ _0831_ _0313_ _0315_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_90_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5398__A3 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7792__A1 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6730_ _1418_ _1875_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3942_ _3477_ _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6661_ net5 _2259_ _2325_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5612_ _0388_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6592_ _1816_ _2259_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5543_ _3673_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5474_ _0727_ _3661_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7213_ _1331_ _2000_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4425_ _0279_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5325__I _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7144_ _2365_ _2790_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4530__A1 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4356_ _3852_ _3854_ _3889_ _3890_ _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7075_ _1613_ _2701_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4287_ _3792_ _3766_ _3822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5086__A2 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6283__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6026_ _1696_ as2650.stack\[0\]\[8\] _1748_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6156__I _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7696__B _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7977_ _0096_ clknet_leaf_33_wb_clk_i as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6586__A2 _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__A3 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7783__A1 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8026__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _2589_ _2587_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ _1689_ _2359_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7535__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5010__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6510__A2 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4521__A1 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5077__A2 _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__B _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4824__A2 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_60 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7774__A1 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_71 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_45_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_82 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4588__A1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_93 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7526__A1 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5001__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5346__S _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7829__A2 _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4210_ _3516_ _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4512__A1 _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1024_ _1025_ _0588_ _0858_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4141_ _3673_ _3676_ _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6265__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4072_ _3543_ _3607_ _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4815__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7900_ _0019_ clknet_leaf_6_wb_clk_i as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7831_ _0803_ _1465_ _1256_ _1507_ _1200_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_97_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6568__A2 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7765__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__A1 _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4974_ _0616_ _0814_ _0817_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7762_ _2899_ _3374_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6713_ _1577_ _2310_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7693_ net38 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6644_ _1571_ _1672_ _2309_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6575_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6740__A2 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5526_ _3541_ _0358_ _3552_ _3810_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5457_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4408_ _3939_ _0261_ _0262_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5388_ _3575_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6595__B _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7127_ _1218_ _2780_ _2783_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4339_ _3873_ _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7058_ _2690_ _2696_ _2716_ _2459_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4806__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6009_ _1738_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6008__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7756__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6559__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5231__A2 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4034__A3 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7508__A1 _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6731__A2 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6495__A1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7113__C _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7747__A1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7909__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4025__A3 _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _0436_ _0538_ _0541_ _3919_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_81_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4733__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6360_ _1338_ _2043_ _2045_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5311_ _1064_ _1088_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6291_ _1986_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8030_ _0149_ clknet_leaf_17_wb_clk_i as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6486__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7304__B _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5173_ _0868_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4124_ _3659_ _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4219__I _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4055_ _3586_ _3587_ _3588_ _3590_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_83_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7738__A1 _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7814_ _1379_ _0883_ _1401_ _2839_ _1319_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6410__A1 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7745_ _3355_ _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4957_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4421__B1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4972__A1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7676_ _1913_ _2736_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4888_ _0737_ _0720_ _3935_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6627_ _1884_ _2294_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _0939_ _1971_ _1786_ _1788_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ _1307_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6489_ _1503_ _2160_ _2166_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6477__A1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6609__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4557__C _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6229__A1 _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4129__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5452__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7729__A1 _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6401__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__A1 as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7175__I _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6180__A3 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6640__A1 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5860_ _1595_ _1631_ _1641_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7196__A2 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _1586_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6943__A2 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7530_ _3147_ _3058_ _3159_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4742_ _0474_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7461_ _3090_ _3092_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4673_ _3634_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6203__B _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4502__I _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6412_ _2089_ _2095_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4706__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7392_ net52 net28 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4706__B2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6343_ _1382_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4182__A2 _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__C _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6459__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5761__C _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6274_ _1558_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4658__B _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8013_ _0132_ clknet_leaf_31_wb_clk_i as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5225_ _1043_ _1044_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6429__I _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5682__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5156_ _3712_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4107_ as2650.psl\[3\] _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ _3708_ _0885_ _0925_ _0839_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ _3558_ _3559_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5489__B _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5198__A1 _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6934__A2 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5989_ as2650.stack\[5\]\[7\] _1724_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7728_ _1624_ _3094_ _3092_ _3349_ _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4945__A1 _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7659_ _1836_ _3252_ _2075_ _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4412__I _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5370__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6767__C _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6622__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6074__I _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7119__B _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6689__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4322__I _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4951__A4 _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A2 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _3664_ _0842_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6861__A1 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7789__B _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6961_ _2464_ _2615_ _2621_ _2475_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5912_ _1672_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3978__A2 _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _2551_ _2494_ _2553_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5843_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6916__A2 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4927__A1 _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5774_ _1572_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7029__B _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7513_ _1479_ _0517_ _3142_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4725_ net1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5328__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7444_ _0317_ _0320_ _0288_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4656_ _0403_ _0306_ _0497_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4587_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7375_ _1981_ _3008_ _2236_ _1822_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6326_ _0289_ _2015_ _2017_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6257_ _1953_ _1896_ _1550_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_103_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6852__A1 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ _3834_ as2650.r123_2\[0\]\[4\] _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5655__A2 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ _1885_ _3587_ _3588_ _3590_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_130_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ _0495_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4091__A1 _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4918__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4394__A2 _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6778__B _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4146__A2 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3981__I _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7453__I _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5701__I _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4317__I _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8082__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5576__C _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7571__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5582__A1 _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ _3934_ _0363_ _3916_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _1295_ _1297_ _1273_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5334__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4441_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4987__I _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4137__A2 _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7160_ as2650.stack\[4\]\[12\] _2814_ _2815_ as2650.stack\[6\]\[12\] _2816_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4372_ _3894_ _3905_ _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _1815_ _1817_ _1818_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7091_ _2740_ _2727_ _2748_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6042_ _1758_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5611__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7993_ _0112_ clknet_leaf_38_wb_clk_i as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6062__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6944_ _2506_ _2602_ _2605_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6875_ _2506_ _2536_ _2537_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7011__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5826_ as2650.pc\[10\] _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5573__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5058__I _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _1555_ _1556_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4708_ _0499_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5688_ _1399_ _1494_ _1410_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7427_ _3020_ _3057_ _3059_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4128__A2 _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _0392_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7358_ _2991_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _1526_ _1335_ _1999_ _2001_ _2002_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7289_ _2870_ _0660_ _2886_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7250__A1 _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3976__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7002__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7942__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4367__A2 _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5564__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4119__A2 as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4600__I _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5867__A2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6816__A1 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7241__A1 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4990_ _3542_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4445__I3 as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3941_ as2650.psl\[4\] _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7358__I _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6660_ _1817_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4358__A2 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5555__A1 _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\] _3481_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5542_ _1196_ _1349_ _3577_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5473_ _0737_ _0727_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6355__I0 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7093__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6211__B _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5606__I _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4424_ _0278_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7212_ _1970_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7143_ as2650.addr_buff\[4\] _2385_ _2499_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4355_ _3630_ _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7074_ _2396_ _2731_ _2381_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4286_ _3808_ _3779_ _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7480__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6283__A2 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6025_ _1603_ _1741_ _1752_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4046__A1 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7976_ _0095_ clknet_leaf_46_wb_clk_i as2650.stack\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7965__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7783__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6927_ _0668_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6172__I _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6858_ _2463_ _2521_ _2045_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7535__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6105__C _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5809_ as2650.pc\[7\] _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_50_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5546__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6789_ _2282_ _2452_ _2453_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5516__I _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7471__A1 _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6347__I _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4285__A1 _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5482__B1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7223__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_61 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7774__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_72 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_83 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7526__A2 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8120__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5537__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6810__I _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5426__I _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ _3674_ _3675_ _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6265__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _3605_ _3606_ _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4276__A1 _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7988__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7830_ _3434_ _3435_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7765__A2 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7761_ _1711_ _3373_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4973_ as2650.r123\[1\]\[5\] _0815_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6206__B _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4505__I _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6712_ _2307_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7692_ _3018_ _3314_ _3315_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6643_ _1537_ _2309_ _1571_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6574_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7037__B _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_22_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5525_ _3628_ _1310_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4240__I _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5456_ _3490_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4407_ _3782_ _3574_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4503__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5700__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5387_ _0820_ _3497_ _3535_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_120_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7126_ _2271_ _2781_ _2782_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _3872_ _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7057_ _2695_ _2707_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4269_ _3803_ _3624_ _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6008_ _1709_ _1740_ _1742_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6008__A2 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7205__A1 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7205__B2 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7756__A2 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7959_ _0078_ clknet_leaf_42_wb_clk_i as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5519__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6630__I _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5690__B _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7692__A1 _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6495__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6077__I _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4325__I _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4025__A4 _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6183__A1 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4733__A2 _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5310_ _1127_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _1279_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5241_ _1065_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8016__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5172_ _0920_ _0955_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_123_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7435__A1 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4123_ _3658_ _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6238__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4054_ as2650.cycle\[6\] _3528_ _3589_ _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_68_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4944__B _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6715__I _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7738__A2 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7813_ _3385_ _2008_ _2007_ _1445_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6946__B1 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6410__A2 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7744_ _3353_ _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4956_ _0801_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4421__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4421__B2 _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7675_ _3257_ _3259_ _2826_ _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _0717_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__I _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6626_ _1673_ _2127_ _2292_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6557_ _2222_ _1865_ _1903_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ _0769_ _1312_ _1315_ _1311_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6488_ _2108_ _2162_ _2165_ _2046_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7674__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_opt_1_1_wb_clk_i_I clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7674__B2 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ as2650.halted _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7426__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6229__A2 _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ _2765_ _2724_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8089_ _0208_ clknet_leaf_4_wb_clk_i as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5988__A1 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6625__I _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5452__A3 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A1 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6401__A2 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4145__I as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6165__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6468__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7665__A1 _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7417__A1 _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6640__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4651__A1 _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4810_ _0564_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ as2650.pc\[4\] _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4741_ _0475_ _0476_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__I _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7460_ _3091_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4672_ _3841_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6203__C _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6411_ _1521_ _2094_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5903__A1 as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4706__A2 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7391_ _3023_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6342_ _2031_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7105__B1 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7656__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6459__A2 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6273_ _1969_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8012_ _0131_ clknet_leaf_31_wb_clk_i as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5224_ _1041_ _1042_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7408__A1 _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ as2650.r123_2\[0\]\[4\] _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4106_ _3641_ _3642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5086_ _0306_ _0889_ _0884_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4037_ _3568_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5198__A2 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A1 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5988_ _1600_ _1717_ _1729_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7727_ _2583_ _3338_ _3348_ _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4945__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4939_ _3659_ _0488_ _0772_ _3895_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6147__A1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7658_ _3034_ _3282_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6609_ _1546_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7589_ _3016_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_1_0_wb_clk_i clknet_3_5_0_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_101_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7647__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7225__B _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5524__I _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3979__I _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6622__A2 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4633__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4936__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7119__C _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6689__A2 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7638__A1 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7638__B2 _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6974__B _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6861__A2 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7789__C _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6613__A2 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7810__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6960_ _2306_ _2620_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5911_ _1536_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6891_ _2551_ _2494_ _2553_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ _1547_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5773_ _1571_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4927__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5609__I _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7512_ _3140_ _3141_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4724_ _0532_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7443_ _1459_ _3898_ _3899_ _3041_ _3042_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XANTENNA__7877__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4655_ _3694_ _0507_ _0403_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7374_ _1789_ _1504_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4586_ _0397_ _0398_ _0437_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_115_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6325_ _2016_ _1446_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6256_ _1352_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _1041_ _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_76_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6187_ as2650.cycle\[7\] _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4863__A1 as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5138_ _0973_ _0974_ _0858_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _0908_ _0867_ _0905_ _3742_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4091__A2 _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__C _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4918__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4423__I _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A2 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7868__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6778__C _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7096__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4606__A1 _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7020__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5582__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ _0294_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4137__A3 _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4371_ _3894_ _3905_ _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6110_ _1498_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7087__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7090_ _2339_ _2720_ _2747_ _2456_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _1709_ _1760_ _1762_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7992_ _0111_ clknet_leaf_31_wb_clk_i as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6598__A1 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6943_ as2650.stack\[1\]\[6\] _2603_ _2604_ as2650.stack\[3\]\[6\] _2605_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4952__B _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5270__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6874_ as2650.stack\[3\]\[5\] _2507_ _2510_ as2650.stack\[2\]\[5\] _2537_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ _1614_ _1568_ _1615_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5022__A1 _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4243__I _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5756_ as2650.cycle\[2\] _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5573__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6879__B _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5687_ _1445_ _1493_ _1394_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7426_ net52 _3058_ _2751_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4638_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7894__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7357_ _2053_ _1385_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4569_ _0418_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6308_ _0860_ _1362_ _1888_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7288_ _2070_ _0679_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5089__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _1871_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6589__A1 _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7250__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4862__B _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6633__I _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7002__A2 _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4153__I _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6761__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3992__I _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7069__A2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4827__B2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4328__I _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7241__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4055__A2 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ net26 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5004__A1 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5610_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6752__A1 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6590_ _2253_ _1852_ _2256_ _1877_ _2257_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5555__A2 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ _1203_ _1247_ _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5472_ _1193_ _1262_ _1278_ _1280_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6355__I1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7211_ _2864_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4423_ _3861_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7142_ _2721_ _2797_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4354_ _3857_ _3874_ _3887_ _3888_ _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6718__I _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7073_ as2650.addr_buff\[2\] _2385_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4285_ _3818_ _3819_ _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5622__I _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6024_ as2650.stack\[0\]\[7\] _1746_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7480__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7975_ _0094_ clknet_leaf_48_wb_clk_i as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4046__A2 _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _1454_ _2587_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6857_ _2476_ _2504_ _2520_ _2293_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout46 net48 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6043__I0 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5808_ _1600_ _1567_ _1601_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6788_ as2650.stack\[3\]\[3\] _2445_ _2287_ as2650.stack\[0\]\[3\] _2453_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5739_ _1538_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7409_ _1459_ _3893_ _3897_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__8072__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__B _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7471__A2 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5482__B2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3987__I _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6363__I _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_62 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_73 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_84 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6982__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6034__I0 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__B1 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__C _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ as2650.addr_buff\[5\] _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4276__A2 _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4058__I _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6273__I _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7765__A3 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7760_ _2230_ _3367_ _3371_ _3372_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4972_ _0521_ _0814_ _0816_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _2060_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7691_ net38 _3217_ _1883_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6642_ _1206_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6725__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5528__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6573_ _1892_ _2225_ _2233_ _2240_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_121_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5617__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8095__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5524_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7150__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_62_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4406_ as2650.holding_reg\[2\] _3872_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5700__A2 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5386_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6448__I _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7125_ as2650.stack\[7\]\[11\] _2342_ _2272_ as2650.stack\[4\]\[11\] _2782_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4337_ _3871_ _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__I0 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7932__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7056_ _2339_ _2690_ _2714_ _2456_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4268_ as2650.holding_reg\[1\] _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6007_ as2650.stack\[0\]\[0\] _1741_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4199_ as2650.idx_ctrl\[1\] _3734_ _3735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7205__A2 _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5216__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7958_ _0077_ clknet_leaf_38_wb_clk_i as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _1593_ _1483_ _2570_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7889_ _0008_ clknet_leaf_61_wb_clk_i as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4431__I _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6495__A3 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6358__I _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__I _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6955__A1 as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A2 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6183__A2 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4194__A1 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7132__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7955__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5240_ _1066_ _1067_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5694__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5171_ _1006_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ _3645_ _3617_ _3654_ _3523_ _3657_ _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_57_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4053_ _3485_ _3486_ _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5997__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4944__C _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7199__A1 _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7199__B2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8135__D _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7812_ _3396_ _3418_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7743_ _0430_ _3354_ _3360_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4955_ _0803_ _3534_ _3841_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4421__A2 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7674_ _1703_ _3024_ _3184_ _3297_ _1319_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4886_ _0717_ _0720_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7048__B _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6625_ _2241_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7371__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4251__I _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6556_ _1359_ _1366_ _2223_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5507_ _1313_ _1314_ _1113_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6487_ _1025_ _2162_ _1797_ _2164_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__7123__A1 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _1246_ _3581_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5685__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4488__A2 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6178__I _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5369_ as2650.r123_2\[1\]\[1\] _1183_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7108_ _2722_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7426__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8088_ _0207_ clknet_leaf_63_wb_clk_i as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8110__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7039_ _2380_ _2694_ _2697_ _1953_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5810__I _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5988__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7230__C _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5031__B _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4426__I _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5685__C _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7362__A1 _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6165__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7978__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__A1 _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4479__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6873__B1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7417__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7421__B _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6928__A1 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7050__B1 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4740_ _0424_ _0477_ _0480_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4671_ _3517_ _0523_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6410_ _1881_ _1959_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7390_ _1232_ _2305_ _2473_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5903__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _2030_ as2650.holding_reg\[4\] _2026_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7105__A1 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6272_ _1968_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8133__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5667__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8011_ _0130_ clknet_leaf_49_wb_clk_i as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5223_ _1056_ _1057_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4714__I0 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5154_ _0948_ _0989_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4955__B _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4105_ _3638_ _3640_ _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5085_ _0288_ _0848_ _0889_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4036_ _3565_ _3567_ _3571_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_37_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4246__I _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5987_ as2650.stack\[5\]\[6\] _1724_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7726_ _1844_ _2057_ _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4938_ _0377_ _0770_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7657_ _2314_ _3260_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6147__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ _3658_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4158__A1 _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6608_ as2650.stack\[4\]\[0\] _2272_ _2275_ as2650.stack\[6\]\[0\] _2276_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7588_ _1691_ _3022_ _3215_ _3056_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_105_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6539_ _1114_ _2182_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5805__I _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7647__A2 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6083__A1 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4633__A2 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7583__A1 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8006__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4397__A1 _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6371__I _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5897__A1 as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5715__I _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6974__C _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A1 _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__A2 _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7810__A2 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5910_ _1671_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6890_ _0577_ _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ _1541_ _3515_ _1563_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7574__A1 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6377__A2 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ _1570_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4927__A3 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7511_ _0386_ _3139_ _3067_ _3068_ _3109_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4723_ _0571_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7442_ _1418_ _3066_ _2984_ _3073_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7877__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4654_ _0506_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7373_ _3005_ _3006_ _1195_ _2304_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4585_ _3521_ _0395_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6324_ _0280_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6657__S _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6255_ _1526_ _1825_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5206_ _3681_ as2650.r123_2\[0\]\[5\] _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4312__A1 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6186_ _1869_ _1880_ _1882_ _1884_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5137_ _3608_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5068_ _3843_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5812__A1 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4019_ as2650.idx_ctrl\[0\] _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4091__A3 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7565__A1 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7709_ _1620_ _2992_ _2338_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7317__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4640__S _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4854__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6366__I _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6056__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7253__B1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7556__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4909__A3 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7308__A1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4790__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6531__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _3688_ _3903_ _3904_ _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7492__B1 _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6040_ as2650.stack\[3\]\[0\] _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7795__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7991_ _0110_ clknet_leaf_45_wb_clk_i as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6598__A2 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _2283_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4952__C _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5270__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6873_ as2650.stack\[1\]\[5\] _2402_ _2535_ as2650.stack\[0\]\[5\] _2536_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5824_ as2650.stack\[2\]\[9\] _1574_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5558__B1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5022__A2 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5755_ as2650.cycle\[3\] _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6879__C _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4781__A1 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4706_ _0514_ _0506_ _0555_ _0372_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5686_ _1447_ _1492_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7056__B _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7425_ _3017_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4637_ _3896_ _0483_ _0487_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6522__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7356_ _1921_ _2985_ _2989_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4568_ _0419_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6895__B _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6307_ _2000_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7078__A3 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7287_ _2885_ _2935_ _2936_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ as2650.holding_reg\[2\] _3503_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6286__A1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6238_ _1925_ _1935_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4836__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ _3770_ _1867_ _1868_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6589__A2 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7538__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4434__I _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6210__A1 _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7710__A1 _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4524__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4524__B2 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7413__C _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6029__A1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__A3 _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5004__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6201__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5376__S _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4763__A1 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _3509_ _1199_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5471_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7701__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ _0270_ _0276_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7210_ _2856_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7141_ _2795_ _2796_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4353_ _3853_ _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6268__A1 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7072_ _2430_ _2720_ _2729_ _1953_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4284_ _3760_ _3786_ _3761_ _3663_ _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_140_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6023_ _1599_ _1740_ _1751_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7768__A1 _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7974_ _0093_ clknet_leaf_39_wb_clk_i as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6925_ as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\] _3482_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6991__A2 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6856_ _2338_ _2467_ _2517_ _2519_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5807_ as2650.stack\[2\]\[6\] _1584_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6787_ as2650.stack\[1\]\[3\] _2451_ _2275_ as2650.stack\[2\]\[3\] _2452_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3999_ _3509_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5546__A3 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4754__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5738_ _1537_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ _1452_ _1464_ _1468_ _1475_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_136_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4506__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7408_ _3665_ _3730_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_102_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7339_ as2650.stack\[7\]\[10\] _2964_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4857__C _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6259__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6259__B2 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5857__I1 as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7759__A1 _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A1 _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_63 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_74 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_85 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4993__A1 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__A3 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6498__B2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5723__I _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4339__I _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5473__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6670__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5225__A2 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ as2650.r123\[1\]\[4\] _0815_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6710_ _2362_ _2374_ _2375_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4984__A1 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7690_ _1703_ _3022_ _3313_ _3056_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6641_ _2307_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6725__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6572_ _1908_ _2234_ _2236_ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5523_ _0311_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__S _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6489__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5454_ _1203_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4405_ _3810_ _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5161__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5385_ _3530_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5633__I _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4336_ _3864_ _3870_ _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7124_ as2650.stack\[5\]\[11\] _2340_ _2343_ as2650.stack\[6\]\[11\] _2781_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7055_ _2112_ _2710_ _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4267_ _3748_ _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6006_ _1739_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6661__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4198_ as2650.idx_ctrl\[0\] _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__I _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6413__A1 _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6413__B2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7957_ _0076_ clknet_leaf_38_wb_clk_i as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6964__A2 _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6908_ as2650.pc\[4\] net9 _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7888_ _0007_ clknet_leaf_58_wb_clk_i as2650.r123\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6839_ _2125_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6716__A2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5519__A3 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4712__I as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7228__C _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6639__I _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5543__I _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4159__I _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6652__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3998__I _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6374__I _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4966__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5718__I _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__A1 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7154__B _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5143__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5694__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5170_ _0987_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4121_ _3655_ _3656_ _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4052_ as2650.cycle\[4\] _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_77_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7199__A2 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5121__C _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7811_ _1414_ _2015_ _2221_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6946__A2 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8062__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7742_ _0299_ _3356_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7673_ _2586_ _3296_ _2731_ _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4885_ _3829_ _0730_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4532__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6624_ _2269_ _2291_ _2126_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7048__C _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7371__A2 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5382__A1 as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6555_ _1887_ _1804_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5506_ _0662_ _0560_ _0492_ _0407_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6486_ _1885_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5437_ _1244_ _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6882__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5685__A2 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5368_ _0874_ _1182_ _1184_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7107_ as2650.pc\[10\] _0669_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4319_ _3853_ _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8087_ _0206_ clknet_3_0_0_wb_clk_i as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5299_ _1066_ _1067_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6634__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5437__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7831__B1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7511__C _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7038_ _2248_ _2690_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_47_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4707__I _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7362__A2 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__A2 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6873__A1 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8085__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6928__A2 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7050__A1 as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4939__A1 _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4939__B2 _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4670_ as2650.r123\[2\]\[4\] _0433_ _0522_ _3634_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7922__CLK clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5364__A1 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6340_ _1843_ _1307_ _2029_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7105__A2 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6271_ _1783_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6864__A1 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8010_ _0129_ clknet_leaf_33_wb_clk_i as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5222_ _1009_ _1049_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5667__A2 _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4714__I1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _0947_ _0949_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5911__I _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4104_ _3489_ _3639_ _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5084_ _0284_ _0848_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6092__A2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4035_ _3506_ _3570_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6742__I _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _1595_ _1717_ _1728_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4690__C _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6395__A3 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7725_ _1921_ _3341_ _3346_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4937_ _3645_ _3716_ _3851_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ net37 _3280_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4868_ _0717_ _3660_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4158__A2 _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6607_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7587_ _2575_ _3195_ _3214_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ _0620_ _0621_ _0648_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6538_ _2185_ _2207_ _2208_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6469_ _3587_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5658__A2 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6917__I _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8139_ _0258_ clknet_leaf_22_wb_clk_i as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6083__A2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4094__A1 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7945__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4397__A2 _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5594__A1 _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4172__I _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7483__I _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6099__I _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7271__A1 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4347__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7023__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5840_ _1627_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6377__A3 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ as2650.pc\[1\] _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4082__I _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7510_ _0387_ _3139_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _0573_ _0554_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7607__B _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8100__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7441_ _3067_ _3070_ _3072_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4653_ _0499_ _3617_ _0502_ _3522_ _0505_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_124_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__I _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7372_ _3846_ _1968_ _1898_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4584_ _0391_ _3616_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5127__B _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6323_ _1383_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4560__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6837__A1 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ _1936_ _1950_ _1951_ _1280_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5205_ _0999_ _1003_ _1001_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4312__A2 _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6185_ _1883_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5641__I _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _3604_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7262__A1 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5067_ _0861_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4076__A1 _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7968__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5812__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4018_ as2650.idx_ctrl\[1\] _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7014__A1 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7565__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5576__A1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _1716_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7708_ _1620_ _1322_ _2479_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7639_ _3219_ _3220_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5816__I _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4000__A1 _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4551__A2 _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7253__A1 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7005__A1 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7556__A2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8123__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5567__A1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A2 _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5726__I _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6819__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7492__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5461__I _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7990_ _0109_ clknet_leaf_40_wb_clk_i as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7795__A2 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6941_ _2286_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5270__A3 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6872_ _1713_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5823_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5558__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5558__B2 _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5754_ _1244_ _1351_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4230__A1 _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4705_ _0275_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4781__A2 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5685_ _1257_ _1451_ _1491_ _1439_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7424_ _1572_ _3022_ _3055_ _3056_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7056__C _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4636_ _0488_ _0401_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7355_ _2137_ _2254_ _2987_ _2988_ _2832_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4567_ _0327_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ _1266_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7286_ _1017_ _2862_ _2751_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _3502_ _3930_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6237_ _1528_ _1926_ _1934_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_131_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6168_ net22 _1867_ _1431_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7235__A1 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _0384_ _0848_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ _1788_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7786__A2 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7538__A2 _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5549__A1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4450__I _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4524__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4288__A1 _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6029__A2 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7226__A1 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A1 as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6326__B _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6201__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5456__I _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ _3519_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _0272_ _3873_ _0274_ _0275_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_126_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5712__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8019__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7140_ as2650.pc\[12\] _1097_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4352_ _3875_ _3881_ _3885_ _3886_ _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7465__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6268__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7465__B2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7071_ _1520_ _2725_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4283_ _3812_ _3817_ _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6022_ as2650.stack\[0\]\[6\] _1746_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7217__A1 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7973_ _0092_ clknet_leaf_39_wb_clk_i as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6924_ _2384_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6855_ _2518_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5806_ _1599_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4203__A1 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6786_ _1546_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3998_ _3533_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5737_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4754__A2 _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5366__I _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5668_ _1469_ _1470_ _1474_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7407_ _0314_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4619_ _0470_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4506__A2 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5703__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5599_ _1406_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7338_ _1732_ _2962_ _2975_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7456__A1 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7269_ _2914_ _0494_ _2162_ _0561_ _2919_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_133_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7530__B _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7208__B2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7759__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_53 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_64 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4442__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_75 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_86 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6660__I _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4180__I _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7695__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_1_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6498__A2 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7440__B _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6670__A2 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4681__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__A2 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4355__I _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4970_ _0808_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4984__A2 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _1930_ _1933_ _1815_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6571_ _1779_ _1226_ _2237_ _2238_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_121_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5522_ _1328_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_117_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ _1225_ _1227_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4404_ _3916_ _3918_ _3936_ _3937_ _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5384_ as2650.psu\[5\] _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7123_ _2679_ _2778_ _2779_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4335_ _3521_ _3869_ _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7054_ _2444_ _2711_ _2712_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4266_ _3518_ _3801_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6005_ _1739_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6661__A2 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _3723_ _3732_ _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7610__A1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7956_ _0075_ clknet_leaf_40_wb_clk_i as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6907_ _2568_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7887_ _0006_ clknet_leaf_58_wb_clk_i as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _2479_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6177__A1 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5519__A4 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6769_ _2331_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5152__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8059__D _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4175__I as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7601__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4966__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6390__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5391__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7668__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7668__B2 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5679__B1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6340__A1 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4120_ _3650_ as2650.r123_2\[1\]\[7\] _3495_ _3551_ _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4051_ as2650.cycle\[5\] _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput5 io_in[5] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7053__C1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4085__I _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7810_ _1154_ _3402_ _1374_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4406__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _0335_ _3354_ _3359_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4953_ _3523_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4813__I _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7672_ net38 _3295_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6159__A1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4884_ _0731_ _0732_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6623_ _1672_ _1264_ _2290_ _2116_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5906__A1 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6554_ _1246_ _1216_ _1356_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_119_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7659__A1 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5505_ _0280_ _3842_ _3715_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6485_ _1920_ _2153_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _3752_ _3499_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6882__A2 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5367_ as2650.r123_2\[1\]\[0\] _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7106_ as2650.pc\[11\] _2589_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4318_ _3620_ _3598_ _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8086_ _0205_ clknet_leaf_3_wb_clk_i as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5298_ _1066_ _1067_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7080__B _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6634__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7037_ _2362_ _2695_ _2375_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7831__A1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4249_ _3762_ _3785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7831__B2 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6398__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7939_ _0058_ clknet_leaf_30_wb_clk_i as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5070__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6570__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4879__B _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5554__I _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5125__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6873__A2 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5920__I1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4884__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6385__I _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7822__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4636__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7050__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4939__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5061__A1 _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5464__I _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6313__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6270_ _1446_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ _1029_ _1048_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6864__A2 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4714__I2 as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5152_ _0947_ _0949_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6295__I _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4103_ _3593_ _3596_ _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5413__B _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7813__A1 _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ _0869_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4034_ _3569_ _3557_ _3540_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_65_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7041__A2 _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5985_ as2650.stack\[5\]\[5\] _1724_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7724_ _2167_ _3338_ _3344_ _3051_ _3345_ _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_40_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6395__A4 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4936_ _3854_ _0775_ _0785_ _3890_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7655_ net50 _3265_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ as2650.holding_reg\[7\] _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6606_ _2273_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7586_ _3085_ _3197_ _3213_ _2833_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6552__A1 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ _0620_ _0621_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6537_ net20 _2178_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7897__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4563__B1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6304__A1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6468_ _2145_ _2146_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5419_ _0802_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6399_ _2067_ _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8138_ _0257_ clknet_leaf_13_wb_clk_i as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6419__B _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4718__I _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8069_ _0188_ clknet_leaf_12_wb_clk_i as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6083__A3 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8072__D _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5594__A2 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7343__I0 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8052__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5282__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6843__I _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_1_0_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _1539_ _1567_ _1569_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A2 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _3498_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7440_ _3067_ _3070_ _3071_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4652_ _0503_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7607__C _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7371_ _1791_ _1827_ _1906_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4583_ _3815_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6322_ _2014_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6837__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6253_ net26 _1936_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5922__I _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5204_ _1033_ _1039_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6184_ _3513_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__I _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5135_ _0445_ _0462_ _0338_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7262__A2 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5066_ _3842_ _3714_ _0867_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_57_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5273__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4076__A2 _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4017_ _3552_ _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7014__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ _1715_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5576__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7707_ _3184_ _3329_ _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4919_ _0400_ _0482_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5899_ as2650.stack\[4\]\[7\] _1660_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7638_ _2887_ _3255_ _3263_ _2984_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5318__B _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7569_ _2569_ _3196_ _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5832__I _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5887__I0 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7252__C _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4448__I _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7912__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7253__A2 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5264__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__B1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7005__A2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5016__A1 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5279__I _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__I _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5567__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6764__A1 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7494__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6819__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7492__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6940_ as2650.stack\[0\]\[6\] _2508_ _2601_ as2650.stack\[2\]\[6\] _2602_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _2533_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5007__A1 _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5822_ _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5558__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5753_ _1550_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8098__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4704_ _0528_ _0485_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6507__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5684_ _1257_ _1476_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7704__B1 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7423_ _1990_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4635_ _3729_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7180__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7354_ net28 _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4566_ _0295_ as2650.r123\[0\]\[1\] _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_25_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6305_ _0698_ _1311_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7285_ _0663_ _1364_ _2926_ _2934_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_143_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4497_ _0346_ _0349_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7072__C _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7935__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6236_ _1930_ _1933_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4541__I0 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6167_ _1440_ _3570_ _1866_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5118_ _0920_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7235__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6098_ _1328_ _1806_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7786__A3 _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6483__I _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5049_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6994__A1 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5099__I _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6746__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5549__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__B2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3980__A1 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__I _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7226__A2 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6393__I _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4748__B1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6201__A3 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5737__I _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7162__A1 as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ _0271_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7958__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4351_ _3856_ _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7465__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7070_ _2247_ _2727_ _2126_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4282_ as2650.holding_reg\[1\] _3816_ _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4279__A2 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ _1594_ _1740_ _1750_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4088__I _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7217__A2 _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7399__I _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6976__A1 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7972_ _0091_ clknet_leaf_41_wb_clk_i as2650.stack\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6923_ _2250_ _2578_ _2582_ _2584_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6728__A1 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6854_ _2113_ _2467_ _1243_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout49 net13 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5805_ _1598_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6785_ _2444_ _2446_ _2449_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5647__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3997_ _3532_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5736_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5667_ _0894_ _3707_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7153__B2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7406_ _1415_ _3032_ _3034_ _3038_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4618_ _0415_ _0469_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5703__A2 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5598_ _0781_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7337_ as2650.stack\[7\]\[9\] _2964_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4549_ _3641_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7268_ _1423_ _1941_ _2918_ _1939_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8113__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5467__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6219_ _3496_ _3489_ _3535_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7199_ _3553_ _3610_ _2852_ _1318_ _2853_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7208__A2 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4726__I _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__A1 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__B2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A3 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_54 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_65 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_76 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6941__I _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_87 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7392__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5557__I _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6162__B _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6195__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4681__A2 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A1 _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4984__A3 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7168__B _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6186__A2 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4197__A1 _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6570_ _1351_ _1982_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5521_ _3673_ _3548_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5452_ _3510_ _1231_ _1233_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8136__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ _3793_ _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5383_ _1156_ _1182_ _1192_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7122_ as2650.stack\[1\]\[11\] _2340_ _2278_ as2650.stack\[3\]\[11\] _2779_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4334_ _3866_ _3868_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _3478_ _3614_
+ _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_113_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5449__A1 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ as2650.stack\[7\]\[9\] _2283_ _2284_ as2650.stack\[6\]\[9\] _1713_ as2650.stack\[4\]\[9\]
+ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_119_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4265_ as2650.r123\[2\]\[0\] _3636_ _3799_ _3800_ _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6004_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4196_ _3719_ _3731_ _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6949__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7955_ _0074_ clknet_leaf_40_wb_clk_i as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6906_ as2650.pc\[6\] _0668_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7886_ _0005_ clknet_leaf_58_wb_clk_i as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _2090_ _2487_ _2496_ _2500_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7374__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4281__I _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6768_ _2308_ _2426_ _2429_ _1873_ _2432_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5719_ _1522_ _1515_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7126__A1 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7592__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6710__B _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6699_ _1942_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5688__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4230__B as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6157__B _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5860__A1 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4456__I _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7601__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__A2 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6671__I _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8009__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7365__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6168__A2 _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5391__A3 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7668__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6876__B1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5679__B2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6340__A2 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6846__I _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4103__A1 _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4050_ as2650.cycle\[7\] _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7840__A2 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 io_in[6] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7053__B1 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7053__C2 as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4406__A2 _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5603__A1 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7740_ _3866_ _3356_ _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4952_ _3693_ _0800_ _3748_ _3841_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7671_ net37 net50 _3265_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7356__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4883_ _0721_ _0732_ _3821_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6159__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _2280_ _2289_ _1204_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5906__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6553_ _3543_ _1355_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5925__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5504_ _1101_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6484_ _2161_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5146__B _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5435_ _3573_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4342__A1 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _1181_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4985__B _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7105_ _2247_ _2755_ _2757_ _2251_ _2761_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4317_ _3691_ _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8085_ _0204_ clknet_leaf_62_wb_clk_i as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5297_ _1085_ _1086_ _1083_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6095__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7036_ _2422_ _2694_ _2690_ _2364_ _2474_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_59_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4248_ _3783_ _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7831__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5842__A1 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4179_ _3714_ _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7044__B1 _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7595__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6398__A2 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7938_ _0057_ clknet_leaf_37_wb_clk_i as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7347__A1 _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7869_ _1419_ _2011_ _3455_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6570__A2 _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5056__B _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6666__I _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7271__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7822__A2 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4636__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7586__A1 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7338__A1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6561__A2 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7165__C _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7510__A1 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6313__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5220_ _0711_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4714__I3 as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ _3712_ _0945_ _0950_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4102_ _3538_ _3552_ _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5082_ _0906_ _0919_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7813__A2 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4096__I _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _3568_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_84_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _1727_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7723_ _1870_ _2868_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7329__A1 as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4935_ _3857_ _0776_ _0784_ _3888_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7654_ _3277_ _3278_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ _0716_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6605_ _1542_ _1710_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7585_ _2986_ _3192_ _3212_ _3116_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4797_ _0644_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6552__A2 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4563__A1 _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4563__B2 _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6536_ _2187_ _0706_ _2206_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6467_ _2145_ _2146_ _2147_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7501__A1 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6304__A2 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4315__A1 _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5418_ _1158_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6398_ _2068_ _1906_ _2081_ _2082_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5349_ _1173_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8137_ _0256_ clknet_leaf_12_wb_clk_i as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5390__I _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6419__C _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7804__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8068_ _0187_ clknet_leaf_15_wb_clk_i net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ _2281_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7017__B1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5594__A3 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7266__B _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5565__I _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7740__A1 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4554__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4402__C _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7343__I1 as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7991__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4857__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7559__A1 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7559__B2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6231__A1 _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _3807_ _3626_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7176__B _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4651_ _3649_ as2650.r123_2\[1\]\[5\] _3494_ _3551_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__6534__A2 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7731__B2 _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4545__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4582_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7370_ _3003_ _1930_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6321_ _2013_ _3803_ _2005_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6298__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6252_ _1937_ _1949_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5203_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6183_ _1881_ _1880_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5134_ _0968_ _0971_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7798__A1 _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _3702_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6470__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4016_ _3551_ _3533_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_84_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _1628_ _1714_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7706_ _2825_ _3318_ _2771_ _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4918_ _0528_ _0568_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5898_ _1600_ _1654_ _1665_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7637_ _3260_ _3262_ _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5385__I _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4849_ _0684_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7568_ _2525_ _3179_ _2572_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _2182_ _0960_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7499_ _2416_ _3119_ _3128_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6289__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7789__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5264__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6461__A1 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8083__D _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6213__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6764__A2 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4775__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4413__B _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7713__A1 _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4527__A1 _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4639__I _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7244__A3 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7887__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4374__I _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6870_ _2362_ _2531_ _2532_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6204__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ as2650.pc\[9\] _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5752_ _3594_ _1499_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4703_ _0529_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ _1467_ _1489_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7704__B2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7422_ _1374_ _3030_ _3050_ _3054_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4634_ _0485_ _0486_ _3895_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7180__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7353_ _2986_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4565_ _0296_ _3743_ _3837_ _3861_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5191__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5933__I _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6304_ _1900_ _1901_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4496_ _0346_ _0349_ _3919_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7284_ _2409_ _0576_ _2933_ _1374_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4549__I _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6235_ _1931_ _1932_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4541__I1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6166_ _3512_ _1235_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_97_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _0951_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6097_ _1802_ _1805_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ _3855_ _0834_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7809__B _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6999_ _1607_ _2658_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8042__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3980__A2 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7544__B _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6939__I _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5182__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5843__I _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5064__B _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4459__I _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6682__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6434__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4408__B _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4996__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6737__A2 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4748__B2 _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5173__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4350_ _3883_ _3884_ _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4281_ _3811_ _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ as2650.stack\[0\]\[5\] _1746_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6584__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7971_ _0090_ clknet_leaf_40_wb_clk_i as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8065__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6922_ _1424_ _2583_ _1853_ _3605_ _2032_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_70_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6853_ _2505_ _2512_ _2516_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6728__A2 _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5928__I _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5804_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6784_ as2650.stack\[4\]\[3\] _2447_ _2448_ as2650.stack\[6\]\[3\] _2449_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3996_ _3531_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_5735_ as2650.pc\[0\] _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5666_ _1472_ _0306_ _1452_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7153__A2 _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7405_ _3035_ _3036_ _3037_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5164__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4617_ _0415_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6900__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5597_ _1375_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7336_ _2974_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4548_ _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7267_ _1379_ _1096_ _2916_ _2917_ _1409_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _0267_ _0324_ _0332_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6664__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5467__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6218_ _1332_ _1914_ _1915_ _1360_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7198_ _3537_ _3562_ _1896_ _1797_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_131_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6708__B _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6149_ _1525_ _1850_ _1831_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7759__A4 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_55 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_66 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_77 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_88 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5838__I _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7392__A2 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6195__A3 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__A2 _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7274__B _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6655__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6407__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4418__B1 _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5949__S _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7080__A1 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5630__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7449__B _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _1309_ _1323_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5146__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5451_ _1243_ _1247_ _1254_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4402_ _3919_ _3925_ _3933_ _3935_ _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5941__I0 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5382_ as2650.r123_2\[1\]\[7\] _1183_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7121_ as2650.stack\[0\]\[11\] _2272_ _2343_ as2650.stack\[2\]\[11\] _2778_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4333_ _3867_ _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5449__A2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7052_ as2650.stack\[5\]\[9\] _2340_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4264_ _3634_ _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _1541_ _1564_ _1651_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4195_ _3730_ _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7203__I _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7954_ _0073_ clknet_leaf_38_wb_clk_i as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6905_ _2566_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7359__B _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7885_ _0004_ clknet_leaf_57_wb_clk_i as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6836_ _2498_ _2499_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6177__A3 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _2430_ _2421_ _2431_ _2381_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3979_ _3514_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5718_ _1362_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6698_ _2363_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7094__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ _1455_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4230__C as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7319_ _1679_ as2650.stack\[7\]\[1\] _2964_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5860__A2 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output43_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7948__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__A3 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5568__I _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7365__A2 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7117__A2 _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5128__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5679__A2 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6876__B2 as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6628__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput7 io_in[7] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4951_ _3584_ _3610_ _0799_ _3613_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_91_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7670_ _3018_ _3293_ _3294_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4882_ _0700_ _0570_ _0688_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7356__A2 _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6621_ _2282_ _2285_ _2288_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7693__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6552_ _1481_ _2086_ _2215_ _2220_ _2131_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5119__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5503_ _1310_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6483_ _1995_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__I _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5434_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7642__B _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__A2 _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5365_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7104_ _2434_ _2759_ _2760_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4316_ _3850_ _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8084_ _0203_ clknet_leaf_3_wb_clk_i as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5296_ _1128_ _1129_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6258__B _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6095__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7292__A1 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ _2691_ _2693_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4247_ _3757_ _3758_ _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5842__A2 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ _3713_ _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__A1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7044__B2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7595__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6398__A3 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7937_ _0056_ clknet_leaf_9_wb_clk_i as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5388__I _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__B1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7868_ _2899_ _3467_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4225__C _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6819_ _2365_ _2466_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6721__B _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7799_ _1284_ _3832_ _3405_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6168__B _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8086__D _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7283__A1 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7035__A1 _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7586__A2 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8126__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7338__A2 _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6149__I0 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7510__A2 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5521__A1 _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5150_ _0952_ _0953_ _0951_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4101_ _3631_ _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7274__A1 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ _0906_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6321__I0 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5824__A2 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4032_ as2650.ins_reg\[2\] _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7026__A1 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7577__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5588__A1 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5983_ _1589_ as2650.stack\[5\]\[4\] _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7722_ _2796_ _3343_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4934_ _3875_ _0780_ _0783_ _3856_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_19_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7329__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7653_ _1608_ _1387_ _3246_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4865_ _0524_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_60_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4840__I _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6604_ _1712_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _3204_ _3211_ _2167_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4012__A1 _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4796_ _0597_ _0645_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6535_ _1380_ _2182_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4563__A2 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5760__A1 _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6466_ _2145_ _2146_ _1431_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7501__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4315__A2 _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _1194_ _1199_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5671__I _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6397_ _1323_ _1465_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8136_ _0255_ clknet_3_2_0_wb_clk_i net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5348_ as2650.r123\[3\]\[0\] _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7265__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8067_ _0186_ clknet_leaf_15_wb_clk_i net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4079__A1 _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5279_ _3645_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7018_ _2444_ _2676_ _2677_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6716__B _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5594__A4 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4003__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7740__A2 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4554__A2 _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5751__A1 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5782__S _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7008__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__I _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4490__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7559__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6231__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A1 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5990__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4650_ _0396_ as2650.r123\[1\]\[5\] _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7731__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 wb_rst_i net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4581_ _3754_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6320_ _1460_ _1307_ _2012_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7495__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7192__B _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6251_ _1440_ _1939_ _1857_ _1947_ _1948_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5202_ _1034_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6182_ _3525_ _3526_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5133_ as2650.r123_2\[2\]\[3\] _0969_ _0970_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _3908_ _0903_ _0869_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4015_ _3550_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7211__I _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6758__B1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5966_ _1713_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7705_ _2869_ _3327_ _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4917_ _0752_ _0753_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5981__A1 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ as2650.stack\[4\]\[6\] _1660_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7636_ _2253_ _3261_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ _0653_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7567_ _1691_ _3024_ _3184_ _3194_ _1319_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5733__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _0390_ _3865_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5733__B2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _2179_ _2191_ _2193_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7814__C _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7498_ as2650.pc\[3\] _0386_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7486__A1 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _2086_ _3546_ _2128_ _2130_ _2131_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_106_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7238__A1 _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8119_ _0238_ clknet_leaf_61_wb_clk_i as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6446__B _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6461__A2 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4472__A1 _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__A2 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5972__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4527__A2 _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7724__C _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7477__A1 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6524__I0 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7229__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6452__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6204__A2 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5820_ _1611_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4215__A1 _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ _3524_ _1466_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4766__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _0400_ _0482_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5682_ as2650.psu\[0\] _1453_ _1480_ as2650.psu\[4\] _1488_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__7165__B1 _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7704__A2 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7421_ _3051_ _3053_ _2833_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4633_ _0370_ _0304_ _0439_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7352_ _1919_ _1794_ _1239_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4564_ _0416_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7468__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6303_ _1365_ _0799_ _1995_ _1996_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7283_ _1271_ _1375_ _2930_ _2932_ _2409_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_116_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4495_ _3917_ _0347_ _0348_ _3813_ _3923_ _0261_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_4
XFILLER_143_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6234_ _0831_ _3779_ _1220_ _1221_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_143_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6140__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7650__B _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _1241_ _1252_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4541__I2 as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5116_ _0952_ _0953_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _1329_ _1803_ _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7640__A1 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5047_ _3874_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_34_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6998_ _1602_ _2563_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7981__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5949_ as2650.stack\[1\]\[9\] _1700_ _1697_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5396__I _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7619_ _2617_ _2652_ _3244_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3980__A3 _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5182__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7459__A1 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6131__A1 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7560__B _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5485__A3 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6434__A2 _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6623__C _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7698__A1 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6370__A1 _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4920__A2 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ _3814_ _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7470__B _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7870__A1 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7622__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7970_ _0089_ clknet_leaf_38_wb_clk_i as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4436__A1 _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _2385_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _2513_ _2514_ _2515_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6189__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5803_ as2650.pc\[6\] _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6783_ _2274_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4739__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3995_ as2650.ins_reg\[1\] _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ _1534_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7689__A1 _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5665_ _1471_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5944__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7404_ _3035_ _3036_ _2981_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4616_ _3681_ _0393_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5164__A2 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5596_ _1379_ _1397_ _1399_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5703__A4 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7335_ _1696_ as2650.stack\[7\]\[8\] _2969_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4547_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7266_ _0707_ _2197_ _2052_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4478_ _3748_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6217_ _1308_ _3600_ _1799_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6664__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7861__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7197_ _1808_ _2851_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4675__A1 _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6708__C _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ _3846_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6416__A2 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6079_ _1787_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_56 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_67 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_78 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7539__C _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_89 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_53_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__A3 _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8089__D _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6104__A1 _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6655__A2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7604__A1 _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6407__A2 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4418__B2 _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__A1 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5450_ _1255_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4401_ _3934_ _3788_ _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5381_ _1191_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5941__I1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7120_ _2246_ _2762_ _2774_ _2090_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_99_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4332_ as2650.r123_2\[0\]\[2\] _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7051_ _2679_ _2708_ _2709_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4263_ _3798_ _3799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6002_ _1737_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4194_ _3724_ _3729_ _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4409__A1 _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7071__A2 _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7953_ _0072_ clknet_leaf_30_wb_clk_i as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5939__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ _2563_ _2565_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7884_ _0003_ clknet_leaf_60_wb_clk_i as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6835_ _1479_ _1817_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6177__A4 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6766_ _2365_ _2415_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3978_ _3512_ _3513_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5717_ _1520_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7375__B _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6697_ _2000_ _1505_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5674__I as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5648_ _1454_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6334__A1 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _1098_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4896__A1 _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7318_ _2959_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_78_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7834__A1 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _2887_ _0376_ _2900_ _1970_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7269__C _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6573__A1 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7285__B _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5128__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6325__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6876__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8055__CLK clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7825__A1 _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 io_in[8] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7053__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5064__A1 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _3629_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7179__C _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4881_ _0721_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6620_ as2650.stack\[1\]\[0\] _2286_ _2287_ as2650.stack\[0\]\[0\] _2288_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6564__A1 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _1529_ _2219_ _1861_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5502_ _3934_ _1309_ _3574_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6482_ _1885_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6316__A1 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5119__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6867__A2 _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5433_ _1237_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5364_ _0820_ _0826_ _0943_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7103_ as2650.addr_buff\[3\] _2663_ _2736_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4315_ _3621_ _3847_ _3849_ _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8083_ _0202_ clknet_leaf_5_wb_clk_i as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _3836_ as2650.r123_2\[0\]\[6\] _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7214__I _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ _2692_ _2655_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4246_ _3752_ _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4177_ _3712_ _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5055__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__A4 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7936_ _0055_ clknet_leaf_9_wb_clk_i as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4802__B2 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7867_ as2650.psu\[3\] _3465_ _3466_ _3461_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6818_ as2650.addr_buff\[4\] _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6555__A1 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6721__C _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7798_ _3805_ _3831_ _3404_ _3795_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ _1576_ as2650.pc\[1\] _1535_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6858__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7807__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7283__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5294__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5579__I _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6546__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6149__I1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4309__B1 _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__A2 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4100_ _3635_ _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ _0917_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7274__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6321__I1 _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5285__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4031_ as2650.ins_reg\[3\] _3566_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7026__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5037__A1 as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6785__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _1716_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_65_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5588__A2 _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7721_ _2794_ _3342_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4933_ _0782_ _3884_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6537__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7652_ _1699_ _0670_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4864_ _0525_ _0713_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6603_ _2270_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7583_ _1456_ _3066_ _1802_ _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ _0595_ _0610_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_59_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4012__A2 _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6534_ _2185_ _2204_ _2205_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5760__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7653__B _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ _1248_ _2133_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7938__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5416_ _1202_ _1213_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6396_ _2070_ _2073_ _2080_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8135_ _0254_ clknet_leaf_12_wb_clk_i as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5347_ _1172_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8066_ _0185_ clknet_leaf_18_wb_clk_i net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7265__A2 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5278_ _1111_ _1112_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4079__A2 _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7017_ as2650.stack\[5\]\[8\] _2277_ _2447_ as2650.stack\[4\]\[8\] _2677_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4229_ _3764_ _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6716__C _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7017__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6776__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7919_ _0038_ clknet_3_4_0_wb_clk_i as2650.r123\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6528__A1 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5200__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4003__A2 _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5751__A2 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6700__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4478__I _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7256__A2 _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5267__A1 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6693__I _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6626__C _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7008__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6067__I0 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6767__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5102__I _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5990__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7192__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _3635_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7319__I0 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5772__I _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6250_ net26 _1900_ _1273_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7495__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5201_ _1000_ _1035_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_131_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6181_ _1871_ _1874_ _1879_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5132_ _0876_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _0855_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4014_ as2650.ins_reg\[0\] _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__6108__I _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6758__B2 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5965_ _1712_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4233__A2 _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7704_ _3319_ _3324_ _3326_ _3085_ _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4916_ _0754_ _0759_ _0765_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_40_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5896_ _1595_ _1654_ _1664_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5981__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7635_ _3257_ _3259_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4847_ _0539_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7183__A1 as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7566_ _2586_ _3192_ _3193_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4778_ _0627_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6517_ net42 _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7497_ _2468_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7486__A2 _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6448_ _1279_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8116__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5497__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6379_ _2061_ _2063_ _1553_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8118_ _0237_ clknet_leaf_60_wb_clk_i as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7238__A2 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6727__B _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8049_ _0168_ clknet_leaf_10_wb_clk_i as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6997__A1 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5421__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5972__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7174__A1 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__A3 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7293__B _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7477__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_4_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6524__I1 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4160__A1 _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7229__A2 _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6988__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5767__I _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4215__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5412__A1 as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _1205_ _3594_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A1 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4701_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5681_ _1481_ _1406_ _0286_ _1482_ _1487_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_124_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7165__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7165__B2 _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7420_ _3052_ _2302_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4632_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7351_ _2870_ _2980_ _2983_ _2984_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4923__B1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4563_ _3834_ _3866_ _0299_ _3712_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4923__C2 _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6302_ _0698_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7282_ _1375_ _2931_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4494_ _3870_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5479__B2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6233_ _1197_ _1222_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6140__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4151__A1 _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6164_ _1862_ _1863_ _1864_ _1280_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_135_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4541__I3 as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6428__B1 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5115_ _0279_ _0866_ _0917_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6095_ _1558_ _1787_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6979__A1 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7222__I _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4454__A2 _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5677__I as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6997_ _2655_ _2656_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5403__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4581__I _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5948_ _1699_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7618_ _2651_ _3196_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6903__A1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7549_ _3031_ _3162_ _3177_ _3049_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6301__I _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7459__A2 _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4142__A1 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6457__B _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5890__A1 as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7395__A1 _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__I _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4491__I _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7147__A1 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6370__A2 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4381__A1 _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7870__A2 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5271__B _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7083__B1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7622__A2 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4436__A2 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6920_ _1521_ _2574_ _2580_ _2581_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ as2650.stack\[7\]\[4\] _2507_ _2508_ as2650.stack\[4\]\[4\] _2515_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7386__A1 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6189__A2 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _1595_ _1567_ _1596_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_opt_1_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3994_ _3529_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6782_ _1712_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7138__A1 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ _1376_ _1515_ _1523_ _1525_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5664_ net8 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7403_ _1458_ _3893_ _3905_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_4615_ _0466_ _0467_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5595_ _1400_ _1401_ _1402_ _0768_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_102_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7334_ _1603_ _2962_ _2973_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4546_ _0392_ _3617_ _0395_ _3522_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_117_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7661__B _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4477_ _3746_ _0331_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7265_ as2650.psu\[4\] _2836_ _2915_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6216_ _1913_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7196_ _3607_ _0973_ _1310_ _1901_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7861__A2 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4675__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _1848_ _1834_ _1849_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6078_ _3545_ _1557_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6416__A3 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5624__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6791__I _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5029_ _0865_ _0867_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_57 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_68 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_79 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7129__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__A4 _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6104__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7301__A1 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4115__A1 _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7852__A2 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5863__A1 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5091__B _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5091__A2 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7540__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4400_ _3808_ _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5380_ _1110_ as2650.r123_2\[1\]\[6\] _1187_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ _3865_ _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5780__I _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7050_ as2650.stack\[1\]\[9\] _2451_ _2448_ as2650.stack\[2\]\[9\] _2709_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7971__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4262_ _3750_ _3797_ _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5854__A1 as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4657__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ _1626_ as2650.stack\[5\]\[12\] _1726_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4396__I _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4193_ _3726_ _3728_ _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7952_ _0071_ clknet_leaf_30_wb_clk_i as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6903_ _1598_ _2564_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7359__A1 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7883_ _0002_ clknet_leaf_61_wb_clk_i as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _2497_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6765_ _2309_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3977_ net10 _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5955__I _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5716_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4593__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7375__C _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6696_ _2247_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5647_ net2 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7531__A1 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6334__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__A1 _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5578_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4896__A2 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7317_ _1709_ _2961_ _2963_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6786__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4529_ _0381_ _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6098__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7248_ _2887_ _0380_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7834__A2 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7179_ _2825_ _3796_ _2829_ _2831_ _2833_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_58_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__B _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7770__A1 as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6573__A2 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4584__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__C _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5086__B _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6325__A2 _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__A1 _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7994__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6696__I _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7825__A2 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5105__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput9 io_in[9] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5064__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5976__S _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4880_ _0691_ _0726_ _0729_ _0453_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7476__B _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6564__A2 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__A1 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4575__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6550_ _2212_ _1353_ _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5501_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7513__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6481_ _1430_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6316__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4327__A1 _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5432_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4878__A2 _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5363_ _1180_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _2758_ _2737_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _3848_ _3603_ _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5294_ _0392_ _0945_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8082_ _0201_ clknet_leaf_30_wb_clk_i as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7033_ _1607_ _1098_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4245_ _3662_ _3764_ _3780_ _3781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ _3711_ _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__A3 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6252__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7935_ _0054_ clknet_3_3_0_wb_clk_i as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A2 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7866_ _3458_ _2024_ _2021_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _1587_ _2480_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7752__A1 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7797_ _0698_ _3852_ _3762_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6555__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4566__A1 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6748_ _2358_ _2413_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5763__B1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6679_ _2281_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4318__A1 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6449__C _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7807__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7341__S _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6491__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7743__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8022__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4004__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4309__A1 _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4309__B2 _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7315__I _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6482__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4030_ as2650.ins_reg\[4\] _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6234__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__C _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5981_ _1723_ _1717_ _1725_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5588__A3 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7720_ _2765_ _2763_ _3308_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7651_ _3020_ _3275_ _3276_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4863_ as2650.r123\[2\]\[6\] _0433_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7734__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6602_ as2650.stack_ptr\[2\] _1649_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7582_ _2981_ _3209_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4794_ _0595_ _0610_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ net19 _2192_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _3588_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5415_ _1214_ _1218_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6395_ _1439_ _2074_ _2076_ _2079_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_28_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8134_ _0253_ clknet_leaf_22_wb_clk_i as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5346_ _1171_ as2650.r123_2\[0\]\[7\] _1161_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8065_ _0184_ clknet_leaf_15_wb_clk_i net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5277_ as2650.r123_2\[2\]\[6\] _0969_ _0970_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6473__A1 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5276__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7016_ as2650.stack\[7\]\[8\] _2278_ _2275_ as2650.stack\[6\]\[8\] _2676_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4323__I1 as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4228_ _3761_ _3763_ _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4159_ _3694_ _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6225__A1 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7918_ _0037_ clknet_3_4_0_wb_clk_i as2650.r123\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7849_ _0803_ _1208_ _1877_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7725__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7844__B _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5751__A3 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5339__I0 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5364__B _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7135__I _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6700__A2 _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4711__A1 _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4494__I _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7413__B1 _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6067__I1 as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__A2 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7716__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7192__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4669__I _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5200_ as2650.r0\[4\] as2650.r123_2\[0\]\[1\] _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4702__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _1254_ _1876_ _1878_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _0827_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5062_ _0879_ _0900_ _0901_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ _3503_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5663__C1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8068__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6758__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ as2650.stack_ptr\[1\] _1711_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6552__C _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7703_ _2763_ _3325_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4915_ _0762_ _0763_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5895_ as2650.stack\[4\]\[5\] _1660_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6124__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7634_ as2650.addr_buff\[0\] _3257_ _3259_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4846_ _0692_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7183__A2 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7565_ _1424_ _2583_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4777_ _0294_ _3859_ as2650.r123\[0\]\[3\] as2650.r123\[0\]\[4\] _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6516_ _2177_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4941__A1 _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7496_ _3020_ _3124_ _3126_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6447_ _1888_ _2129_ _2046_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6694__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5497__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6378_ _1969_ _2050_ _2062_ _1944_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8117_ _0236_ clknet_leaf_61_wb_clk_i as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5329_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6727__C _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6446__A1 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8048_ _0167_ clknet_leaf_13_wb_clk_i as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6749__A2 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7558__C _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__C _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5421__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output11_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7174__A2 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7574__B _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5185__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4489__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6685__A1 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4160__A2 _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6988__A2 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7928__CLK clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5412__A2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _0435_ _0534_ _0549_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A2 _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5680_ as2650.psu\[3\] _1472_ _1483_ as2650.psu\[5\] _1486_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__7165__A2 _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7484__B _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5176__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4631_ _0370_ _0303_ _0439_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_129_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6912__A2 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7350_ _1802_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4923__A1 _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4923__B2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4562_ _0325_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _1823_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7281_ _1400_ _0706_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4493_ _3864_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6232_ _0576_ _0667_ _0780_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_89_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4151__A2 _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6163_ net24 _1862_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5114_ _0915_ _0916_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__B2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6094_ _3586_ _1794_ _1239_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5045_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7659__B _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__I _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6996_ _2650_ _2654_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6282__C _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6600__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5403__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5947_ as2650.pc\[9\] _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3965__A2 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5878_ _1628_ _1651_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7156__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7394__B _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7617_ _3219_ _3061_ _3243_ _2948_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4829_ _0316_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_43_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4914__A1 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7548_ _3114_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7479_ _3067_ _3068_ _3109_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6667__A1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4142__A2 _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3941__I as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6419__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6457__C _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4258__B _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7092__A1 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7092__B2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7395__A2 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6920__C _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7147__A2 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6699__I _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6370__A3 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6658__A1 _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7323__I _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7479__B _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5778__I as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6850_ as2650.stack\[5\]\[4\] _2402_ _2510_ as2650.stack\[6\]\[4\] _2514_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ as2650.stack\[2\]\[5\] _1584_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6781_ as2650.stack\[5\]\[3\] _2277_ _2445_ as2650.stack\[7\]\[3\] _2446_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3993_ _3525_ _3526_ _3527_ _3528_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5732_ _1533_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7138__A2 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5727__B _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5663_ _3667_ _3852_ _0402_ _0976_ _1096_ _1269_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7402_ _3665_ _3739_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6897__A1 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6402__I _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4614_ _0391_ as2650.r123\[0\]\[0\] _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6897__B2 _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5594_ _3816_ _0887_ _0307_ _0449_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_129_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7333_ as2650.stack\[7\]\[7\] _2967_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4545_ _0397_ _0398_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6649__A1 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7264_ _3650_ _2878_ _1392_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4476_ _3840_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6113__A3 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6215_ _1885_ _1800_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5321__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7195_ _1327_ _2845_ _2847_ _2849_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7233__I _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6146_ _3605_ _1831_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7074__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6077_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5624__A2 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6821__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _0868_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I wb_rst_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_58 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_69 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7377__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ _2513_ _2638_ _2639_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4060__A1 _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6888__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5560__A1 _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6104__A3 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7301__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4115__A2 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5863__A2 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4823__B1 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6040__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6222__I _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6879__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5926__I0 as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7540__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4354__A2 _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__A1 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4330_ as2650.r123\[0\]\[2\] _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6378__B _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5303__A1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4677__I _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _3751_ _3796_ _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6351__I0 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ _1736_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A2 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4192_ _3727_ as2650.addr_buff\[5\] _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7056__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7951_ _0070_ clknet_leaf_40_wb_clk_i as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6902_ _1689_ _2523_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7882_ _0001_ clknet_leaf_60_wb_clk_i as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7359__A2 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4290__A1 _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6833_ _1232_ _1975_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6031__A2 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _1840_ _2427_ _2428_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3976_ as2650.halted _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5715_ _1206_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4593__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6695_ _1577_ _2360_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5646_ _3667_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_108_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5542__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5577_ _1194_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7316_ as2650.stack\[7\]\[0\] _2962_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4896__A3 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4528_ _3689_ _3706_ _3878_ _3930_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_104_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5192__B _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4587__I _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6098__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7247_ _2044_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4459_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7178_ _2832_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6129_ _1830_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6022__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7770__A2 _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4584__A2 _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__A2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__A1 _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7286__A1 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__A2 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7038__A1 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6261__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4165__C _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7757__B _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4024__A1 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7761__A2 _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5500_ _3566_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ _1503_ _2150_ _2158_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7513__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5431_ _3671_ _1239_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4327__A2 _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5791__I _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ as2650.r123\[3\]\[7\] _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7101_ as2650.addr_buff\[3\] _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7277__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _3542_ _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8081_ _0200_ clknet_leaf_25_wb_clk_i as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5293_ _1077_ _1087_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7032_ _1612_ _0669_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4244_ _3753_ _3779_ _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4175_ as2650.r0\[0\] _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6788__B1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6252__A2 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7934_ _0053_ clknet_leaf_5_wb_clk_i as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7865_ _2022_ _3450_ _3455_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5966__I _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _1581_ _2425_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7796_ _0456_ _0457_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ _2359_ _2412_ _2159_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4566__A2 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5763__A1 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3959_ _3494_ _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5763__B2 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ _2271_ _2341_ _2344_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4318__A2 _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5629_ _0338_ _0731_ _1435_ _0739_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5634__C _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7268__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4097__A4 _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6491__A2 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4254__A1 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5876__I _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7296__C _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7961__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4557__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4309__A2 _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5506__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7259__A1 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5560__B _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6482__A2 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7431__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6234__A2 _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5980_ as2650.stack\[5\]\[3\] _1724_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4931_ net3 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6391__B _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5786__I _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7650_ net50 _3217_ _3125_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4862_ _3802_ _0683_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_60_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7734__A2 _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6601_ _2246_ _2265_ _2266_ _1672_ _2268_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7581_ _3205_ _3208_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4793_ _0622_ _0625_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_105_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6532_ _1017_ _2181_ _2203_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7498__A1 as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6463_ _2086_ _1555_ _2132_ _2144_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5414_ _1195_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6394_ _1407_ _2071_ _2078_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8133_ _0252_ clknet_leaf_5_wb_clk_i as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _1153_ _1155_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4720__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8064_ _0183_ clknet_leaf_15_wb_clk_i net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5276_ _0935_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7015_ _2478_ _2660_ _2674_ _2532_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7670__A1 _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4227_ _3502_ _3724_ _3760_ _3762_ _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5681__B1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4158_ _3693_ _3583_ _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4086__B _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7422__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6225__A2 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ _3624_ _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7917_ _0036_ clknet_3_4_0_wb_clk_i as2650.r123\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7848_ _2035_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7725__A2 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7779_ _1444_ _2033_ _3386_ _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5339__I1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7416__I _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6161__A1 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__A2 as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4475__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6990__I _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7413__A1 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7413__B2 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4227__A1 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4015__I _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5555__B _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7326__I _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5274__C _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4702__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5130_ _0935_ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5061_ _3900_ _0838_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5663__B1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5663__C2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4012_ _3545_ _3547_ _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5963_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4634__B _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7702_ _2764_ _3310_ _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4914_ _3645_ _3745_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5894_ _1663_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7707__A2 _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7633_ _2844_ _3258_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _0534_ _0537_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6341__S _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7564_ net34 _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4776_ _0294_ as2650.r123\[0\]\[3\] _0393_ _3859_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5194__A2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6391__A1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6515_ _2187_ _2188_ _2190_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7495_ net31 _3058_ _3125_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4941__A2 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6143__A1 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6446_ _1996_ _1336_ _2119_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6377_ _1385_ _1930_ _1933_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_88_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8116_ _0235_ clknet_3_3_0_wb_clk_i net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5328_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7643__A1 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6446__A2 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8047_ _0166_ clknet_leaf_13_wb_clk_i as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5259_ _1092_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8012__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5654__B1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__A3 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4544__B _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6382__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6050__I _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7590__B _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4696__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7634__A1 as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6437__A2 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6934__B _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5660__A3 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5269__C _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4630_ _0439_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6373__A1 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ as2650.r0\[1\] _0298_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4923__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _1987_ _1994_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7280_ _2927_ _2929_ _1400_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4492_ _0345_ _0343_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6231_ _3881_ _0494_ _1927_ _1928_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7873__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8035__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _1434_ _1322_ _1809_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7625__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5113_ _0946_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6428__A2 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6093_ _1799_ _1801_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _3598_ _0835_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6336__S _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _2650_ _2654_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _1698_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5877_ _1650_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7616_ _3239_ _3242_ _3014_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4828_ _0678_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4375__B1 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7547_ _3168_ _3175_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4914__A2 _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ _0595_ _0597_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_105_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6116__A1 _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7478_ _0287_ _0270_ _0276_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_107_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6667__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ _1217_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4678__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_12_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6419__A2 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4850__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7585__B _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5884__I _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5953__I1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8058__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6658__A2 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7855__A1 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7607__A1 _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7083__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5800_ _1594_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6780_ _1650_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3992_ _3488_ _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6594__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7495__B _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5731_ _3787_ _1511_ _1523_ _1425_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5794__I _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5662_ _1406_ _3661_ _0960_ _0286_ _0699_ _1098_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_136_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7401_ _3033_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4613_ _0416_ _0420_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6897__A2 _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5593_ _3661_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7332_ _1599_ _2961_ _2972_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4544_ _3649_ as2650.r123_2\[1\]\[4\] _3494_ _3863_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_102_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6649__A2 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7263_ _2858_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7846__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _0325_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6214_ _1366_ _1876_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5321__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7194_ _1819_ _2304_ _2848_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6145_ _1456_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5034__I _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7074__A2 _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6076_ _1244_ _1784_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5085__A1 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6282__B1 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _3511_ _0833_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6821__A2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4832__A1 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xwrapped_as2650_59 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7377__A3 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6978_ as2650.stack\[5\]\[7\] _2603_ _2535_ as2650.stack\[4\]\[7\] _2639_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ _1676_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6888__A2 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4899__A1 _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__A2 _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7837__A1 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7918__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5312__A2 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__I _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6503__I _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6879__A2 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5926__I1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5551__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4958__I _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6378__C _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4260_ _3795_ _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6500__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__I1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4191_ as2650.addr_buff\[6\] _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7056__A2 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6394__B _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7950_ _0069_ clknet_leaf_46_wb_clk_i as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4814__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6901_ as2650.pc\[6\] _1688_ _2523_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7881_ _0000_ clknet_leaf_60_wb_clk_i as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4290__A2 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _2492_ _2495_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6567__A1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _1841_ _1875_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3975_ _3491_ _3510_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5714_ _1511_ _1517_ _1518_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6319__A1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6694_ _1570_ _1537_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5645_ _0802_ _1206_ _3674_ _3815_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5917__I1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5576_ _1229_ _1315_ _1381_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5542__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7315_ _2960_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4527_ _3498_ _3876_ _0370_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7295__A2 _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7246_ _2296_ _2898_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4458_ _3600_ _3607_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_85_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7177_ _1328_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4389_ _3792_ _3766_ _3922_ _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_86_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6128_ as2650.addr_buff\[1\] _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6059_ _1696_ as2650.stack\[3\]\[8\] _1768_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7847__C _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6558__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6323__I _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6573__A4 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6730__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__A2 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6089__A3 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7890__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6494__B1 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7038__A2 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5402__I _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6261__A3 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7757__C _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6549__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5430_ _1238_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7492__C _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6721__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5361_ _1179_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7100_ _1620_ _2756_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _3846_ _3607_ _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8080_ _0199_ clknet_leaf_34_wb_clk_i as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7277__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5292_ _1065_ _1075_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5288__A1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7031_ _1700_ _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4243_ _3508_ _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4174_ _3642_ _3664_ _3709_ _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7933_ _0052_ clknet_leaf_5_wb_clk_i as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7864_ _3463_ _3464_ _2688_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _2333_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7201__A2 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7795_ _0737_ _1996_ _3401_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_51_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6746_ _2361_ _2376_ _2411_ _2127_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6960__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3958_ _3493_ _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5763__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6677_ as2650.stack\[7\]\[1\] _2342_ _2343_ as2650.stack\[6\]\[1\] _2344_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5628_ _3829_ _0730_ _0734_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_104_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8119__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5559_ _0359_ _1245_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7268__A2 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7229_ _2116_ _3881_ _2882_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6318__I _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7728__B1 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6400__B1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6951__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5754__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7259__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5690__A1 as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6228__I _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5132__I _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7431__A2 _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4245__A2 _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5442__A1 _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4930_ _0777_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _3749_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7195__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6600_ _2254_ _2267_ _2106_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7580_ _3165_ _3206_ _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4792_ _0637_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6531_ _2180_ _1096_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7498__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6462_ _1946_ _2140_ _2143_ _1442_ _1861_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5413_ _1220_ _1221_ _0822_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6393_ _2077_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5344_ _1170_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4181__A1 _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8132_ _0251_ clknet_leaf_10_wb_clk_i as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8063_ _0182_ clknet_leaf_15_wb_clk_i net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5275_ _1055_ _0830_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7014_ _2479_ _2673_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4226_ as2650.holding_reg\[0\] _3501_ _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4367__B _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5681__A1 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6138__I _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5681__B2 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4157_ _3638_ _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7422__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4088_ _3623_ _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_71_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5433__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_37_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7916_ _0035_ clknet_opt_2_0_wb_clk_i as2650.r123\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7186__A1 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7847_ _3447_ _3448_ _3449_ _2132_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7778_ _3385_ _1268_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6729_ _2118_ _2394_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8091__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7860__C _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6449__B1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7110__A1 _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7413__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6492__B _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4227__A2 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A2 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6511__I _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5555__C _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6667__B _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _3843_ _0880_ _0882_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7652__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5663__A1 _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4011_ as2650.cycle\[3\] _3546_ _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5663__B2 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5797__I as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4218__A2 _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5415__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5962_ as2650.stack_ptr\[0\] _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7701_ _3114_ _3323_ _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ _0598_ _0603_ _0635_ _0637_ _0642_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__7168__A1 _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5893_ _1589_ as2650.stack\[4\]\[4\] _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4206__I _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7632_ _1115_ _0773_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6915__A1 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ _0550_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7563_ net51 _3147_ _3149_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ _0598_ _0603_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6391__A2 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7517__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6514_ _2189_ _2187_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7494_ _0807_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6445_ _2108_ _2115_ _2124_ _2127_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7340__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6143__A2 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6376_ _1850_ _2059_ _1959_ _3526_ _2060_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8115_ _0234_ clknet_leaf_27_wb_clk_i net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5327_ _1158_ _1159_ _0826_ _0907_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_142_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7951__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7643__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8046_ _0165_ clknet_3_0_0_wb_clk_i as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5258_ _1089_ _1091_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5654__A1 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6851__B1 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__B2 _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4209_ _3744_ _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5189_ _3849_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4825__B _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5406__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5500__I _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__A1 _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3955__I _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6382__A2 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A1 _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6331__I _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7634__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5645__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6934__C _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5410__I as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__C _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6070__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7570__A1 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6373__A2 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6241__I _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4560_ _0326_ _0327_ _0328_ _0325_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4384__A1 _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4491_ _0341_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7974__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6230_ _0284_ _0384_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7873__A2 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6161_ _1853_ _1858_ _1860_ _1861_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_124_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7086__B1 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _0947_ _0948_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6092_ _3586_ _1800_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5636__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _3852_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5320__I _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6994_ _2573_ _2651_ _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ as2650.stack\[1\]\[8\] _1696_ _1697_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5876_ _1649_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7615_ _1602_ _3001_ _3241_ _2621_ _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4827_ _0488_ _0664_ _0657_ _0377_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_119_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7546_ _1846_ _1024_ _2827_ _3174_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4758_ _0604_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7691__B _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7477_ _1421_ _3040_ _3107_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6116__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4689_ _0531_ _0539_ _0436_ _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_134_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ _1527_ _2052_ _1853_ _1857_ _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4678__A2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7077__B1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7616__A2 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8029_ _0148_ clknet_leaf_17_wb_clk_i as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_52_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_130_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7866__B _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7585__C _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7001__B1 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4366__A1 _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7997__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7304__A1 as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4118__A1 _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7855__A2 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5405__I _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7607__A2 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5618__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5341__S _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5140__I _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4184__C _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3991_ _3487_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7791__A1 _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ _1531_ _1532_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5661_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7400_ _0315_ _1913_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4357__A1 _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ _0435_ _0462_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5592_ _1378_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7331_ as2650.stack\[7\]\[6\] _2967_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4543_ _0396_ as2650.r123\[1\]\[4\] _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7262_ _2866_ _0972_ _2869_ _2912_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4474_ _0326_ _0327_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ _1327_ _1906_ _1908_ _1910_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7193_ _3787_ _1266_ _1365_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6144_ _1846_ _1834_ _1847_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6657__I0 as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _3771_ _1339_ _3524_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_135_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5085__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6282__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5026_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6282__B2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5050__I _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7377__A4 _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ as2650.stack\[7\]\[7\] _2604_ _2601_ as2650.stack\[6\]\[7\] _2638_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ _1588_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7534__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5859_ as2650.stack\[6\]\[5\] _1637_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4899__A2 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7529_ _1430_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4520__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5076__A2 _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4284__B1 _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4823__A2 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6025__A1 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7773__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8025__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7525__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4304__I _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4190_ as2650.addr_buff\[6\] _3725_ _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7350__I _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6900_ _2522_ _2562_ _2045_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7880_ _2899_ _3476_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6016__A1 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6831_ _2493_ _2494_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7937__D _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6567__A2 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__B2 _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6762_ _1968_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3974_ _3497_ _3509_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5713_ _3497_ _1515_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6693_ _2242_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7516__A1 _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5378__I0 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5644_ _1159_ _1449_ _1450_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5575_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7314_ _2960_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4526_ _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4750__A1 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7245_ _2016_ _2885_ _2897_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5045__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4457_ _0311_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7176_ _2830_ _3740_ _2825_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4388_ _3812_ _3817_ _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_113_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6127_ _1453_ _1832_ _1835_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6255__A1 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6058_ _1603_ _1761_ _1772_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5009_ _3708_ _0844_ _0847_ _0849_ _0842_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8048__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__A2 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7755__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7507__A1 _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__I _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3963__I _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6730__A2 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6089__A4 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6494__A1 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6494__B2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7746__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6549__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5558__C as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4980__A1 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__I _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ as2650.r123\[3\]\[6\] _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4311_ as2650.addr_buff\[7\] _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5291_ _1058_ _1094_ _1092_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6485__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7030_ _1606_ _2658_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4242_ _3663_ _3765_ _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _3670_ _3696_ _3708_ _3695_ _3642_ _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__A1 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6788__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4209__I _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7932_ _0051_ clknet_leaf_5_wb_clk_i as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7863_ _2030_ _3461_ _3459_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7737__A1 _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6814_ _2477_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7908__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7794_ _1996_ _1401_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6745_ _2374_ _2399_ _2407_ _2410_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3957_ _3492_ _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6676_ _2274_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5627_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5558_ _1365_ _0799_ _1334_ _3490_ as2650.halted _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_133_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4509_ _0339_ _0340_ _3502_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5489_ _1292_ _0718_ _1296_ _0572_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_132_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6476__A1 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7228_ _1416_ _2875_ _2880_ _2881_ _2373_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_133_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7159_ _1674_ _1544_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5503__I _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4334__S0 _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7728__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7728__B2 _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6951__A2 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4962__A1 _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5506__A3 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4190__A2 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_7_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6219__A1 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5690__A2 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6244__I _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ _0704_ _0709_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7195__A2 _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4791_ _0639_ _0640_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6530_ _2179_ _2201_ _2202_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6461_ _1926_ _1974_ _2136_ _2141_ _2142_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4705__A1 _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5412_ as2650.psl\[6\] _0820_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6392_ _1919_ _1795_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8131_ _0250_ clknet_leaf_9_wb_clk_i as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5343_ _1110_ as2650.r123_2\[0\]\[6\] _1161_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8062_ _0181_ clknet_leaf_15_wb_clk_i net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _0876_ _1095_ _1106_ _1108_ _0871_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_102_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7013_ _2434_ _2664_ _2672_ _2377_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7024__B _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4225_ _3624_ _3688_ _3756_ _3760_ _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5681__A2 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4156_ _3679_ _3691_ _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6355__S _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4087_ _3568_ as2650.ins_reg\[3\] _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6225__A4 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5433__A2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7915_ _0034_ clknet_leaf_54_wb_clk_i as2650.r123\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7846_ _1292_ _3447_ _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5197__A1 _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5993__I _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7777_ _1258_ _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4989_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _2392_ _2328_ _2390_ _2391_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4944__A1 _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6659_ _1412_ _2259_ _2325_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6449__A1 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6449__B2 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6329__I _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5121__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6621__A1 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5408__I _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6688__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6667__C _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6239__I _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6860__A1 as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5663__A2 _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4010_ as2650.cycle\[2\] _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6612__A1 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5415__A2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _1538_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7700_ _1841_ _3321_ _3322_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4912_ _0625_ _0760_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5892_ _1653_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7168__A2 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7631_ _3205_ _3208_ _3256_ _3228_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _0531_ _3549_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6376__B1 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6915__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7562_ _3189_ _3190_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4774_ _0605_ _0623_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5974__I0 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6513_ _0908_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7493_ _1683_ _3022_ _3123_ _3056_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4222__I _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6444_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6858__B _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7340__A2 _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _1786_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8114_ _0233_ clknet_leaf_26_wb_clk_i net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5326_ _3534_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8045_ _0164_ clknet_leaf_1_wb_clk_i as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5103__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5257_ _1089_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5053__I _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7689__B _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4208_ _3743_ _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ _3571_ _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5406__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3968__A2 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7829_ as2650.overflow _3430_ _3159_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6906__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4560__C _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7331__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3971__I _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7095__A1 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5645__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6070__A2 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6723__S _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4908__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7570__A2 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6373__A3 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4384__A2 _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5581__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7858__B1 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4490_ _0341_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5582__B _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5333__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7353__I _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6160_ _1248_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5111_ as2650.r0\[2\] as2650.r123_2\[0\]\[1\] _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6091_ _1793_ _1794_ _1238_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5636__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6833__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5042_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4926__B _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7302__B _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5601__I _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6993_ _2617_ _2652_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6061__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4217__I _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ _1676_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4072__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5875_ as2650.stack_ptr\[1\] as2650.stack_ptr\[0\] _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_90_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7010__A1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7614_ _1694_ _3094_ _3092_ _3240_ _2337_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4826_ _3895_ _0655_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7561__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7545_ _3169_ _3172_ _3173_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4757_ _0607_ _0608_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7476_ _3044_ _3106_ _2075_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ _0539_ _0507_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6427_ _1556_ _2109_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7263__I _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6358_ _3519_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7077__A1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7077__B2 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5309_ _1130_ _1131_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ _1280_ _1966_ _1985_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6824__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8028_ _0147_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5511__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3966__I _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7001__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4366__A2 _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7304__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5315__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_opt_2_0_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7173__I _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7068__A1 _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5618__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6961__B _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4037__I _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7240__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ _3486_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7791__A2 _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _1228_ _1465_ _1466_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7941__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4611_ _0434_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5591_ _1398_ _0776_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7330_ _1594_ _2961_ _2971_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4542_ _3478_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7261_ _2872_ _2910_ _2911_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4473_ _0278_ _3835_ _3744_ _3838_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__6201__B _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6212_ _1505_ _1508_ _1909_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7192_ _1779_ _0572_ _2846_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6143_ _3606_ _1831_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6657__I1 as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6074_ _3548_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5025_ _3684_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6282__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4375__C _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__A1 _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7231__B2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6976_ _2599_ _2615_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6590__C _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5093__I0 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7782__A2 _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5927_ _1684_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5858_ _1640_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7534__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5545__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5789_ _1583_ _1567_ _1585_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7528_ _1588_ _3002_ _3157_ _1937_ _3014_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6345__I0 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7459_ _2991_ _2994_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6111__B _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4520__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7470__A1 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4284__A1 _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4284__B2 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6025__A2 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4036__A1 _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7964__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__B1 _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7773__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6981__B1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7525__A2 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6800__I _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7289__A1 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__I0 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7461__A1 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6247__I _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6264__A2 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__A2 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7213__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6830_ _2488_ _2438_ _2491_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4027__A1 _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6761_ _1582_ _2425_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4578__A2 _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3973_ _3499_ _3504_ _3508_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5712_ _1416_ _1512_ _1513_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6692_ _1578_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5527__A1 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5643_ as2650.psl\[7\] _1407_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5574_ _3491_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7313_ _2959_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4525_ _0377_ _0373_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6327__I0 _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5326__I _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7244_ _2862_ _2891_ _2896_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _3585_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7175_ _2070_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4387_ _3920_ _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6126_ _1833_ _1834_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6255__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6057_ as2650.stack\[3\]\[7\] _1766_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4266__A1 _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7987__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _3692_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4805__A3 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__A2 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__A3 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7755__A2 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6959_ _2616_ _2619_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4405__I _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7507__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6191__A1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7691__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7443__A1 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__A1 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__A1 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__A2 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A1 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4732__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4310_ _3841_ _3844_ _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5290_ _0879_ _1122_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7682__A1 _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4241_ _3776_ _3691_ _3756_ _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7361__I _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4172_ _3707_ _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__A2 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7931_ _0050_ clknet_leaf_11_wb_clk_i as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7310__B _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7862_ as2650.psu\[4\] _3462_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5748__A1 _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6813_ _2088_ _2323_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6945__B1 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7793_ _3400_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6744_ _2408_ _2361_ _2409_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3956_ as2650.ins_reg\[1\] _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _1650_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__S _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5626_ _1332_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5557_ _3618_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4508_ _3780_ _0355_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _0736_ _1282_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7122__B1 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7673__A1 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4439_ as2650.r0\[3\] _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7227_ _1400_ _0960_ _1940_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4487__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8015__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7158_ _1543_ _1544_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _1499_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7089_ _2112_ _2743_ _2746_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4334__S1 _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7220__B _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6615__I _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5451__A3 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7728__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4135__I _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6400__A2 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A4 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6467__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7664__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7181__I _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6219__A2 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7719__A2 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4650__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4790_ _0564_ _3744_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4402__A1 _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5585__B _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6460_ _1408_ _1322_ _2049_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6155__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5411_ _1219_ _3496_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6391_ _1850_ _2071_ _2075_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8038__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8130_ _0249_ clknet_leaf_11_wb_clk_i as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5342_ _1169_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7655__A1 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8061_ _0180_ clknet_leaf_15_wb_clk_i net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6458__A2 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5273_ _0907_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4469__A1 _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__I _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7012_ _2001_ _2666_ _2669_ _2378_ _2671_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4224_ _3757_ _3758_ _3759_ _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__7024__C _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5130__A2 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _3690_ _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _3584_ _3610_ _3613_ _3621_ _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_55_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6435__I _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7914_ _0033_ clknet_leaf_54_wb_clk_i as2650.r123\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4641__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7845_ _0908_ _2036_ _3440_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5197__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7776_ _1843_ _3382_ _3384_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4988_ _0825_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6727_ _2390_ _2391_ _2392_ _2328_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4944__A2 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6146__A1 _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ _3882_ _2324_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _0286_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_46_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6697__A2 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6589_ _3666_ _0939_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7646__A1 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5514__I _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5657__B1 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5121__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4880__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__A2 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6080__I _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6137__A1 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4699__A1 _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__I _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5415__A3 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5960_ _1708_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _0622_ _0643_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5891_ _1583_ _1654_ _1661_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7630_ _0782_ _0773_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4842_ _0358_ _0506_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6376__A1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6376__B2 _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6915__A3 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7561_ net51 _3058_ _3159_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4773_ _0607_ _0608_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4926__A2 _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6512_ _3816_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7492_ _1582_ _1812_ _2914_ _3103_ _3122_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6443_ _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6374_ _1817_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4659__B _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8113_ _0232_ clknet_leaf_27_wb_clk_i net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7628__A1 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5325_ _0803_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6300__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ _1032_ _1046_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8044_ _0163_ clknet_leaf_1_wb_clk_i as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5103__A2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ as2650.r123\[0\]\[0\] _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6851__A2 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5187_ _3847_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4138_ _3567_ _3674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4069_ as2650.addr_buff\[6\] _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4614__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7828_ _3426_ _3427_ _3433_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4917__A2 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7759_ _3612_ _1356_ _1506_ _1976_ _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7867__A1 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7867__B2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4550__B1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6803__I _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A2 _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5419__I _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5581__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7858__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7858__B2 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _0295_ _3684_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7086__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6090_ _3590_ _3602_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5097__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__I0 as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _0852_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6833__A2 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6597__A1 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6992_ _1693_ _1454_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5943_ _1609_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4072__A2 _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6349__A1 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5874_ _1648_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ _1449_ _3221_ _2118_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _0662_ _3637_ _3851_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5329__I _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7544_ _3169_ _3172_ _0314_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4756_ _0498_ _3743_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7849__A1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7475_ _0388_ _0380_ _3105_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4687_ _0359_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6426_ _3564_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6521__A1 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5324__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6357_ _2036_ _1334_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5308_ _1134_ _1135_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _1937_ _1965_ _1984_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5088__A1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6824__A2 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8027_ _0146_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _1072_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4835__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6588__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4063__A2 _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7001__A2 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_61_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5012__A1 _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6760__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3982__I _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__C _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5315__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7893__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7068__A2 _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5079__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5618__A3 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__A1 _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6579__A1 _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7240__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4054__A2 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5251__A1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4610_ _0441_ _0444_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_90_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5590_ _1378_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6751__A1 as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4541_ _0394_ as2650.r123_2\[0\]\[4\] as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\]
+ _3647_ _3493_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__4988__I _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4472_ _3861_ _3743_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5306__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7260_ _2830_ _0517_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6211_ _1331_ _1808_ _1878_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7191_ _1236_ _1895_ _1344_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6142_ _1483_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4937__B _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6073_ _1504_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5612__I _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _3742_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7231__A2 _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6975_ _2478_ _2615_ _2635_ _2532_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6443__I _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5926_ as2650.stack\[1\]\[3\] _1683_ _1677_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5857_ _1589_ as2650.stack\[6\]\[4\] _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _0514_ _0653_ _0655_ _3903_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5545__A2 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5788_ as2650.stack\[2\]\[3\] _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7527_ _2833_ _3152_ _3156_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4739_ _0369_ _0559_ _0590_ _0267_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_108_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7298__A2 _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7458_ _2386_ _3089_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6111__C _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6345__I1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ _2089_ _2092_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7389_ _3021_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4808__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__B2 _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7470__A2 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4138__I _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5233__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3977__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4036__A2 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__B2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6733__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5536__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7289__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6336__I1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5432__I _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7461__A2 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4027__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6760_ _1535_ _3573_ _1576_ _1570_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_50_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3972_ _3505_ _3507_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6972__A1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ _1511_ _1514_ _1516_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6691_ _2297_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5642_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6724__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5527__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7308__B _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4735__B1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5573_ _1380_ _1229_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5607__I _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7312_ _1628_ _2400_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7027__C _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4524_ _0318_ _0305_ _0371_ _0319_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6327__I1 _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7243_ _2858_ _0284_ _2859_ _0887_ _2895_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4455_ _0280_ _3716_ _0281_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4386_ as2650.holding_reg\[2\] _3872_ _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7174_ _2828_ _3731_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4667__B _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6125_ _1830_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6438__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6056_ _1599_ _1760_ _1771_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5007_ _3677_ _0835_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5498__B _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5215__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6173__I _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6558__A4 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7755__A3 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6958_ _2617_ _2618_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6963__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ _1626_ as2650.stack\[4\]\[12\] _1662_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6889_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _3482_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6191__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8094__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7140__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6348__I _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6792__B _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4257__A2 _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5206__A1 _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5757__A2 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6811__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6706__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7128__B _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6182__A2 _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7131__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4240_ _3775_ _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4496__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5693__A1 _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4171_ _3706_ _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5445__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7930_ _0049_ clknet_leaf_13_wb_clk_i as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4934__C _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7861_ _1423_ _3450_ _3456_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7198__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6812_ _2464_ _2467_ _2472_ _2475_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6945__A1 as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7792_ _1884_ _3398_ _3399_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5748__A2 _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6945__B2 as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _1854_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3955_ _3490_ _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ as2650.stack\[5\]\[1\] _2340_ _1714_ as2650.stack\[4\]\[1\] _2341_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5625_ _1321_ _1429_ _1432_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7370__A1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4184__A1 _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5556_ _1309_ _1265_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4507_ _3772_ _0357_ _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5487_ _0736_ _1282_ _1290_ _1291_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7954__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7226_ _1395_ _0883_ _2877_ _2879_ _3582_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4438_ _3648_ as2650.r123_2\[1\]\[3\] _3493_ _3863_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4487__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7157_ as2650.stack\[5\]\[12\] _2811_ _2812_ as2650.stack\[7\]\[12\] _2813_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4369_ _3554_ _3734_ _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6108_ _1816_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7088_ _2444_ _2744_ _2745_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5436__A1 _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _1759_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5800__I _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__A4 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6936__A1 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6936__B2 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7462__I _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__A2 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5427__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7352__A1 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6155__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ as2650.psl\[7\] _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7977__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6390_ _1799_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5341_ _1053_ _0501_ _1161_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7104__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5093__S _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8060_ _0179_ clknet_leaf_18_wb_clk_i as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5272_ _0660_ _0856_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4469__A2 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5666__A1 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7011_ _1608_ _2670_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_114_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4223_ as2650.holding_reg\[0\] _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4154_ _3689_ _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5418__A1 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4085_ _3620_ _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6091__A1 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout51_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7913_ _0032_ clknet_leaf_52_wb_clk_i as2650.r123\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4236__I _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7844_ _1460_ _2023_ _3438_ _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7775_ _1434_ _3382_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7591__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6394__A2 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6726_ _3883_ _2324_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6146__A2 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6657_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\] _0396_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5067__I _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5608_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6588_ _1519_ _2254_ _2255_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5539_ _1322_ _1327_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7646__A2 _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5657__A1 _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5016__B _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7209_ _2296_ _2863_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5657__B2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8189_ net47 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_15_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5530__I _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A1 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7582__A1 _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3985__I _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6361__I _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__A1 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__A1 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7406__B _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5705__I _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6845__B1 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5112__A3 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4320__A1 _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4871__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4910_ _0622_ _0643_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5890_ as2650.stack\[4\]\[3\] _1660_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5596__B _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4841_ _0684_ _0569_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6376__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8005__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ _3183_ _3188_ _3061_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4772_ _0606_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6511_ _0974_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7325__A1 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7491_ _3115_ _3117_ _3121_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6442_ _1957_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6373_ _2057_ _1326_ _1859_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5615__I _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4659__C _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8112_ _0231_ clknet_leaf_27_wb_clk_i net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5324_ _0828_ _1156_ _1157_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8043_ _0162_ clknet_leaf_14_wb_clk_i as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5255_ _0994_ _1047_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5103__A3 _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4206_ _3715_ _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5186_ _1017_ _0880_ _0882_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4137_ _3671_ _3672_ _3564_ _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_110_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4068_ _3600_ _3603_ _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4614__A2 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7827_ _3430_ _3432_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7564__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7758_ _3368_ _2323_ _2228_ _3370_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _2125_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6119__A2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7689_ _2726_ _3298_ _3312_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7867__A2 _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5645__A4 _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A1 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7307__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7858__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6530__A2 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5435__I _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5341__I0 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ _0840_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6991_ _2568_ _2616_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_92_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6597__A2 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7794__A1 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5942_ _1695_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7546__A1 _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6349__A2 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5873_ _1626_ as2650.stack\[6\]\[12\] _1639_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7612_ _3062_ _3234_ _3238_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8133__D _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4824_ _3632_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7543_ _3131_ _3170_ _3132_ _3171_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4755_ _0605_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7474_ _3075_ _3076_ _3104_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7849__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4686_ _0535_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6425_ _2107_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6356_ _2042_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ _1137_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7077__A3 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6287_ _1967_ _1983_ _1522_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6285__A1 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8026_ _0145_ clknet_leaf_32_wb_clk_i as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5238_ as2650.r0\[6\] _3684_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6176__I _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5169_ _0988_ _0996_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6588__A2 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7785__A1 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4852__C _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7537__A1 _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4424__I _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6760__A2 _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6276__A1 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7776__A1 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6579__A2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4054__A3 _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5251__A2 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7528__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7528__B2 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6751__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4762__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4471_ _3836_ _3838_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7700__A1 _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6210_ _3581_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4514__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7190_ _1886_ _2844_ _1330_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6141_ _1843_ _1834_ _1845_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7380__I _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6267__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _1780_ _1252_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_112_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5023_ _0857_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8128__D _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _1945_ _2628_ _2634_ _2246_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_65_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ as2650.pc\[3\] _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5856_ _1630_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _3737_ _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5787_ _1566_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7555__I _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7526_ _1587_ _2993_ _3155_ _1433_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4738_ _0585_ _0589_ _0369_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7457_ _2074_ _3064_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4669_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6408_ _2090_ _2091_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7388_ _1990_ _2161_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6339_ _2028_ _2011_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7290__I _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6258__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4808__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8009_ _0128_ clknet_leaf_37_wb_clk_i as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5233__A2 _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6981__A2 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4744__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6497__A1 _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6809__I _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6249__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7749__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6421__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3971_ _3506_ _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6972__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5710_ _1158_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6690_ _2296_ _2356_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4999__I _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5641_ _1406_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6724__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4735__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5572_ _0661_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7308__C _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4735__B2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7311_ _1114_ _2865_ _2958_ _2948_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4523_ _3728_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_117_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6488__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7242_ _0289_ _2875_ _2893_ _2894_ _1938_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _3854_ _3708_ _0291_ _0308_ _3631_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__A1 _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7173_ _2827_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6719__I _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5623__I _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4385_ _3773_ _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6124_ as2650.addr_buff\[0\] _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4239__I _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6055_ as2650.stack\[3\]\[6\] _1766_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5006_ _3666_ _0846_ _0844_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5498__C _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5215__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6412__A1 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4649__S1 _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7755__A4 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6957_ _2569_ _2573_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7883__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4974__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5908_ _1670_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6888_ _0495_ _2489_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5839_ _1626_ as2650.stack\[2\]\[12\] _1590_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7509_ _0372_ _0373_ _3138_ _0374_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_136_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7140__A2 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5151__A1 _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6629__I _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6792__C _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6364__I _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6403__A1 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5909__S _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6706__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7128__C _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7131__A2 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5142__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6890__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ _3705_ _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5445__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4653__B1 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6274__I _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7860_ _1485_ _3457_ _3460_ _3461_ _1986_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_36_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7198__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6811_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7791_ _3396_ _3389_ _1457_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6945__A2 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5819__S _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4956__A1 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6742_ _2051_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3954_ _3489_ _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6673_ _1546_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5624_ _1388_ _1372_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7370__A2 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5555_ _3676_ _1358_ _1360_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4506_ _0339_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5486_ _1292_ _0718_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7122__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5133__A1 as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7225_ as2650.psu\[1\] _2878_ _3597_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4437_ _3479_ as2650.r123\[1\]\[3\] _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6881__A1 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A2 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7156_ _1543_ _1711_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4368_ _3735_ _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _1548_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7087_ as2650.stack\[5\]\[10\] _2451_ _2287_ as2650.stack\[4\]\[10\] _2745_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4299_ _3699_ _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5436__A2 _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6038_ _1759_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6184__I _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7989_ _0108_ clknet_leaf_45_wb_clk_i as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8061__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4432__I _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5372__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5124__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6624__A1 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A2 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4938__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5374__S _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5340_ _1168_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5115__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5271_ _1104_ _1105_ _0856_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7010_ _1694_ _2623_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4222_ _3686_ _3758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5666__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4153_ _3688_ _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5418__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4084_ _3619_ _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6218__B _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7912_ _0031_ clknet_leaf_2_wb_clk_i as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8084__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7843_ _3444_ _3446_ _2688_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7040__A1 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4986_ _0822_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7774_ _1840_ _3382_ _3383_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6725_ _0285_ _2389_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _1872_ _1975_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7921__CLK clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5607_ _0894_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6587_ _1537_ _1519_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _1330_ _1337_ _1343_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_105_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6303__B1 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5469_ _1264_ _1277_ _1262_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6854__A1 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7208_ _2834_ _2841_ _2861_ _2862_ _0865_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__5657__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5016__C _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8188_ net47 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7139_ _2655_ _2691_ _2792_ _2794_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_59_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5811__I _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7231__C _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A2 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A1 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6909__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6642__I _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4162__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__A2 _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7406__C _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4320__A2 _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7270__A1 _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7022__A1 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ _3780_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7944__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4771_ _0604_ _0609_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6781__B1 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6510_ _2179_ _2184_ _2186_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7490_ _2099_ _3120_ _2867_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5336__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6441_ _2116_ _2117_ _2123_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7383__I _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6372_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8111_ _0230_ clknet_leaf_26_wb_clk_i net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7089__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5323_ as2650.r123_2\[2\]\[7\] _0875_ _0877_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8042_ _0161_ clknet_leaf_14_wb_clk_i as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5254_ _1061_ _1064_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_138_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4205_ _3720_ _3733_ _3740_ _3723_ _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_87_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5185_ _0561_ _0886_ _1020_ _0898_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5631__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ _3488_ _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7261__A1 _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4067_ _3590_ _3602_ _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_71_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7013__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7013__B2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7826_ _2068_ _2018_ _3431_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4378__A2 _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _0805_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7757_ _2473_ _3369_ _2098_ _1326_ _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6708_ _2364_ _2361_ _2372_ _2373_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7688_ _3305_ _3306_ _3311_ _2137_ _2832_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7316__A2 _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6119__A3 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__A1 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _2305_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5806__I _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__A2 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7226__C _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7252__A1 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4157__I _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7967__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5802__A2 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3996__I _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7004__A1 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6372__I _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5917__S _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7417__B _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5318__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5869__A2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7491__A1 _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__I _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5341__I1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7243__A1 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7243__B2 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6990_ _2649_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7794__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5941_ as2650.stack\[1\]\[7\] _1694_ _1686_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5872_ _1647_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7546__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7611_ _2616_ _3236_ _3237_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _3642_ _0663_ _0672_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8122__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7542_ _1478_ _0490_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4754_ _0391_ _3837_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7473_ _0287_ _0317_ _0320_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ _0463_ _0447_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5626__I _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6424_ _2106_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6355_ _2041_ _0737_ _2004_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5306_ _1070_ _1138_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_88_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6286_ _1979_ _1980_ _1982_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8025_ _0144_ clknet_leaf_32_wb_clk_i as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5237_ _1069_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4296__A1 _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ _0997_ _1004_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_84_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4119_ _3480_ as2650.r123\[1\]\[7\] _3655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4048__A1 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5099_ _0312_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7785__A2 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6192__I _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7537__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5548__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7809_ _1154_ _3402_ _3414_ _3415_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_125_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6745__B1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4440__I _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__A1 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__B2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6367__I _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6276__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A2 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7225__A1 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__A1 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7776__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7528__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5539__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4211__A1 _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5446__I _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4762__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4470_ _3681_ as2650.r123\[0\]\[2\] _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6140_ _1844_ _1837_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7464__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6267__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ _1779_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5181__I _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _3740_ _0859_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7610__B _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7767__A2 _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6973_ _2630_ _2632_ _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ _1682_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5855_ _1583_ _1631_ _1638_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _0569_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5786_ _1582_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7525_ _2373_ _1528_ _3154_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4737_ _0316_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7456_ _3062_ _3087_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7152__B1 _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4668_ _3802_ _0465_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6896__B _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6407_ _1272_ _1971_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5702__A1 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7387_ _3017_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8018__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4599_ _0436_ _0448_ _0451_ _3919_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ _0492_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6258__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6269_ net25 _1965_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4269__A1 _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8008_ _0127_ clknet_leaf_36_wb_clk_i as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7758__A2 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__B1 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A2 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6194__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4744__A2 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5266__I _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4170__I _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6497__A2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5215__B _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6249__A2 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5930__S _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3970_ as2650.ins_reg\[7\] _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4983__A2 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ _1113_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5571_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4735__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4522_ _0275_ _0371_ _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7310_ _2951_ _2957_ _2864_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__A2 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7605__B _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4453_ _3857_ _0307_ _3888_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7241_ _2839_ _2188_ _2197_ _1398_ _1940_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7391__I _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4499__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7172_ _2826_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6001__S _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5160__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4384_ _3917_ _3874_ _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_113_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7437__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6123_ _1831_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6054_ _1594_ _1760_ _1770_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__A1 _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6956_ _1597_ _1454_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ _1622_ as2650.stack\[4\]\[11\] _1662_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6887_ _2308_ _2544_ _2546_ _1873_ _2549_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5838_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5769_ as2650.stack\[2\]\[0\] _1568_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7508_ _0275_ _0371_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7125__B1 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7676__A1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7515__B _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7439_ _2844_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4858__C _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5151__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6100__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7250__B _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6651__A2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6403__A2 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7600__A1 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4414__A1 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__A1 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6706__A3 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7667__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__I _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7419__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4653__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4653__B2 _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4075__I _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7198__A3 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6810_ _2473_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7790_ _1434_ _0972_ _3397_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6741_ _2401_ _2403_ _2406_ _1264_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_90_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3953_ _3485_ _3486_ _3487_ _3488_ _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__6290__I _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6158__A1 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7355__B1 _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6672_ _2051_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5623_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5554_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7658__A1 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4505_ _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5485_ _0705_ _0718_ _0723_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ _3678_ _0284_ _0290_ _3694_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7224_ _2835_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6330__A1 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4367_ _3719_ _3900_ _3901_ _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7155_ _1674_ _1711_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ _1265_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7086_ as2650.stack\[7\]\[10\] _2445_ _2448_ as2650.stack\[6\]\[10\] _2744_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ _3832_ _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4694__B _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6037_ _1758_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7988_ _0107_ clknet_leaf_49_wb_clk_i as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6939_ _2284_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4947__A2 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5809__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7649__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__B2 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5544__I _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3999__I _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6375__I _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7821__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6388__A1 _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4938__A2 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5060__A1 _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7352__A3 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6560__A1 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5454__I _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7104__A3 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5270_ _1024_ _1025_ _0679_ _0858_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4221_ _3683_ _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4152_ _3687_ _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__B _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7812__A1 _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4083_ _3483_ _3514_ _3618_ _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_95_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__C _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7911_ _0030_ clknet_leaf_2_wb_clk_i as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7842_ _3438_ _3445_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6379__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7040__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__A2 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7773_ _2108_ _3382_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4985_ _0800_ _0824_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4533__I _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6724_ _0285_ _2389_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7879__A1 as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7879__B2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6655_ _2062_ _2299_ _2321_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5606_ _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6551__A1 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _1536_ _3665_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7065__B _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5537_ _1214_ _1237_ _1212_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6303__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6303__B2 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5468_ _1268_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7207_ _2857_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4419_ _3872_ _0273_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_8187_ net47 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4865__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5399_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7138_ as2650.pc\[11\] _1097_ _2793_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4708__I _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7803__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7069_ _2364_ _2720_ _2726_ _2107_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A3 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6790__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7896__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6845__A2 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4608__A1 _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5959__I1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4353__I _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4770_ _0592_ _0612_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6440_ _2120_ _2122_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6533__A1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6371_ _1816_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8110_ _0229_ clknet_leaf_27_wb_clk_i net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5322_ _1153_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8041_ _0160_ clknet_leaf_50_wb_clk_i net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _1077_ _1087_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5912__I _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4204_ _3739_ _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5184_ _0706_ _0890_ _0891_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4135_ _3487_ _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ as2650.cycle\[7\] _3601_ _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5272__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6743__I _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7013__A2 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7825_ _3385_ _2017_ _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4263__I _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7756_ _1214_ _1560_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _0430_ _0806_ _0813_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6707_ _2106_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7687_ _3309_ _3310_ _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4899_ _3714_ as2650.r123\[0\]\[7\] _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6119__A4 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5327__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6638_ _1815_ _2304_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6569_ _1210_ _1786_ _1825_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_106_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4838__A1 _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7242__C _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7252__A2 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6763__A1 _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7417__C _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5318__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8074__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5732__I _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4348__I _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7911__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7243__A2 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5940_ _1693_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ _1622_ as2650.stack\[6\]\[11\] _1639_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5006__A1 _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7610_ _2616_ _3236_ _2099_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ _3695_ _3660_ _0403_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6754__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7541_ _1478_ _0490_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4753_ _0472_ _0473_ _0470_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4811__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7472_ _1683_ _1233_ _2721_ _3102_ _2035_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4684_ _0442_ _0458_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6423_ _2053_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6354_ _1447_ _2040_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5305_ _0278_ _0501_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6285_ _1981_ _1504_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5642__I _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8024_ _0143_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7482__A2 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5236_ _1036_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5493__A1 _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _0999_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4118_ _3646_ _3651_ _3653_ _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5098_ _0434_ _0346_ _0365_ _0366_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5245__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4048__A2 _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ _3499_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7808_ _1055_ _0723_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6745__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5548__A2 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7739_ _3913_ _3354_ _3358_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6422__B _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5817__I _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4220__A2 _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8097__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__B1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7225__A2 _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4039__A2 _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6383__I _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6984__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5539__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4211__A2 _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7161__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5462__I _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _0831_ _0938_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A1 _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4078__I _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5021_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7389__I _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6972_ _2216_ _2493_ _2498_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6975__A1 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5923_ as2650.stack\[1\]\[2\] _1681_ _1677_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5854_ as2650.stack\[6\]\[3\] _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4805_ _0400_ _0482_ _0506_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5785_ _1581_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5637__I _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4202__A2 _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7524_ _2245_ _2471_ _2995_ _3153_ _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4736_ _0587_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7455_ _3065_ _3086_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4667_ _0479_ _0481_ _0519_ _0333_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7152__A1 _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6896__C _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7957__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6406_ _1818_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7386_ _3015_ _3019_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5702__A2 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _0356_ _0449_ _0450_ _0436_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6337_ _2027_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7455__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6268_ _1903_ _1935_ _1964_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_130_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8007_ _0126_ clknet_leaf_43_wb_clk_i as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5219_ _1016_ _1054_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6199_ _1819_ _1341_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7758__A3 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__A2 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__A1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__B2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4451__I _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3952__A1 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__A1 as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8112__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6841__I _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4983__A3 _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5457__I _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4196__A1 _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _1376_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4521_ _0372_ _0373_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7134__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7240_ as2650.overflow _1231_ _2892_ _1444_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4452_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4499__A2 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5696__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ _1799_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4383_ as2650.holding_reg\[2\] _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6122_ _1830_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7437__A2 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7621__B _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ as2650.stack\[3\]\[5\] _1766_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4120__A1 _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5004_ _3572_ _0824_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4536__I as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6948__A1 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6955_ as2650.pc\[7\] net2 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5620__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5906_ _1617_ _1655_ _1669_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6886_ _2430_ _2528_ _2547_ _2548_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5837_ _1624_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5768_ _1566_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7507_ _1480_ _3040_ _3134_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _3541_ _3876_ _0485_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5699_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7676__A2 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7438_ _3068_ _3069_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6723__I1 as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5687__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_49_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8135__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6198__I _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7369_ _1194_ _1926_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5830__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6100__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7250__C _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4414__A2 _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7364__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__A2 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7116__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7667__A2 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5941__S _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7419__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4350__A1 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__I as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4102__A1 _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4653__A2 _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7198__A4 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8008__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6740_ as2650.stack\[3\]\[2\] _1651_ _2400_ as2650.stack\[2\]\[2\] _2405_ _2406_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ as2650.cycle\[3\] as2650.cycle\[2\] _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6671_ _2337_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7355__A1 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5187__I _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6158__A2 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7355__B2 _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4169__A1 _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ _3513_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5905__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7107__A1 as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5553_ _3672_ _1250_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6012__S _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4504_ _3503_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5484_ as2650.psl\[1\] _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5669__A1 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7223_ _1292_ _2876_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4435_ _0289_ _3678_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5851__S _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4341__A1 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7154_ _2798_ _2809_ _1898_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4366_ _3621_ _3721_ _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6105_ _1810_ _1811_ _1813_ _1360_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7085_ _2679_ _2741_ _2742_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4297_ _3806_ _3831_ _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _1543_ _1675_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4644__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7987_ _0106_ clknet_leaf_33_wb_clk_i as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6481__I _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6938_ _2599_ _2567_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7346__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6869_ _2125_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5380__I0 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7821__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4176__I _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7585__A1 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6388__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4399__A1 _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5735__I as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6560__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4220_ as2650.holding_reg\[0\] _3623_ _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4874__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4151_ _3683_ _3686_ _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_95_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5470__I _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4082_ _3617_ _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7812__A2 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7910_ _0029_ clknet_leaf_62_wb_clk_i as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7841_ _2020_ _1967_ _3440_ _2022_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7576__A1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7772_ _0860_ _1871_ _1512_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4984_ _3484_ _0823_ _3562_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6723_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _3480_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7879__A2 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6654_ _2308_ _2312_ _2320_ _2060_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5605_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6585_ _2252_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6250__B _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4562__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ _1203_ _1247_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5467_ as2650.psu\[5\] _1271_ _1273_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6303__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__A1 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7206_ _2857_ _2860_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4418_ _3757_ _3758_ _3701_ _3704_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8186_ net46 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ _1206_ _3674_ _3935_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7137_ _2764_ _2723_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _3668_ _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7068_ _2721_ _2725_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7803__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6019_ _1749_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7016__B1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__B2 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6790__A2 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A2 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4599__C _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6386__I _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6058__A1 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7255__B1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7558__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7558__B2 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6230__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6781__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7730__A1 _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__B2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4544__A1 _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _2051_ _2052_ _1895_ _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5321_ _1154_ _0871_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6297__B2 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8040_ _0159_ clknet_leaf_46_wb_clk_i net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7990__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5252_ _1085_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_114_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4203_ _3724_ _3738_ _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__I _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5183_ _0576_ _0892_ _0893_ _1018_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6049__A1 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ _3667_ _3669_ _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4065_ as2650.cycle\[5\] _3588_ _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5272__A2 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7549__A1 _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7824_ _2068_ _3428_ _3394_ _3429_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4967_ as2650.r123\[1\]\[3\] _0809_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7755_ _2430_ _2473_ _2548_ _1818_ _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6899__C _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6706_ _1383_ _2090_ _2371_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7686_ _3307_ _3308_ _2765_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4898_ _0392_ _0299_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6637_ _1821_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4535__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6568_ _1367_ _1341_ _2235_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5519_ _0312_ _1324_ _1247_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6499_ _1995_ _1781_ _2174_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__6288__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7788__A1 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6460__A1 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6763__A2 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7712__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6279__A1 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7779__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__I _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6451__A1 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5870_ _1617_ _1632_ _1646_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6203__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4821_ _3669_ _0667_ _0671_ _3886_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6754__A2 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7540_ _0580_ _0588_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4752_ _0598_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4765__A1 as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7471_ _2048_ _2421_ _3101_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4683_ _0530_ _0533_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6506__A2 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _2087_ _2105_ _2045_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4517__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5190__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6353_ _1525_ _1529_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5304_ as2650.r0\[7\] _0866_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6284_ _0781_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8023_ _0142_ clknet_leaf_36_wb_clk_i as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4539__I as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5235_ _0498_ _3867_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6690__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5166_ _1001_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4117_ _3533_ _3652_ _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ _0822_ _0826_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4048_ _3572_ _3583_ _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_37_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7886__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7807_ _0711_ _0723_ _3411_ _3412_ _3413_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4205__B1 _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6745__A2 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5999_ _1622_ as2650.stack\[5\]\[11\] _1726_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4756__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7738_ _3839_ _3356_ _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7669_ net37 _3217_ _3125_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4508__A1 _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5833__I _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7709__B _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8041__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4211__A3 _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7444__B _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6839__I _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4359__I _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _3484_ _3537_ _0860_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6574__I _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6971_ _2583_ _2631_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _1578_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4986__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ _1630_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4738__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ _0569_ _0654_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5784_ as2650.pc\[3\] _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7523_ _2427_ _3150_ _2485_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _0488_ _0507_ _0555_ _0377_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_7454_ _1795_ _3082_ _3084_ _3085_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7688__B1 _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _0412_ _0512_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6405_ _3525_ _2047_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5163__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7385_ _2988_ _3018_ _2159_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5653__I _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4597_ _0443_ _0356_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6336_ _2025_ _0339_ _2026_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _1376_ _1908_ _1956_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6663__A1 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5466__A2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8006_ _0125_ clknet_leaf_37_wb_clk_i as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5218_ _0935_ _1053_ _0970_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6198_ _1784_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6484__I _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ _0920_ _0955_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5218__A2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__A2 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8064__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4977__A1 as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4729__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7901__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4888__B _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7143__A2 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7264__B _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4179__I _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6654__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5209__A2 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4128__B _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6957__A2 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4968__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4642__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7382__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__A2 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5393__A1 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _0272_ _0340_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_117_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4451_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6893__A1 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5696__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7170_ _2384_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4382_ _3809_ _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ _1798_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5448__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6052_ _1769_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _0843_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4817__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8087__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4120__A2 as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7070__A1 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5849__S _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4959__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6954_ _2614_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5905_ as2650.stack\[4\]\[10\] _1657_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__I _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6885_ _1210_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4552__I _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5836_ as2650.pc\[12\] _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7924__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5767_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7506_ _3044_ _3135_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4718_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5698_ _1500_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7125__A2 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7437_ _1417_ _0277_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4649_ _0500_ _0501_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _3479_ _3494_
+ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_135_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _3001_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6319_ _0908_ _2011_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7299_ _2044_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_18_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4727__I _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6942__I _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7364__A2 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__A3 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__I _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5127__A1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5507__B _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6875__A1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6627__A1 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4102__A2 _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7947__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ as2650.cycle\[7\] as2650.cycle\[6\] as2650.cycle\[5\] as2650.cycle\[4\] _3487_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6670_ _0937_ _1870_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7355__A2 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _1372_ _1428_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4169__A2 _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5552_ _1359_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4503_ _0356_ _0305_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5483_ _0692_ _0731_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5669__A2 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4434_ _0288_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7222_ _1230_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7153_ _2266_ _2791_ _2808_ _2246_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4365_ _3898_ _3899_ _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4341__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ _3514_ _1812_ _1782_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7084_ as2650.stack\[1\]\[10\] _2451_ _2448_ as2650.stack\[2\]\[10\] _2742_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4296_ _3810_ _3813_ _3828_ _3830_ _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_112_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6248__B _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4547__I _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7291__A1 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6035_ _1757_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5841__A2 _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__A1 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6762__I _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7986_ _0105_ clknet_leaf_34_wb_clk_i as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6937_ _2337_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6868_ _2474_ _2529_ _2530_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8102__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5819_ _1610_ as2650.stack\[2\]\[8\] _1590_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6799_ _1588_ _2359_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7526__C _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__A1 _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6937__I _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5380__I1 as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4457__I _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7282__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6672__I _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7585__A2 _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5596__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7337__A2 _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7717__B _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6560__A3 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6848__A1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5520__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ as2650.ins_reg\[0\] _3685_ _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__A2 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7273__A1 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4081_ _3616_ _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4087__A1 _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7840_ _3443_ _3438_ as2650.psl\[3\] _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8125__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7771_ _3375_ _3380_ _3381_ _2948_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6784__B1 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4983_ _3483_ _0823_ _3552_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_51_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ _2378_ _2379_ _2382_ _2387_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6653_ _1438_ _2316_ _2319_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5604_ _3666_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4011__A1 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6584_ as2650.addr_buff\[0\] _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ _1338_ _1263_ _1340_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_106_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5466_ _1270_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7362__B _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4417_ _0271_ _3904_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7205_ _2858_ _3692_ _2859_ _3784_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4314__A2 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8185_ net46 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5397_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5661__I _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7136_ _2722_ _2763_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4348_ _3882_ _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7264__A1 _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7067_ _2722_ _2724_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4279_ _3808_ _3771_ _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _1685_ as2650.stack\[0\]\[4\] _1748_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7969_ _0088_ clknet_leaf_40_wb_clk_i as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5836__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5750__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4305__A2 _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5502__A1 _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6058__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4187__I _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7255__A1 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7255__B2 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7007__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6230__A2 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A1 _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7447__B _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7730__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4544__A2 as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5320_ _0741_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6297__A2 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ _0278_ _0992_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4202_ _3735_ _3737_ _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5182_ _0580_ _0977_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7246__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4133_ _3668_ _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__A2 _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ as2650.addr_buff\[7\] _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__S _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5009__B1 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7549__A2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7823_ _2107_ _1445_ _3391_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5857__S _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7754_ _2992_ _2226_ _2995_ _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4966_ _0335_ _0806_ _0812_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4232__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6705_ _2365_ _2369_ _2370_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7685_ _2765_ _3307_ _3308_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_123_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4897_ _0279_ _0500_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6636_ _2301_ _2302_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5327__A4 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6567_ _1361_ _1917_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5518_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6498_ _1318_ _1326_ _1856_ _1815_ _0860_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5449_ _3497_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7237__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7119_ _2363_ _2755_ _2775_ _2474_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8099_ _0218_ clknet_leaf_43_wb_clk_i as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7788__A2 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5566__I _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7476__A1 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6279__A2 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__B1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7228__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7779__A2 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__A3 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6451__A2 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7400__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6203__A2 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4820_ _0670_ _3875_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A1 _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4751_ _0601_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5476__I _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7470_ _1421_ _2057_ _2995_ _3100_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4682_ _0530_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6421_ _1340_ _2097_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6352_ _2039_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5190__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7467__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ as2650.r123_2\[0\]\[7\] _1132_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6283_ net25 _1526_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8022_ _0141_ clknet_leaf_36_wb_clk_i as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7219__A1 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5165_ _0294_ as2650.r123_2\[0\]\[1\] _3867_ as2650.r0\[2\] _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5493__A3 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4116_ as2650.r123\[2\]\[7\] as2650.r123_2\[2\]\[7\] _3479_ _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _0828_ _0933_ _0934_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6978__B1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4047_ _3577_ _3582_ _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7806_ _0552_ _0694_ _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _1734_ _1718_ _1735_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__B2 _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7737_ _3798_ _3354_ _3357_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4949_ _0798_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5386__I _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7668_ _1700_ _3021_ _3288_ _1991_ _3292_ _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_123_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6619_ _1712_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7599_ _3223_ _3224_ _3225_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7458__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6130__A1 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6681__A2 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4692__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8084__D _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7630__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6197__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7980__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4747__A2 _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5795__I1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7449__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7621__A1 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6970_ _2588_ _2593_ _2629_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4435__A1 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5921_ _1680_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6188__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5852_ _1636_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ _0528_ _0484_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5783_ _1580_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7522_ _3051_ _3130_ _3151_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4734_ _0319_ _0556_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7688__A1 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7688__B2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7453_ _2078_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4665_ _3909_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _2000_ _1934_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7384_ _3017_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6360__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ _0440_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6335_ _2004_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6112__A1 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6266_ _1912_ _1961_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _0124_ clknet_leaf_31_wb_clk_i as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6663__A2 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5217_ _1028_ _1051_ _1052_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7860__A1 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7860__B2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4674__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6197_ _1265_ _3536_ _1199_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5148_ _0517_ _0903_ _0943_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7612__A1 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5079_ _0279_ _0866_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6179__A1 _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7376__B1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6005__I _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7679__A1 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7280__B _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7851__A1 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4968__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5090__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6590__A1 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6590__B2 _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4450_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4381_ _3518_ _3915_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ _1807_ _1809_ _1814_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7842__A1 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6051_ _1685_ as2650.stack\[3\]\[4\] _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _3583_ _0824_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4408__A1 _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6948__A3 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7070__A2 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _1693_ _2563_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4959__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5929__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5904_ _1614_ _1655_ _1668_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5620__A3 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6026__S _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6884_ _1520_ _2524_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5835_ _1623_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5865__S _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6581__A1 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5766_ _1565_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7505_ _3131_ _3133_ _3132_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4717_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5664__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5697_ _3515_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ _0270_ _0276_ _0287_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4648_ as2650.r123_2\[0\]\[5\] _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6333__A1 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6884__A2 _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7367_ _1870_ _1364_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4579_ _3518_ _0432_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4895__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ _2006_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7298_ _2940_ _2946_ _2865_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7833__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _1812_ _1941_ _1945_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_58_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6572__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7899__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5574__I _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A2 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7521__B1 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7824__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7052__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5749__I _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3950_ as2650.cycle\[0\] _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ _1374_ _1405_ _1411_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6563__A1 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5551_ _1308_ _1209_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _3776_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6315__A1 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _0535_ _0536_ _1287_ _1288_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_133_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7221_ _3675_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4433_ _0287_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6866__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8054__CLK clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7152_ _1446_ _2804_ _2806_ _2251_ _2807_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4364_ _3894_ _3897_ _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ _3674_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4828__I _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7083_ as2650.stack\[3\]\[10\] _2445_ _2447_ as2650.stack\[0\]\[10\] _2741_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4295_ _3782_ _3817_ _3829_ _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7204__I _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6094__A3 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7291__A2 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6034_ _1707_ as2650.stack\[0\]\[12\] _1748_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5841__A3 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7985_ _0104_ clknet_leaf_49_wb_clk_i as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6936_ _2478_ _2567_ _2597_ _2503_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4801__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6867_ _2266_ _2524_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5818_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6554__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6798_ _1583_ _2244_ _2462_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4565__B1 _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4512__B _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5394__I _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5749_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7419_ _1535_ net5 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7823__B _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6439__B _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7034__A2 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__I _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6793__A1 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4859__A1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5520__A2 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ _3615_ _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7273__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4087__A2 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5284__A1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4383__I as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7770_ as2650.stack_ptr\[2\] _3375_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6784__A1 as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ as2650.halted _3519_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6784__B2 as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6721_ _2383_ _2384_ _1233_ _2386_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_3_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _1211_ _2317_ _2318_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5603_ _1408_ _1410_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6583_ _2060_ _2250_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5534_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5465_ _3553_ _1208_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7204_ _2161_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4416_ _3736_ _3555_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8184_ net46 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5396_ _3573_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7135_ _2790_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4347_ net6 _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7264__A2 _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7066_ _2655_ _2691_ _2723_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4278_ _3812_ _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5275__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _1739_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7016__A2 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A1 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6775__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7968_ _0087_ clknet_leaf_41_wb_clk_i as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6919_ _2548_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7818__B _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7899_ _0018_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4250__A2 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7724__B1 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__A2 _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5750__A2 _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7937__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4305__A3 _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5502__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8087__D _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7255__A2 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7007__A2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5018__A1 _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6766__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4241__A2 _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4931__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7191__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5250_ _1083_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ _3736_ _3555_ _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5181_ _0560_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4132_ _3638_ _3572_ _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4063_ _3592_ _3598_ _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5009__A1 _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4480__A2 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7822_ _1419_ _2015_ _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7753_ _0795_ _3361_ _3366_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4965_ as2650.r123\[1\]\[2\] _0809_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4232__A2 _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6704_ _2367_ _2368_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6509__A1 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6034__S _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7684_ _3277_ _3246_ _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4896_ _3842_ as2650.r123\[0\]\[6\] _0598_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6635_ as2650.pc\[1\] net6 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7182__A1 _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__S _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _1324_ _1216_ _1907_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7373__B _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5517_ _3611_ _1215_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5672__I _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6497_ _3676_ _1360_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5448_ _1228_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6288__A3 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5496__A1 _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5379_ _1190_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7118_ _2305_ _2768_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8098_ _0217_ clknet_leaf_39_wb_clk_i as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7049_ as2650.stack_ptr\[2\] as2650.stack\[3\]\[9\] _2447_ as2650.stack\[0\]\[9\]
+ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A3 _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4471__A2 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5971__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6920__A1 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8115__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__B2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7730__C _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6987__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6451__A3 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4462__A2 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6739__A1 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7400__A2 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A2 _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5411__A1 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _0295_ _3865_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3973__A1 _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4681_ _0531_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7164__A1 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6420_ _2098_ _2102_ _2103_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_122_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _2038_ _0700_ _2026_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5190__A3 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ _3713_ as2650.r123_2\[0\]\[7\] _1132_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7467__A2 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6282_ _1812_ _1856_ _1946_ _1970_ _1978_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8021_ _0140_ clknet_leaf_36_wb_clk_i as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5233_ _0498_ _3702_ _3868_ _0390_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7219__A2 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ _0949_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4115_ _3650_ as2650.r123\[0\]\[7\] _3495_ _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ as2650.r123_2\[2\]\[2\] _0875_ _0877_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7212__I _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _3578_ _3581_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__A2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7805_ _3403_ _0465_ _0552_ _0694_ _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ as2650.stack\[5\]\[10\] _1720_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7736_ _3745_ _3356_ _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4948_ _0524_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7667_ _2422_ _2694_ _3291_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4879_ _0717_ _0727_ _0691_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6618_ _1545_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6902__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7598_ _3223_ _3224_ _1023_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8138__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6549_ as2650.psu\[7\] _1408_ _1353_ _2217_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5469__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6130__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4141__A1 _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7630__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6197__A2 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5577__I _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4481__I _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7146__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7697__A2 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7449__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4380__A1 as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4380__B2 _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4132__A1 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4435__A2 _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ as2650.stack\[1\]\[1\] _1679_ _1677_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ _1579_ as2650.stack\[6\]\[2\] _1634_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7385__A1 _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6188__A2 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4802_ _0564_ _3618_ _0566_ _3523_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_94_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5782_ _1579_ as2650.stack\[2\]\[2\] _1574_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7521_ _1921_ _3146_ _3150_ _1800_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4733_ _0560_ _3637_ _3851_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7137__A1 _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7452_ _2368_ _3083_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4664_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6403_ _2086_ _3525_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7383_ _3016_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4595_ _0445_ _0447_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6334_ _2021_ _2024_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _1263_ _1395_ _1906_ _1237_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_103_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6112__A2 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8004_ _0123_ clknet_leaf_30_wb_clk_i as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5216_ _0553_ _0942_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6267__B _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6196_ _1780_ _1893_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4674__A2 _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5147_ _0491_ _0882_ _0879_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5078_ _0915_ _0916_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4029_ _3527_ _3528_ _3564_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_37_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5397__I _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7376__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7376__B2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7719_ _1801_ _3338_ _3340_ _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7128__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6887__B1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4362__A1 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7561__B _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7300__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7851__A2 _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A1 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4665__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5614__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7367__A1 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5100__I _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7119__A1 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6640__B _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6590__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4380_ as2650.r123\[2\]\[1\] _3636_ _3914_ _3800_ _3915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A1 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _1759_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input7_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5001_ _3640_ _0824_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4656__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4408__A2 _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6952_ _2298_ _2612_ _2613_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5903_ as2650.stack\[4\]\[9\] _1657_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6883_ _3725_ _2327_ _2545_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5620__A4 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6106__I _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5834_ _1622_ as2650.stack\[2\]\[11\] _1590_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7646__B _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5765_ _1541_ _1547_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6581__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7504_ _3131_ _3132_ _3133_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4716_ _0562_ _0563_ _0565_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7365__C _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5696_ _1500_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7435_ _1459_ _3906_ _3907_ _3035_ _3036_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4647_ as2650.r123\[0\]\[5\] _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6333__A2 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7366_ _2990_ _2999_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4578_ as2650.r123\[2\]\[3\] _3636_ _0431_ _3800_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4895__A2 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6317_ _3759_ _2005_ _2010_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7297_ _2914_ _0667_ _2859_ _0775_ _2945_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6097__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7970__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7294__B1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7833__A2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ _1250_ _1557_ _0937_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _1877_ _1325_ _1859_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7597__A1 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7061__A3 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7349__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4245__B _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6021__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_27_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7521__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7521__B2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6686__I _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4886__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6088__A1 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7588__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6260__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _3529_ _3673_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7185__C _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _0344_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5481_ _0695_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6315__A2 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7220_ _2866_ _3833_ _2869_ _2873_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4432_ _0286_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5374__I0 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7993__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7151_ _2477_ _2791_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4363_ _3894_ _3897_ _3898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ _1785_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7082_ _2121_ _2735_ _2739_ _2442_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _3788_ _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A2 _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _1756_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5005__I _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7579__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7984_ _0103_ clknet_leaf_35_wb_clk_i as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6251__A1 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _1945_ _2585_ _2596_ _2479_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6866_ _2267_ _2528_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_50_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5817_ _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6797_ _2243_ _2460_ _2461_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7751__A1 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6554__A2 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4565__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4565__B2 _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5748_ _3545_ _3547_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7503__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5679_ _1484_ _3883_ _0670_ _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7418_ _2078_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4868__A2 _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5624__B _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7349_ _1413_ _2982_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6439__C _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6490__A1 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6793__A2 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7286__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7742__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4859__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5808__A1 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4167__S0 _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5284__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4664__I _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__A1 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4981_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6784__A2 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6720_ _1417_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6651_ _2309_ _2299_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6536__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5602_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8021__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6582_ _1385_ _1934_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5533_ _3671_ _1239_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5464_ _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7203_ _1819_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4415_ _3904_ _0268_ _0269_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_8183_ net46 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5395_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7215__I _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7134_ _1624_ _2789_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4346_ _3707_ _3880_ _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7065_ _1699_ _1606_ _2589_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4277_ as2650.holding_reg\[1\] _3811_ _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6016_ _1723_ _1740_ _1747_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6472__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7889__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7967_ _0086_ clknet_leaf_40_wb_clk_i as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6775__A2 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6918_ _2579_ _2566_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6722__C _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7898_ _0017_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7724__A1 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6849_ _2270_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6527__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7834__B _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4305__A4 _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5502__A3 _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4710__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4149__S0 as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__A1 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4484__I _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_42_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6766__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__A2 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7715__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7191__A2 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4200_ _3554_ _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5180_ as2650.r123_2\[2\]\[5\] _0969_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4131_ _3666_ _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4062_ _3594_ _3530_ _3597_ _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4465__B1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5662__C1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5009__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6206__A1 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7821_ _1442_ _0731_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4964_ _3913_ _0806_ _0811_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7752_ as2650.r123\[0\]\[7\] _3362_ _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6703_ _2367_ _2368_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7683_ _2723_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7706__A1 _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4895_ _0560_ _3866_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6634_ as2650.pc\[0\] net5 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7182__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6565_ _1961_ _2227_ _2229_ _2232_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_121_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5516_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7373__C _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6496_ _3570_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5447_ _1207_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5496__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5378_ _1053_ as2650.r123_2\[1\]\[5\] _1187_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7117_ _2770_ _2773_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4329_ _3532_ _3858_ _3862_ _3863_ _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_86_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8097_ _0216_ clknet_leaf_37_wb_clk_i as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6445__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7048_ _2377_ _2703_ _2706_ _2442_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8067__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7829__B _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6733__B _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4253__B _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7904__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5184__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6381__B1 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6920__A2 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7283__C _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6684__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6436__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4998__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4147__C _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4462__A3 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6643__B _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5411__A2 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__S _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3973__A2 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4680_ _0529_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6869__I _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5773__I _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7905__D _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6350_ _1380_ _2036_ _2037_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4922__A1 _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5301_ _1068_ _1073_ _1071_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6281_ _1972_ _1974_ _1977_ _1780_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7467__A3 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5232_ _0296_ _0944_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8020_ _0139_ clknet_leaf_43_wb_clk_i as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5163_ as2650.r0\[3\] as2650.r123_2\[0\]\[2\] _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4114_ _3649_ _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5094_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6978__A2 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4045_ _3580_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6109__I _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6045__S _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7804_ _3403_ _0465_ _3409_ _3410_ _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7927__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _1616_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7735_ _3355_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _0525_ _0795_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7666_ _1700_ _3094_ _3092_ _3290_ _2337_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4878_ _0356_ _3660_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7155__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6617_ as2650.stack\[3\]\[0\] _2283_ _2284_ as2650.stack\[2\]\[0\] _2285_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6902__A2 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7597_ _1981_ _0790_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4913__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6548_ _1159_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4299__I _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6479_ _2151_ _2154_ _2156_ _2157_ _2046_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5469__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7831__C _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4141__A2 _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__A1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7091__A1 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__B _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6197__A3 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7146__A2 _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5593__I _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4380__A2 _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5542__B _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4132__A2 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__A1 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7082__A1 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5768__I _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4672__I _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5850_ _1635_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7385__A2 _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6188__A3 _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4801_ _0562_ _0563_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5781_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7520_ _3147_ _3149_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4732_ _3854_ _0561_ _0583_ _3890_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5148__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7451_ _3052_ _2302_ _2366_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4663_ _3904_ _0483_ _0513_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6896__A1 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _1861_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4594_ _0344_ _0354_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7382_ _3004_ _3012_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6333_ _2022_ _2023_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6648__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6264_ _1958_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8003_ _0122_ clknet_leaf_32_wb_clk_i as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5215_ _0876_ _1050_ _0871_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6195_ _1886_ _1806_ _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_97_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5146_ _0492_ _0880_ _0975_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7073__A1 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _3713_ _3868_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7612__A3 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6820__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4028_ _3485_ as2650.cycle\[0\] _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6179__A3 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8105__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5387__A1 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5979_ _1716_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7718_ _1844_ _3322_ _3321_ _3339_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7128__A2 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7649_ _1609_ _3021_ _3270_ _1991_ _3274_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6887__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6302__I _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6887__B2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5934__I0 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4362__A2 _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7300__A2 _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5862__A2 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7064__A1 as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5614__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7289__B _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7367__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7119__A2 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6878__A1 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5550__A1 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__A1 _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7055__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6802__A1 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6951_ _1691_ _2357_ _2461_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8128__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5902_ _1667_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6882_ _1269_ _2056_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5833_ _1621_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6030__A2 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7646__C _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4041__A1 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5764_ _3515_ _1563_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7503_ _1479_ _0491_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4715_ _3521_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4592__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5695_ _1251_ _1358_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7218__I _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6122__I _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7434_ _2981_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4646_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7530__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7662__B _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5541__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7365_ _1673_ _2993_ _2998_ _1433_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4577_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5961__I _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6316_ _2005_ _2009_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7296_ _1424_ _1941_ _2944_ _1939_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_89_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4577__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7294__B2 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _1944_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6341__I0 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7833__A3 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _1789_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7046__A1 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5129_ _0936_ _0942_ _0966_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7597__A2 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6021__A2 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6572__A3 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6309__B1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7521__A2 _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7291__C _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6088__A2 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7285__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4099__A1 _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6260__A2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__A1 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7466__C _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7760__A2 _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _3920_ _3927_ _0353_ _0261_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5480_ _0445_ _0534_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4431_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5781__I _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4362_ _3724_ _3895_ _3896_ _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7150_ _1624_ _2805_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6101_ _1783_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7081_ _2737_ _2738_ _2498_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4293_ _3815_ _3820_ _3827_ _3828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _1705_ as2650.stack\[0\]\[11\] _1748_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7579__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7983_ _0102_ clknet_leaf_35_wb_clk_i as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6787__B1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6251__A2 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6934_ _1848_ _2586_ _2434_ _2595_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5021__I _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6865_ _2525_ _2527_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6561__B _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7200__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _1607_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6796_ _1430_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6554__A3 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5747_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5678_ net27 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7503__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7417_ _3031_ _3025_ _3048_ _3049_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4629_ _3783_ _3811_ _3871_ _0302_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_117_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7348_ _2981_ _3740_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7267__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ as2650.psu\[5\] _2836_ _2928_ _1395_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6490__A2 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7411__I _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4253__A1 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7742__A2 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5753__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__A1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7258__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5106__I as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__A2 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4167__S1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7430__A1 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6233__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _0820_ _3533_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4680__I _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6650_ _1942_ _2303_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7960__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5601_ _3675_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6581_ _1538_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5532_ _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5463_ _1195_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7202_ _2856_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4414_ _3784_ _3811_ _3871_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_114_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5394_ _3576_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7249__A1 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7133_ _1619_ _2753_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4345_ _3877_ _3690_ _3879_ _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7064_ as2650.pc\[10\] _2589_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4276_ _3701_ _3704_ _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_87_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6015_ as2650.stack\[0\]\[3\] _1746_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4855__I _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6472__A2 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__A1 _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5680__B1 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5887__S _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6224__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4235__A1 _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7966_ _0085_ clknet_leaf_30_wb_clk_i as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6917_ _2248_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7897_ _0016_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4590__I as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6848_ _2506_ _2509_ _2511_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7185__B1 _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7724__A2 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6779_ _2270_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4149__S1 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6466__B _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7660__A1 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A2 _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4005__I _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4130_ _3665_ _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7651__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4061_ _3596_ _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4465__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5662__B1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4465__B2 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5662__C2 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6206__A2 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7820_ _1436_ _3402_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7751_ _0713_ _3361_ _3365_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4963_ as2650.r123\[1\]\[1\] _0809_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6702_ as2650.pc\[2\] net7 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7682_ _2987_ _3296_ _3116_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4894_ _0742_ _0641_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6633_ _2299_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6564_ _1811_ _1974_ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5515_ _3530_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6495_ _1900_ _1808_ _2138_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5446_ _1211_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ _1189_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7116_ _1233_ _2772_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4328_ _3550_ _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_134_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8096_ _0215_ clknet_leaf_37_wb_clk_i as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6286__B _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7642__A1 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ _2498_ _2705_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4259_ _3755_ _3765_ _3791_ _3794_ _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__C _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7949_ _0068_ clknet_leaf_48_wb_clk_i as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5708__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A1 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__A1 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6684__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7633__A1 _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8011__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3973__A3 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _1132_ _1133_ _1074_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6280_ _1553_ _1976_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7490__B _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5231_ _3711_ as2650.r123_2\[0\]\[6\] _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7872__A1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6885__I _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__A1 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4113_ _3648_ _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_110_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6427__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5093_ _0266_ _0931_ _0829_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4044_ _3568_ _3500_ _3579_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7803_ _0363_ _0936_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4354__B _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5995_ _1732_ _1718_ _1733_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6125__I _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7734_ _0807_ _3353_ _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4946_ as2650.r123\[2\]\[7\] _0433_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7665_ _2699_ _3289_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4877_ _3776_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6616_ _2273_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7596_ _3198_ _3201_ _3222_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6547_ _1448_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6115__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6478_ _1307_ _1550_ _2151_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7863__A1 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5429_ _3528_ _3544_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8034__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7615__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7615__B2 _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8079_ _0198_ clknet_3_6_0_wb_clk_i as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4429__A1 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7091__A2 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6744__B _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6354__A1 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4953__I _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _0267_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6593__A1 _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _3857_ _0570_ _0582_ _3888_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5784__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7450_ _3074_ _3081_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4662_ _0514_ _0401_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5148__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6401_ _1987_ _2085_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7381_ _1937_ _3000_ _3002_ _1673_ _3014_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _0341_ _0363_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8057__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ _1272_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7845__A1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6648__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6263_ _3564_ _1959_ _1943_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8002_ _0121_ clknet_leaf_47_wb_clk_i as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5214_ _1009_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6194_ _1888_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5145_ _0841_ _0980_ _0981_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5024__I _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7073__A2 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5076_ _3835_ _3702_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5084__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6820__A2 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4027_ _3538_ _3562_ _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4831__A1 _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5387__A2 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5978_ _1582_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7717_ _2758_ _1914_ _1844_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4929_ _0573_ _0770_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7648_ _2503_ _3273_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6887__A2 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5934__I1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7579_ _0578_ _0558_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7836__A1 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3942__I _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5135__S _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5311__A2 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7064__A2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A3 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7524__B1 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4889__A1 _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4013__I _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5550__A2 _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7827__A1 _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7917__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__A2 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5779__I _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5066__A1 _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6950_ _2576_ _2598_ _2600_ _2611_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5901_ _1610_ as2650.stack\[4\]\[8\] _1662_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6881_ _1593_ _2543_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _1620_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6566__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5728__B _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5763_ _1549_ _1551_ _1553_ _1562_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4041__A2 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7502_ _0387_ _0379_ _3075_ _3076_ _3104_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4714_ as2650.r123\[0\]\[6\] as2650.r123_2\[0\]\[6\] as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\]
+ _3647_ _3614_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_5694_ _1205_ _1499_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7433_ _2987_ _3064_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4645_ as2650.r0\[5\] _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5019__I _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7662__C _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7364_ _2107_ _1528_ _2997_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4576_ _3749_ _0368_ _0411_ _0429_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__5541__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7818__A1 _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6315_ _2007_ _2008_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7295_ _2942_ _2943_ _1409_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7294__A2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6246_ _1943_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6341__I1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ _1875_ _1242_ _1859_ _1501_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_97_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _0943_ _0956_ _0965_ _0942_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5057__A1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5059_ _0883_ _0886_ _0897_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4804__A1 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6741__C _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6572__A4 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__A1 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6309__B2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7809__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7285__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4099__A2 _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7037__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__I _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4436__C _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4271__A2 _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6548__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6223__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ net7 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7482__C _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6720__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6379__B _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5283__B _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4361_ as2650.addr_buff\[6\] _3725_ _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_99_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6100_ _1331_ _1808_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7080_ _2314_ _2704_ _2383_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4292_ _3821_ _3823_ _3824_ _3826_ _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5287__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6031_ _1734_ _1741_ _1755_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4334__I0 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A4 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7003__B _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7982_ _0101_ clknet_leaf_34_wb_clk_i as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6787__A1 as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__B2 as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _2592_ _2594_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6251__A3 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _1586_ _0976_ _2526_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6539__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6561__C _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5815_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6003__A3 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6795_ _2415_ _2424_ _2458_ _2459_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6554__A4 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5746_ _1545_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7673__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5677_ as2650.psu\[1\] _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7416_ _1796_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4628_ _3746_ _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7347_ _3736_ _3734_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4559_ _3840_ _0330_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7267__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7278_ _1457_ _2878_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6229_ _3579_ _3692_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6778__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5450__A1 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__C _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5087__C _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5753__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7583__B _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6702__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5505__A2 _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5269__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5122__I _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4244__A2 _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7194__A1 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5600_ _1407_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6580_ _1519_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5531_ _3593_ _3499_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5792__I _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ _1270_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7201_ _2843_ _2850_ _2855_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4413_ _3689_ _3705_ _3929_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5393_ _1195_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7249__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7132_ _2296_ _2788_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4344_ _3690_ _3878_ _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7063_ _2305_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ _3808_ _3809_ _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6014_ _1739_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4357__B _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5680__A1 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5680__B2 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7421__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7965_ _0084_ clknet_leaf_30_wb_clk_i as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4235__A2 _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6916_ _1597_ _2577_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7896_ _0015_ clknet_leaf_58_wb_clk_i as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7185__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6847_ as2650.stack\[1\]\[4\] _2402_ _2510_ as2650.stack\[2\]\[4\] _2511_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7185__B2 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6932__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6778_ _2377_ _2433_ _2441_ _2442_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5729_ _1271_ _1523_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4111__I _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6747__B _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6999__A1 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4474__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6038__I _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4226__A2 _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5423__A1 _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__B1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7297__C _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7176__A1 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6923__A1 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6923__B2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6501__I _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6151__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8090__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5561__B _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6149__S _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7100__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6376__C _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4060_ _3595_ _3580_ _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4465__A2 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5662__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5662__B2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7403__A2 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5787__I _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5414__A1 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6611__B1 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7750_ as2650.r123\[0\]\[6\] _3362_ _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4962_ _3798_ _0806_ _0810_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6701_ _2301_ _2302_ _2366_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7681_ _3114_ _3304_ _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4893_ _0639_ _0640_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7167__A1 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6632_ _1570_ _1536_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6563_ _0311_ _2230_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5514_ _1255_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6494_ _3591_ _1807_ _2167_ _1330_ _2170_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_133_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5445_ _1248_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5376_ _1013_ as2650.r123_2\[1\]\[4\] _1187_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7115_ _2440_ _2771_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4327_ _3861_ _3614_ _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6059__S _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8095_ _0214_ clknet_leaf_41_wb_clk_i as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7046_ _2314_ _2704_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7642__A2 _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4258_ _3792_ _3793_ _3755_ _3794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6850__B1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4189_ as2650.addr_buff\[5\] _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5697__I _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7948_ _0067_ clknet_leaf_32_wb_clk_i as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7879_ as2650.psu\[0\] _3474_ _3475_ _3461_ _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4106__I _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3945__I _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6381__A2 _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4392__A1 _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6669__B1 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7330__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6477__B _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5644__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7397__A1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5400__I _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5230_ _1034_ _1037_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5883__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5161_ _0390_ as2650.r123_2\[0\]\[0\] _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4112_ _3647_ _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7624__A2 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5092_ _0920_ _0922_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ as2650.ins_reg\[4\] _3558_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7388__A1 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7802_ _0363_ _0936_ _3406_ _3407_ _3408_ _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6406__I _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5994_ as2650.stack\[5\]\[9\] _1720_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7733_ _3353_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4945_ _3751_ _0741_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7664_ _2493_ _3281_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4876_ _0721_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ _1649_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7595_ _0670_ _0679_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6546_ _1113_ _1196_ _2213_ _2214_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7312__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6115__A2 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6477_ _0973_ _2155_ _2138_ _1440_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7973__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5428_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7863__A2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4596__I _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5359_ _1178_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8078_ _0197_ clknet_leaf_28_wb_clk_i as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7615__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7029_ _2648_ _2687_ _2688_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5220__I _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6760__B _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4601__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6354__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7303__A1 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4117__A1 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6935__B _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6654__C _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4730_ _3669_ _0576_ _0581_ _3886_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4661_ _3738_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7542__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6400_ _2046_ _2047_ _1254_ _2084_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4356__A1 _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7996__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7380_ _3013_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4592_ _0442_ _0444_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6331_ _1421_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7932__D _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6262_ _3671_ _3547_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7845__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4659__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ _1029_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8001_ _0120_ clknet_leaf_47_wb_clk_i as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6193_ _1816_ _1889_ _1890_ _1804_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_97_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5144_ _0307_ _0842_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5075_ _0828_ _0913_ _0914_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5084__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4026_ _3543_ _3548_ _3561_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4831__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5977_ _1722_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7781__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7716_ net40 _3337_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4928_ _0719_ _0573_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7647_ _1608_ _2993_ _3271_ _3272_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4859_ _0435_ _0685_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7578_ _0578_ _0558_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4898__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6529_ net45 _2192_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7836__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5847__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7049__B1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5075__A2 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A4 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4822__A2 _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7586__B _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7772__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__A1 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6649__C _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4510__A1 _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5066__A2 _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6263__A1 _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5900_ _1604_ _1655_ _1666_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6880_ _1587_ _2480_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5831_ _1619_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6566__A2 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8024__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5762_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4041__A3 _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7501_ _0387_ _0379_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_6_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4713_ _0564_ _3616_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7515__A1 _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5693_ _3779_ _1498_ _0821_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4329__A1 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7432_ _3060_ _3063_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _3875_ _0494_ _0496_ _3886_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7363_ _2333_ _2254_ _2995_ _2996_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_116_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4575_ _0412_ _0427_ _0428_ _0333_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5541__A3 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6314_ _1413_ _1439_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7294_ _1398_ _1101_ _0663_ _1392_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5829__A1 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _1942_ _1818_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6176_ _0939_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5127_ _0376_ _0856_ _0869_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6067__S _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5058_ _0839_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4804__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4009_ _3527_ _3544_ _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6557__A2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7754__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7506__A1 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4114__I _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7809__A2 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5048__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6245__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8047__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4733__B _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6548__A2 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7760__A4 _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5508__B1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6720__A2 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ _3726_ _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4291_ _3549_ _3707_ _3825_ _3771_ _3826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6030_ as2650.stack\[0\]\[10\] _1743_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4334__I1 _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6236__A1 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7981_ _0100_ clknet_leaf_43_wb_clk_i as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6787__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6932_ _2427_ _2593_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6863_ _2468_ _2470_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7736__A1 _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5814_ as2650.pc\[8\] _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6794_ _2126_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5211__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5745_ _1543_ _1544_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5676_ net1 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7415_ _3039_ _3046_ _3047_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4869__I _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4627_ _0428_ _0478_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7346_ _1413_ _2979_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _3539_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4489_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7277_ _1392_ _0449_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6475__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6228_ _1552_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6159_ _1854_ _1859_ _1330_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_112_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6227__A1 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7424__B1 _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4789__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5450__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7727__A1 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6324__I _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7907__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7864__B _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4961__A1 as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6702__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5505__A3 _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4713__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput40 net40 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7718__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7194__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4952__A1 _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5530_ _3512_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5461_ _1269_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4412_ _3516_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7200_ _2171_ _2854_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4704__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4343_ _3566_ _3560_ _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7131_ _1621_ _2298_ _2787_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7062_ _1702_ _2719_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4274_ _3770_ _3506_ _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6013_ _1745_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6209__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5680__A2 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6345__S _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7964_ _0083_ clknet_leaf_40_wb_clk_i as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6915_ _1688_ _1586_ _2480_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7709__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7895_ _0014_ clknet_leaf_58_wb_clk_i as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6846_ _2284_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7185__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _1505_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3989_ as2650.cycle\[1\] _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5728_ _1503_ _1522_ _1530_ _1214_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_108_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5659_ _3542_ _3814_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7329_ as2650.stack\[7\]\[5\] _2967_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6999__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output44_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5423__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A4 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7176__A2 _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4302__I as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6687__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6687__B2 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6439__A1 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5662__A2 _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5289__B _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ as2650.r123\[1\]\[0\] _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ as2650.pc\[1\] _3882_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7680_ _3299_ _3300_ _3301_ _3303_ as2650.addr_buff\[2\] _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_127_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7167__A2 _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4892_ _0639_ _0640_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5178__A1 as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6631_ _2297_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6562_ _1788_ _1973_ _1552_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7009__B _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5513_ _1302_ _1306_ _1317_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6493_ _1778_ _2168_ _2169_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__6678__A1 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5444_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5375_ _1188_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7114_ _1841_ _2327_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4326_ _3860_ _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8094_ _0213_ clknet_leaf_37_wb_clk_i as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6139__I as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7045_ as2650.addr_buff\[0\] _2663_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4257_ _3782_ _3788_ _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5043__I _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6850__B2 as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4188_ _3688_ _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5978__I _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6602__A1 as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8108__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7947_ _0066_ clknet_leaf_32_wb_clk_i as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7878_ _3458_ _2008_ _2007_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6829_ _1810_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4831__B _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A2 _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6669__B2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3961__I _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6477__C _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5644__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6512__I _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7771__C _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5160_ _3834_ _0944_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5999__S _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7085__A1 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4111_ _3477_ _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_111_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5091_ _0277_ _0859_ _0862_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4042_ _3507_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7388__A2 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7801_ _0265_ _0353_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5993_ _1613_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4207__I as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7732_ _1158_ _1159_ _0412_ _0801_ _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_40_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _3517_ _0767_ _0793_ _3751_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4071__A1 _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7663_ _3049_ _3279_ _3287_ _2939_ _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4651__B _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4875_ _0692_ _0696_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7518__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6899__A1 _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6614_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7594_ _3219_ _3220_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7560__A2 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6545_ _2015_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _3591_ _2154_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7312__A2 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4877__I _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5323__A1 as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4126__A2 as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _1235_ _3848_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7863__A3 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ as2650.r123\[3\]\[5\] _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7076__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4309_ _3843_ _3745_ _3839_ _3742_ _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8077_ _0196_ clknet_leaf_28_wb_clk_i as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5289_ _0774_ _0879_ _0862_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6823__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6823__B2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7028_ _2044_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5501__I _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7379__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4062__A1 _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6760__C _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7428__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6332__I _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5937__I0 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5562__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7303__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5314__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4117__A2 _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6935__C _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4455__C _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A2 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__I _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4660_ _0485_ _0486_ _3903_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7542__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7782__B _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5553__A1 _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _0443_ _0401_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6330_ _2020_ _2011_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5305__A1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6261_ _1957_ _1501_ _1553_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8000_ _0119_ clknet_leaf_44_wb_clk_i as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5212_ _0994_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7006__C _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6192_ _1803_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7058__A1 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7058__B2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5143_ _0663_ _0890_ _0891_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5069__B1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5074_ as2650.r123_2\[2\]\[1\] _0875_ _0877_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4025_ _3549_ _3553_ _3556_ _3560_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__6281__A2 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4292__A1 _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7230__A1 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7230__B2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__A1 _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5976_ _1579_ as2650.stack\[5\]\[2\] _1720_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7781__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7715_ net39 _3317_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4595__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4927_ _3877_ _0664_ _0654_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6152__I _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7646_ _2586_ _3267_ _3091_ _2668_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7940__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4858_ _3939_ _0705_ _0708_ _0338_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7577_ _1455_ _0659_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4789_ _0499_ _3837_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6528_ _2028_ _2181_ _2200_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__A1 _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7297__B2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _1970_ _1971_ _1926_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A2 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7049__A1 as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8129_ _0248_ clknet_leaf_10_wb_clk_i as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4556__B _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6024__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7586__C _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4035__A1 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7772__A2 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6980__B1 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__A2 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7288__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4510__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6665__C _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4649__I0 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6263__A2 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4274__A1 _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6015__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ as2650.pc\[11\] _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4026__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7963__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5761_ _1554_ _1559_ _1560_ _0547_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7500_ _3127_ _3129_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ as2650.r0\[6\] _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5692_ _1234_ _3566_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7515__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7431_ net52 _2988_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5526__A1 _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _0495_ _3884_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7362_ _2988_ _2427_ _2257_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4574_ _0413_ _0426_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7279__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6313_ _0865_ _2006_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7293_ _1388_ _1231_ _2941_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5829__A2 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6244_ _3569_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6175_ _1375_ _1873_ _1367_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _0380_ _0838_ _0855_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4376__B _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5051__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5057_ _0887_ _0890_ _0891_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4265__A1 as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4265__B2 _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4008_ _3485_ as2650.cycle\[0\] _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7754__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5959_ as2650.stack\[1\]\[12\] _1707_ _1676_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7629_ _3252_ _3254_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5517__A1 _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4130__I _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7690__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6493__A2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7442__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__A2 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5508__A1 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__B2 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__A1 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4731__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ _3803_ _3549_ _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7130__B1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7681__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A1 _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7433__A1 _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6236__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7980_ _0099_ clknet_leaf_33_wb_clk_i as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6931_ _2591_ _2555_ _2588_ _2590_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__5995__A1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _1592_ _0577_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7736__A2 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5813_ _1604_ _1568_ _1605_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8141__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6793_ _2423_ _2443_ _2457_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5744_ as2650.stack_ptr\[0\] _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5675_ as2650.psu\[2\] _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7414_ _1919_ _1890_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6430__I _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4626_ _0428_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7345_ _1023_ _3731_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4557_ _0369_ _0376_ _0410_ _0267_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7276_ _2923_ _2924_ _2869_ _2925_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7121__B1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4488_ as2650.holding_reg\[3\] _0304_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5490__B _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7672__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6227_ _1894_ _1904_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6158_ _3578_ _3570_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7424__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _3699_ _3867_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6089_ _1778_ _1781_ _1792_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A1 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4789__A2 _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7727__A2 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4125__I _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4961__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6163__A1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4713__A2 _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput30 net30 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6466__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7663__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7171__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__A1 _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8014__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6218__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__A1 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7194__A3 _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4401__A1 _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5460_ _0579_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6154__A1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _0265_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4704__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _3536_ _1196_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_114_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7130_ _2503_ _2755_ _2777_ _2786_ _2297_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4342_ _3540_ _3876_ _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7654__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6457__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7061_ _1699_ _1606_ _2658_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4273_ _3807_ _3808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4468__A1 _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _1681_ as2650.stack\[0\]\[2\] _1743_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
.ends

