* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuD

* Black-box entry subcircuit for timers abstract view
.subckt timers addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] bus_cyc bus_we data_in[0]
+ data_in[1] data_in[2] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7] data_out[0]
+ data_out[1] data_out[2] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7]
+ irq1 irq2 irq5 pwm0 pwm1 pwm2 rst tmr0_clk tmr0_o tmr1_clk tmr1_o vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for avali_logo abstract view
.subckt avali_logo vss vdd
.ends

* Black-box entry subcircuit for sid_top abstract view
.subckt sid_top DAC_clk DAC_dat_1 DAC_dat_2 DAC_le addr[0] addr[1] addr[2] addr[3]
+ addr[4] bus_cyc bus_in[0] bus_in[1] bus_in[2] bus_in[3] bus_in[4] bus_in[5] bus_in[6]
+ bus_in[7] bus_out[0] bus_out[1] bus_out[2] bus_out[3] bus_out[4] bus_out[5] bus_out[6]
+ bus_out[7] bus_we clk rst vdd vss
.ends

* Black-box entry subcircuit for gpios abstract view
.subckt gpios DAC_clk DAC_d1 DAC_d2 DAC_le RXD TXD addr[0] addr[1] addr[2] addr[3]
+ bus_cyc bus_we data_in[0] data_in[1] data_in[2] data_in[3] data_in[4] data_in[5]
+ data_in[6] data_in[7] data_out[0] data_out[1] data_out[2] data_out[3] data_out[4]
+ data_out[5] data_out[6] data_out[7] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] irq0 irq6 irq7 la_data_out[0] la_data_out[1] la_data_out[2]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] pwm0
+ pwm1 pwm2 rst tmr0_clk tmr0_o tmr1_clk tmr1_o vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for serial_ports abstract view
.subckt serial_ports RXD TXD addr[0] addr[1] addr[2] bus_cyc bus_we data_in[0] data_in[1]
+ data_in[2] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7] data_out[0] data_out[1]
+ data_out[2] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7] io_in io_oeb[0]
+ io_oeb[1] io_oeb[2] io_out[0] io_out[1] io_out[2] irq3 rst vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for boot_rom abstract view
.subckt boot_rom WEb_raw bus_in[0] bus_in[1] bus_in[2] bus_in[3] bus_in[4] bus_in[5]
+ bus_in[6] bus_in[7] bus_out[0] bus_out[1] bus_out[2] bus_out[3] bus_out[4] bus_out[5]
+ bus_out[6] bus_out[7] cs_port[0] cs_port[1] cs_port[2] le_hi_act le_lo_act ram_end[0]
+ ram_end[10] ram_end[11] ram_end[12] ram_end[13] ram_end[14] ram_end[15] ram_end[1]
+ ram_end[2] ram_end[3] ram_end[4] ram_end[5] ram_end[6] ram_end[7] ram_end[8] ram_end[9]
+ ram_start[0] ram_start[10] ram_start[11] ram_start[12] ram_start[13] ram_start[14]
+ ram_start[15] ram_start[1] ram_start[2] ram_start[3] ram_start[4] ram_start[5] ram_start[6]
+ ram_start[7] ram_start[8] ram_start[9] rom_enabled rst vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for wrapped_as2650 abstract view
.subckt wrapped_as2650 RAM_end_addr[0] RAM_end_addr[10] RAM_end_addr[11] RAM_end_addr[12]
+ RAM_end_addr[13] RAM_end_addr[14] RAM_end_addr[15] RAM_end_addr[1] RAM_end_addr[2]
+ RAM_end_addr[3] RAM_end_addr[4] RAM_end_addr[5] RAM_end_addr[6] RAM_end_addr[7]
+ RAM_end_addr[8] RAM_end_addr[9] RAM_start_addr[0] RAM_start_addr[10] RAM_start_addr[11]
+ RAM_start_addr[12] RAM_start_addr[13] RAM_start_addr[14] RAM_start_addr[15] RAM_start_addr[1]
+ RAM_start_addr[2] RAM_start_addr[3] RAM_start_addr[4] RAM_start_addr[5] RAM_start_addr[6]
+ RAM_start_addr[7] RAM_start_addr[8] RAM_start_addr[9] WEb_raw boot_rom_en bus_addr[0]
+ bus_addr[1] bus_addr[2] bus_addr[3] bus_addr[4] bus_addr[5] bus_cyc bus_data_out[0]
+ bus_data_out[1] bus_data_out[2] bus_data_out[3] bus_data_out[4] bus_data_out[5]
+ bus_data_out[6] bus_data_out[7] bus_in_gpios[0] bus_in_gpios[1] bus_in_gpios[2]
+ bus_in_gpios[3] bus_in_gpios[4] bus_in_gpios[5] bus_in_gpios[6] bus_in_gpios[7]
+ bus_in_serial_ports[0] bus_in_serial_ports[1] bus_in_serial_ports[2] bus_in_serial_ports[3]
+ bus_in_serial_ports[4] bus_in_serial_ports[5] bus_in_serial_ports[6] bus_in_serial_ports[7]
+ bus_in_sid[0] bus_in_sid[1] bus_in_sid[2] bus_in_sid[3] bus_in_sid[4] bus_in_sid[5]
+ bus_in_sid[6] bus_in_sid[7] bus_in_timers[0] bus_in_timers[1] bus_in_timers[2] bus_in_timers[3]
+ bus_in_timers[4] bus_in_timers[5] bus_in_timers[6] bus_in_timers[7] bus_we_gpios
+ bus_we_serial_ports bus_we_sid bus_we_timers cs_port[0] cs_port[1] cs_port[2] io_in[0]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8]
+ io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[1] io_out[2]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1]
+ irq[2] irqs[0] irqs[1] irqs[2] irqs[3] irqs[4] irqs[5] irqs[6] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] le_hi_act
+ le_lo_act reset_out rom_bus_in[0] rom_bus_in[1] rom_bus_in[2] rom_bus_in[3] rom_bus_in[4]
+ rom_bus_in[5] rom_bus_in[6] rom_bus_in[7] rom_bus_out[0] rom_bus_out[1] rom_bus_out[2]
+ rom_bus_out[3] rom_bus_out[4] rom_bus_out[5] rom_bus_out[6] rom_bus_out[7] vdd vss
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_stb_i wbs_we_i
.ends

.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xtimers bus_addr\[0\] bus_addr\[1\] bus_addr\[2\] bus_addr\[3\] bus_addr\[4\] bus_addr\[5\]
+ bus_cyc bus_we_timers bus_data_out\[0\] bus_data_out\[1\] bus_data_out\[2\] bus_data_out\[3\]
+ bus_data_out\[4\] bus_data_out\[5\] bus_data_out\[6\] bus_data_out\[7\] bus_data_timers\[0\]
+ bus_data_timers\[1\] bus_data_timers\[2\] bus_data_timers\[3\] bus_data_timers\[4\]
+ bus_data_timers\[5\] bus_data_timers\[6\] bus_data_timers\[7\] irq1 irq2 irq5 pwm0
+ pwm1 pwm2 reset tmr0_clk tmr0_o tmr1_clk tmr1_o vdd vss wb_clk_i timers
Xavali_logo vss vdd avali_logo
Xsid DAC_clk DAC_d1 DAC_d2 DAC_le bus_addr\[0\] bus_addr\[1\] bus_addr\[2\] bus_addr\[3\]
+ bus_addr\[4\] bus_cyc bus_data_out\[0\] bus_data_out\[1\] bus_data_out\[2\] bus_data_out\[3\]
+ bus_data_out\[4\] bus_data_out\[5\] bus_data_out\[6\] bus_data_out\[7\] bus_data_sid\[0\]
+ bus_data_sid\[1\] bus_data_sid\[2\] bus_data_sid\[3\] bus_data_sid\[4\] bus_data_sid\[5\]
+ bus_data_sid\[6\] bus_data_sid\[7\] bus_we_sid wb_clk_i reset vdd vss sid_top
Xgpios DAC_clk DAC_d1 DAC_d2 DAC_le RXD TXD bus_addr\[0\] bus_addr\[1\] bus_addr\[2\]
+ bus_addr\[3\] bus_cyc bus_we_gpios bus_data_out\[0\] bus_data_out\[1\] bus_data_out\[2\]
+ bus_data_out\[3\] bus_data_out\[4\] bus_data_out\[5\] bus_data_out\[6\] bus_data_out\[7\]
+ bus_data_gpios\[0\] bus_data_gpios\[1\] bus_data_gpios\[2\] bus_data_gpios\[3\]
+ bus_data_gpios\[4\] bus_data_gpios\[5\] bus_data_gpios\[6\] bus_data_gpios\[7\]
+ io_in[19] io_in[29] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[20]
+ io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28]
+ io_oeb[19] io_oeb[29] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_out[19] io_out[29] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28]
+ irq0 irq6 irq7 la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] pwm0 pwm1 pwm2 reset tmr0_clk tmr0_o
+ tmr1_clk tmr1_o vdd vss wb_clk_i gpios
Xserial_ports RXD TXD bus_addr\[0\] bus_addr\[1\] bus_addr\[2\] bus_cyc bus_we_serial_ports
+ bus_data_out\[0\] bus_data_out\[1\] bus_data_out\[2\] bus_data_out\[3\] bus_data_out\[4\]
+ bus_data_out\[5\] bus_data_out\[6\] bus_data_out\[7\] bus_data_serial_ports\[0\]
+ bus_data_serial_ports\[1\] bus_data_serial_ports\[2\] bus_data_serial_ports\[3\]
+ bus_data_serial_ports\[4\] bus_data_serial_ports\[5\] bus_data_serial_ports\[6\]
+ bus_data_serial_ports\[7\] io_in[37] io_oeb[35] io_oeb[36] io_oeb[37] io_out[35]
+ io_out[36] io_out[37] irq3 reset vdd vss wb_clk_i serial_ports
Xboot_rom WEb_raw rom_bus_out\[0\] rom_bus_out\[1\] rom_bus_out\[2\] rom_bus_out\[3\]
+ rom_bus_out\[4\] rom_bus_out\[5\] rom_bus_out\[6\] rom_bus_out\[7\] rom_bus_in\[0\]
+ rom_bus_in\[1\] rom_bus_in\[2\] rom_bus_in\[3\] rom_bus_in\[4\] rom_bus_in\[5\]
+ rom_bus_in\[6\] rom_bus_in\[7\] cs_port\[0\] cs_port\[1\] cs_port\[2\] le_hi_act
+ le_lo_act RAM_end_addr\[0\] RAM_end_addr\[10\] RAM_end_addr\[11\] RAM_end_addr\[12\]
+ RAM_end_addr\[13\] RAM_end_addr\[14\] RAM_end_addr\[15\] RAM_end_addr\[1\] RAM_end_addr\[2\]
+ RAM_end_addr\[3\] RAM_end_addr\[4\] RAM_end_addr\[5\] RAM_end_addr\[6\] RAM_end_addr\[7\]
+ RAM_end_addr\[8\] RAM_end_addr\[9\] RAM_start_addr\[0\] RAM_start_addr\[10\] RAM_start_addr\[11\]
+ RAM_start_addr\[12\] RAM_start_addr\[13\] RAM_start_addr\[14\] RAM_start_addr\[15\]
+ RAM_start_addr\[1\] RAM_start_addr\[2\] RAM_start_addr\[3\] RAM_start_addr\[4\]
+ RAM_start_addr\[5\] RAM_start_addr\[6\] RAM_start_addr\[7\] RAM_start_addr\[8\]
+ RAM_start_addr\[9\] boot_rom_en reset vdd vss wb_clk_i boot_rom
Xwrapped_as2650 RAM_end_addr\[0\] RAM_end_addr\[10\] RAM_end_addr\[11\] RAM_end_addr\[12\]
+ RAM_end_addr\[13\] RAM_end_addr\[14\] RAM_end_addr\[15\] RAM_end_addr\[1\] RAM_end_addr\[2\]
+ RAM_end_addr\[3\] RAM_end_addr\[4\] RAM_end_addr\[5\] RAM_end_addr\[6\] RAM_end_addr\[7\]
+ RAM_end_addr\[8\] RAM_end_addr\[9\] RAM_start_addr\[0\] RAM_start_addr\[10\] RAM_start_addr\[11\]
+ RAM_start_addr\[12\] RAM_start_addr\[13\] RAM_start_addr\[14\] RAM_start_addr\[15\]
+ RAM_start_addr\[1\] RAM_start_addr\[2\] RAM_start_addr\[3\] RAM_start_addr\[4\]
+ RAM_start_addr\[5\] RAM_start_addr\[6\] RAM_start_addr\[7\] RAM_start_addr\[8\]
+ RAM_start_addr\[9\] WEb_raw boot_rom_en bus_addr\[0\] bus_addr\[1\] bus_addr\[2\]
+ bus_addr\[3\] bus_addr\[4\] bus_addr\[5\] bus_cyc bus_data_out\[0\] bus_data_out\[1\]
+ bus_data_out\[2\] bus_data_out\[3\] bus_data_out\[4\] bus_data_out\[5\] bus_data_out\[6\]
+ bus_data_out\[7\] bus_data_gpios\[0\] bus_data_gpios\[1\] bus_data_gpios\[2\] bus_data_gpios\[3\]
+ bus_data_gpios\[4\] bus_data_gpios\[5\] bus_data_gpios\[6\] bus_data_gpios\[7\]
+ bus_data_serial_ports\[0\] bus_data_serial_ports\[1\] bus_data_serial_ports\[2\]
+ bus_data_serial_ports\[3\] bus_data_serial_ports\[4\] bus_data_serial_ports\[5\]
+ bus_data_serial_ports\[6\] bus_data_serial_ports\[7\] bus_data_sid\[0\] bus_data_sid\[1\]
+ bus_data_sid\[2\] bus_data_sid\[3\] bus_data_sid\[4\] bus_data_sid\[5\] bus_data_sid\[6\]
+ bus_data_sid\[7\] bus_data_timers\[0\] bus_data_timers\[1\] bus_data_timers\[2\]
+ bus_data_timers\[3\] bus_data_timers\[4\] bus_data_timers\[5\] bus_data_timers\[6\]
+ bus_data_timers\[7\] bus_we_gpios bus_we_serial_ports bus_we_sid bus_we_timers cs_port\[0\]
+ cs_port\[1\] cs_port\[2\] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[1] io_oeb[2] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8]
+ io_out[9] user_irq[0] user_irq[1] user_irq[2] irq0 irq1 irq2 irq3 irq5 irq6 irq7
+ la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9]
+ le_hi_act le_lo_act reset rom_bus_in\[0\] rom_bus_in\[1\] rom_bus_in\[2\] rom_bus_in\[3\]
+ rom_bus_in\[4\] rom_bus_in\[5\] rom_bus_in\[6\] rom_bus_in\[7\] rom_bus_out\[0\]
+ rom_bus_out\[1\] rom_bus_out\[2\] rom_bus_out\[3\] rom_bus_out\[4\] rom_bus_out\[5\]
+ rom_bus_out\[6\] rom_bus_out\[7\] vdd vss wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i wbs_we_i wrapped_as2650
.ends

